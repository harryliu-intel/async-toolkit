// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

// vim: noai : ts=3 : sw=3 : expandtab : ft=systemverilog

//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors.  The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//   Author        : Dhivya Sankar
//   Project       : Madison Bay
//------------------------------------------------------------------------------

//
`timescale 1ps/1ps

// Module: mby_mesh_tb_top
// Mesh testbench module
// Description :
//   This top module will:
//   1. Instance 1 RTL Unit
//   2. Control Dumping features for FSDB/DVE.

module mby_mesh_tb_top();
   
   import uvm_pkg::*;
   `include "uvm_macros.svh"


   // =============================================== 
   // Clock block instance
   // ===============================================

   logic         fabric_clk;                             // Fabric Clock - 1.2 Ghz
   logic         mclk; 
   shdv_clk_gen  fabric_clk_gen(fabric_clk);
   shdv_clk_gen  mclk_gen(mclk);
   wire          tb_reset;
   wire          ref_clk;


   initial begin

      mclk_gen.period           = 555555fs; //1.8 GHz mesh clock
      mclk_gen.jitter           = 0ps;
      fabric_clk_gen.period     = 833333fs; //1.2 GHz core clock
      fabric_clk_gen.jitter     = 0ps;

   end

   // ===============================================
   // =                FSDB variable                =
   // ===============================================
   string       fsdb_file = "dump";
   int          fsdb_config_file;
   longint      fsdb_on,fsdb_off;
   int          fsdb_file_size = 1800;
   string       str;

   mby_mesh_tb_if mesh_tb_if();
 
 
   assign mesh_tb_if.fab_clk  = fabric_clk;
   assign mesh_tb_if.mclk     = mclk;

   assign ref_clk  = fabric_clk;
   assign tb_reset = mesh_tb_if.chard_reset;


   
   //MGP --> Msh write wb
   mby_mgp_rreq_if      rreq_wb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_req           ()
   );

   //MGP --> Msh Read eb
   mby_mgp_rreq_if      rreq_eb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_req           ()
   );
   // MGP --> Msh write wb
   mby_mgp_wreq_if      wreq_wb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .wr_req           ()
   );

   //MGP --> Msh write eb
   mby_mgp_wreq_if      wreq_eb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .wr_req           ()
   );

   //MGP --> Msh rsp wb
   mby_mgp_rsp_if       rsp_wb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_rsp           ()
   );

   //MGP --> Msh rsp eb
   mby_mgp_rsp_if       rsp_eb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_rsp           ()
   );


   //MGP --> Msh read sb
   mby_mgp_rreq_if      rreq_sb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_req           ()
   );

   //MGP --> Msh Read nb
   mby_mgp_rreq_if      rreq_nb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_req           ()
   );
   // MGP --> Msh write sb
   mby_mgp_wreq_if      wreq_sb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .wr_req           ()
   );

   //MGP --> Msh write nb
   mby_mgp_wreq_if      wreq_nb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .wr_req           ()
   );

   //MGP --> Msh rsp sb
   mby_mgp_rsp_if       rsp_sb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_rsp           ()
   );

   //MGP --> Msh rsp nb
   mby_mgp_rsp_if       rsp_nb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .rd_rsp           ()
   );

   //MGP --> Msh wrdata eb
   mby_mgp_data_if      wrdata_eb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data         ()
   );

   //MGP --> Msh wrdata wb
   mby_mgp_data_if      wrdata_wb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data         ()
   );

   //MGP --> Msh wrdata sb
   mby_mgp_data_if      wrdata_sb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data         ()
   );

   //MGP --> Msh wrdata nb
   mby_mgp_data_if      wrdata_nb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data         ()
   );

   //MGP --> Msh rddata eb
   mby_mgp_data_if      rddata_eb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data         ()
   );

   //MGP --> Msh rddata wb
   mby_mgp_data_if      rddata_wb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data         ()
   );

   //MGP --> Msh rddata sb
   mby_mgp_data_if      rddata_sb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data          ()
   );

   //MGP --> Msh rddata nb
   mby_mgp_data_if      rddata_nb_if (
      .cclk             (ref_clk),
      .reset            (tb_reset),
      .req_data         ()
   );
   //-----------------------------------------------------------------------------
   // Verification Test Island
   //-----------------------------------------------------------------------------
   mby_mesh_ti #(
   ) mesh_ti(
       .mby_mesh_tb_if               (mesh_tb_if),
       .rreq_eb_if                   (rreq_eb_if),
       .rreq_wb_if                   (rreq_wb_if),
       .wreq_eb_if                   (wreq_eb_if),
       .wreq_wb_if                   (wreq_wb_if),
       .rsp_eb_if                    (rsp_eb_if),
       .rsp_wb_if                    (rsp_wb_if),
       .rreq_sb_if                   (rreq_sb_if),
       .rreq_nb_if                   (rreq_nb_if),
       .wreq_sb_if                   (wreq_sb_if),
       .wreq_nb_if                   (wreq_nb_if),
       .rsp_sb_if                    (rsp_sb_if),
       .rsp_nb_if                    (rsp_nb_if),
       .wrdata_eb_if                 (wrdata_eb_if),
       .wrdata_wb_if                 (wrdata_wb_if),
       .wrdata_sb_if                 (wrdata_sb_if),
       .wrdata_nb_if                 (wrdata_nb_if),
       .rddata_eb_if                 (rddata_eb_if),
       .rddata_wb_if                 (rddata_wb_if),
       .rddata_sb_if                 (rddata_sb_if),
       .rddata_nb_if                 (rddata_nb_if)
 
   );


   //////////////////////////////////////////////
   // Hierarchy-Based RTL File List Dumping ////
   /////////////////////////////////////////////

   `include  "std_ace_util.vic"

   initial begin
      dump_hier();
   end

   initial begin
      dump_vcd();
   end

   initial begin
      dump_fsdb();
   end

   initial begin
      if ($test$plusargs("vpd")) begin                                      // Plusarg to Enable VPD dump of all signals in the design
         $vcdpluson();
         $vcdplusmemon();
      end

      if($test$plusargs("fsdb")) begin                                      // Plusarg to enable FSDB dump
         if ($value$plusargs("FSDB_ON=%s",str)) begin                       // Plusarg to enable a start sample time after a delay
            fsdb_on = convert_time(str);                                    // Time to start (Converted time via plusarg)
            $display("FSDB DUMP:  Waiting %s before starting fsdb dump", str);
            #fsdb_on;                                                       // Wait - time before start
         end else begin
            fsdb_on = 0;                                                    // Time to start (no specified Time, so start at 0)
         end

         if ($value$plusargs("FSDB_SIZE=%d",fsdb_file_size)) begin               // Plusarg to specify a FSDB dump file size Limit
            if (fsdb_file_size<32) begin                                         // Must be at least 32
               fsdb_file_size = 32;
            end
         end

         $value$plusargs("FSDB_FILE=%s",fsdb_file);                         // Plusarg to specify user defined FSDB dump file name

         $fsdbAutoSwitchDumpfile(fsdb_file_size,fsdb_file,0,{fsdb_file,"_vf.log"}); // Enablement of Auto file switching

         if ($test$plusargs("fsdb_config")) begin                           // Plusarg to indicate a FSDB.dump.config file will be used. It indicates which modules to sample.
            $fsdbDumpvarsToFile ("fsdb.dump.config");
         end else begin
            $fsdbDumpvars(0,mby_mesh_tb_top,"+all");                         // Default - FSDB dump of all signals in the design
         end

         if ($value$plusargs("FSDB_OFF=%s",str)) begin                      // Plusarg to Enable a stop time of sampling
            fsdb_off = convert_time(str) - fsdb_on;                         // Overall Time to stop, not a length of time. (Converted time via plusarg, subtract Start time)
            $display("FSDB DUMP:  Stopping FSDB dump in %s", str);
            if (fsdb_off>0) begin                                           // calculated difference must be greater than 0, else stop immediately
               #fsdb_off;                                                   // Wait - time before stop
            end
            $fsdbDumpoff();                                                 // Turn off FSDB dumping
            $display("FSDB DUMP :  Stopped FSDB dump");
            fsdb_on = -1; //fsdb is off
         end
      end // if ($test$plusargs("fsdb"))
   end // initial begin
   

   function automatic longint convert_time(string in);
      longint out = in.atoi();

      case (in.substr(in.len()-2, in.len()-1))
         "ms": out *= 1000000000; // ONE BILLION ps steps in a ms unit
         "us": out *= 1000000;    // ONE MILLION ps steps in a us unit
         "ns": out *= 1000;       // ONE THOUSAND ps steps in a ns unit
      endcase //case suffix

      return out;
   endfunction //convert_time()

   // ===============================================
   // Verification Test Library
   // ===============================================
   mby_mesh_test_lib test();

   // MBY Mesh Dut
   // ===============================================
   // ===============================================
  
   wire       w_dummy [mby_mgp_bfm_pkg::NUM_MSH_ROWS-1:0][mby_msh_pkg::NUM_MSH_ROW_PORTS-1:0];
   generate
   for (genvar gv_row=0; gv_row < mby_mgp_bfm_pkg::NUM_MSH_ROWS; gv_row++) begin
       for (genvar ports=0; ports < mby_msh_pkg::NUM_MSH_ROW_PORTS; ports++) begin
	  assign w_dummy[gv_row][ports] = 0;
       end
   end
   endgenerate
   mby_msh #(.NUM_MSH_ROWS(mby_mgp_bfm_pkg::NUM_MSH_ROWS) , .NUM_MSH_COLS(mby_mgp_bfm_pkg::NUM_MSH_COLS)) msh(
       .cclk                    (mesh_tb_if.fab_clk),
       .mclk                    (mesh_tb_if.mclk),
       .chreset                 (mesh_tb_if.chard_reset),
       .mhreset                 (mesh_tb_if.mhard_reset),
       .csreset                 (mesh_tb_if.chard_reset),
       .msreset                 (mesh_tb_if.mhard_reset),
       .i_igr_eb_wreq           (wreq_eb_if.wr_req),
       .i_igr_eb_wr_data        (wrdata_eb_if.req_data),
       .i_igr_wb_wreq           (wreq_wb_if.wr_req),
       .i_igr_wb_wr_data        (wrdata_wb_if.req_data),
       .i_egr_eb_rreq           (rreq_eb_if.rd_req),
       .i_egr_wb_rreq           (rreq_wb_if.rd_req),
//       .i_gmn_sb_wreq           (wreq_sb_if.wr_req[0]),
//       .i_gmn_sb_wr_data        (wrdata_sb_if.req_data[0]),
//       .i_gms_nb_wreq           (wreq_nb_if.wr_req[0]),
//       .i_gms_nb_wr_data        (wrdata_nb_if.req_data[0]),
//       .i_gmn_sb_rreq           (rreq_sb_if.rd_req[0]),
//       .i_gms_nb_rreq           (rreq_nb_if.rd_req[0]),
       .o_egr_wb_rrsp		(),			      
       .o_egr_wb_rd_data        (),
       .o_egr_eb_rrsp           (),
       .o_egr_eb_rd_data        (),
//       .o_gmn_nb_rrsp           (),
//       .o_gmn_nb_rd_data        (),
//       .o_gms_sb_rrsp           (),
//       .o_gms_sb_rd_data        (),
       .o_igr_eb_wr_lat_sat     (),
       .o_igr_crdt_rtn_for_eb_wreq (),
       .o_igr_mcast_crdt_rtn_for_eb_wreq (),
       .o_igr_wb_wr_lat_sat     (),
       .o_igr_crdt_rtn_for_wb_wreq (),
       .o_igr_mcast_crdt_rtn_for_wb_wreq (),
       .o_egr_eb_rd_lat_sat     (),
       .o_egr_crdt_rtn_for_eb_rreq (),
       .o_egr_mcast_crdt_rtn_for_eb_rreq (),
       .o_egr_wb_rd_lat_sat     (),
       .o_egr_crdt_rtn_for_wb_rreq (),
       .o_egr_mcast_crdt_rtn_for_wb_rreq (),
       .i_egr_crdt_rtn_for_wb_rrsp (w_dummy),
       .i_egr_mcast_crdt_rtn_for_wb_rrsp (w_dummy),
       .i_egr_crdt_rtn_for_eb_rrsp (w_dummy),
       .i_egr_mcast_crdt_rtn_for_eb_rrsp (w_dummy),
       .o_gmn_sb_wr_lat_sat (),
       .o_gmn_crdt_rtn_for_sb_wreq (),
       .o_gmn_mcast_crdt_rtn_for_sb_wreq ()
//       .o_gms_nb_wr_lat_sat (),
//       .o_gms_crdt_rtn_for_nb_wreq (),
//       .o_gms_mcast_crdt_rtn_for_nb_wreq (),
//       .o_gmn_sb_rd_lat_sat (),
//       .o_gmn_crdt_rtn_for_sb_rreq (),
//       .o_gmn_mcast_crdt_rtn_for_sb_rreq (),
//       .o_gms_nb_rd_lat_sat (),
//       .o_gms_crdt_rtn_for_nb_rreq (),
//       .o_gms_mcast_crdt_rtn_for_nb_rreq (),
//       .i_gmn_crdt_rtn_for_nb_rrsp (w_dummy[0]),
//       .i_gmn_mcast_crdt_rtn_for_nb_rrsp (w_dummy[0]),
//       .i_gms_crdt_rtn_for_sb_rrsp (w_dummy[0]),
//       .i_gms_mcast_crdt_rtn_for_sb_rrsp (w_dummy[0])		      
       );
endmodule
