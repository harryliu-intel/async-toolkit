magic
tech scmos
timestamp 969938295
<< ndiffusion >>
rect -16 142 -8 143
rect -16 138 -8 139
rect -64 123 -61 127
rect -56 123 -51 127
rect -48 123 -45 127
rect -24 105 -8 106
rect -24 97 -8 102
rect -24 93 -8 94
<< pdiffusion >>
rect 8 142 16 143
rect 8 138 16 139
rect 23 134 27 143
rect 46 140 58 141
rect 46 131 58 132
rect 23 127 27 130
rect 46 127 58 128
rect 54 122 58 127
rect 8 105 24 106
rect 8 97 24 102
rect 8 93 24 94
<< ntransistor >>
rect -16 139 -8 142
rect -61 123 -56 127
rect -51 123 -48 127
rect -24 102 -8 105
rect -24 94 -8 97
<< ptransistor >>
rect 8 139 16 142
rect 23 130 27 134
rect 46 128 58 131
rect 8 102 24 105
rect 8 94 24 97
<< polysilicon >>
rect -61 127 -56 141
rect -20 139 -16 142
rect -8 139 -4 142
rect -51 129 -33 132
rect -51 127 -48 129
rect 4 139 8 142
rect 16 139 20 142
rect 18 130 23 134
rect 27 131 29 134
rect 62 131 65 139
rect 27 130 31 131
rect 18 128 21 130
rect -61 119 -56 123
rect -51 119 -48 123
rect -28 125 21 128
rect 42 128 46 131
rect 58 128 65 131
rect -28 102 -24 105
rect -8 102 8 105
rect 24 102 28 105
rect -28 94 -24 97
rect -8 94 -4 97
rect 4 94 8 97
rect 24 94 28 97
<< ndcontact >>
rect -16 143 -8 151
rect -16 130 -8 138
rect -72 119 -64 127
rect -45 119 -37 127
rect -24 106 -8 114
rect -24 85 -8 93
<< pdcontact >>
rect 8 143 16 151
rect 22 143 30 151
rect 8 130 16 138
rect 46 132 58 140
rect 23 119 31 127
rect 46 119 54 127
rect 8 106 24 114
rect 8 85 24 93
<< psubstratepcontact >>
rect -46 136 -38 144
<< nsubstratencontact >>
rect 46 141 58 149
<< polycontact >>
rect -64 141 -56 149
rect -33 128 -25 136
rect -4 134 4 142
rect 29 131 37 139
rect 62 139 70 147
rect -36 102 -28 110
rect -4 89 4 97
<< metal1 >>
rect -64 141 -56 145
rect -45 145 -21 151
rect -45 144 -8 145
rect -46 143 -8 144
rect 21 145 58 151
rect 8 143 58 145
rect -46 137 -38 143
rect -69 136 -38 137
rect -16 136 -8 138
rect -69 131 -39 136
rect -33 132 -8 136
rect -69 127 -64 131
rect -33 128 -25 132
rect -16 130 -8 132
rect -4 127 4 142
rect 8 136 16 138
rect 29 136 37 139
rect 8 132 37 136
rect 46 132 58 143
rect 62 139 70 145
rect 8 130 16 132
rect 29 131 37 132
rect -72 119 -64 127
rect -45 123 -37 127
rect -45 121 -4 123
rect 23 123 31 127
rect 46 123 54 127
rect 4 121 54 123
rect -45 119 54 121
rect -4 114 4 119
rect -36 102 -28 109
rect -24 107 24 114
rect -24 106 -8 107
rect 8 106 24 107
rect -24 91 -8 93
rect -24 85 -21 91
rect -4 89 4 97
rect 8 91 24 93
rect 21 85 24 91
<< m2contact >>
rect -64 145 -56 151
rect -21 145 -8 151
rect 8 145 21 151
rect 62 145 70 151
rect -4 121 4 127
rect -36 109 -28 115
rect -4 97 4 103
rect -21 85 -8 91
rect 8 85 21 91
<< metal2 >>
rect -64 145 -27 151
rect 27 145 70 151
rect -6 121 6 127
rect -36 109 0 115
rect -6 97 6 103
<< m3contact >>
rect -21 145 -8 151
rect 8 145 21 151
rect -21 85 -8 91
rect 8 85 21 91
<< metal3 >>
rect -21 82 -3 154
rect 3 82 21 154
<< labels >>
rlabel m2contact -12 89 -12 89 1 GND!
rlabel metal1 -12 110 -12 110 5 x
rlabel metal1 22 89 22 89 1 Vdd!
rlabel metal2 -6 97 -6 103 3 a
rlabel metal2 6 97 6 103 7 a
rlabel metal2 0 109 0 115 7 b
rlabel space 24 85 29 114 3 ^p
rlabel space -40 84 -24 116 7 ^n
rlabel metal2 -32 112 -32 112 1 b
rlabel metal1 0 93 0 93 1 a
rlabel metal1 26 147 26 147 5 Vdd!
rlabel metal1 -68 123 -68 123 3 GND!
rlabel polysilicon -60 128 -60 128 3 _SReset!
rlabel metal1 27 122 27 122 5 x
rlabel metal1 -41 123 -41 123 3 x
rlabel metal2 -60 148 -60 148 5 _SReset!
rlabel ndcontact -12 147 -12 147 5 GND!
rlabel pdcontact 12 147 12 147 5 Vdd!
rlabel metal1 11 110 11 110 5 x
rlabel metal2 -6 121 -6 127 3 x
rlabel metal2 6 121 6 127 7 x
rlabel metal1 0 138 0 138 1 x
rlabel metal1 -42 140 -42 140 1 GND!
rlabel metal1 50 136 50 136 6 Vdd!
rlabel polysilicon 59 130 59 130 7 _PReset!
rlabel metal2 66 148 66 148 5 _PReset!
rlabel metal1 52 143 52 143 1 Vdd!
<< end >>
