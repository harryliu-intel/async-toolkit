magic
tech scmos
timestamp 965070645
<< ndiffusion >>
rect 26 5 34 6
rect 26 1 34 2
rect 26 -8 34 -7
rect 26 -12 34 -11
rect 26 -21 34 -20
rect 26 -25 34 -24
rect 26 -34 34 -33
rect 26 -38 34 -37
rect 26 -47 34 -46
rect 26 -51 34 -50
rect 26 -60 34 -59
rect 26 -64 34 -63
<< pdiffusion >>
rect 50 -5 58 -4
rect 50 -13 58 -8
rect 50 -21 58 -16
rect 50 -25 58 -24
rect 50 -34 58 -33
rect 50 -42 58 -37
rect 50 -50 58 -45
rect 50 -54 58 -53
<< ntransistor >>
rect 26 2 34 5
rect 26 -11 34 -8
rect 26 -24 34 -21
rect 26 -37 34 -34
rect 26 -50 34 -47
rect 26 -63 34 -60
<< ptransistor >>
rect 50 -8 58 -5
rect 50 -16 58 -13
rect 50 -24 58 -21
rect 50 -37 58 -34
rect 50 -45 58 -42
rect 50 -53 58 -50
<< polysilicon >>
rect 22 2 26 5
rect 34 2 48 5
rect 45 -5 48 2
rect 45 -8 50 -5
rect 58 -8 62 -5
rect 22 -11 26 -8
rect 34 -11 39 -8
rect 36 -13 39 -11
rect 36 -16 50 -13
rect 58 -16 62 -13
rect 22 -24 26 -21
rect 34 -24 50 -21
rect 58 -24 62 -21
rect 22 -37 26 -34
rect 34 -37 50 -34
rect 58 -37 62 -34
rect 36 -45 50 -42
rect 58 -45 62 -42
rect 36 -47 39 -45
rect 22 -50 26 -47
rect 34 -50 39 -47
rect 45 -53 50 -50
rect 58 -53 62 -50
rect 45 -60 48 -53
rect 22 -63 26 -60
rect 34 -63 48 -60
<< ndcontact >>
rect 26 6 34 14
rect 26 -7 34 1
rect 26 -20 34 -12
rect 26 -33 34 -25
rect 26 -46 34 -38
rect 26 -59 34 -51
rect 26 -72 34 -64
<< pdcontact >>
rect 50 -4 58 4
rect 50 -33 58 -25
rect 50 -62 58 -54
<< metal1 >>
rect 26 6 46 14
rect 26 -7 34 1
rect 38 -12 46 6
rect 50 -4 58 4
rect 26 -20 46 -12
rect 38 -25 46 -20
rect 26 -33 34 -25
rect 38 -33 58 -25
rect 38 -38 46 -33
rect 26 -46 46 -38
rect 26 -59 34 -51
rect 38 -64 46 -46
rect 50 -62 58 -54
rect 26 -72 46 -64
<< labels >>
rlabel metal1 30 -16 30 -16 1 x
rlabel polysilicon 59 -23 59 -23 7 a
rlabel polysilicon 59 -15 59 -15 7 b
rlabel polysilicon 25 -10 25 -10 1 b
rlabel polysilicon 25 -23 25 -23 1 a
rlabel polysilicon 59 -7 59 -7 7 c
rlabel metal1 30 10 30 10 5 x
rlabel polysilicon 25 3 25 3 1 c
rlabel metal1 54 -29 54 -29 5 x
rlabel metal1 30 -42 30 -42 5 x
rlabel metal1 30 -68 30 -68 1 x
rlabel polysilicon 59 -36 59 -36 7 c
rlabel polysilicon 59 -44 59 -44 7 b
rlabel polysilicon 59 -52 59 -52 7 a
rlabel polysilicon 25 -49 25 -49 1 b
rlabel polysilicon 25 -62 25 -62 1 a
rlabel polysilicon 25 -36 25 -36 1 c
rlabel metal1 54 -58 54 -58 1 Vdd!
rlabel metal1 54 0 54 0 1 Vdd!
rlabel metal1 30 -3 30 -3 1 GND!
rlabel metal1 30 -29 30 -29 1 GND!
rlabel metal1 30 -55 30 -55 1 GND!
rlabel space 21 -72 26 14 7 ^n
rlabel space 58 -62 63 4 3 ^p
<< end >>
