module dpb_tb;
endmodule
