///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_mapper_map.sv                                      
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_mapper_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_FF
`define RTLGEN_MBY_PPE_MAPPER_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_FF

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF
`define RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_MAPPER_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_FF_RSTD


module rtlgen_mby_ppe_mapper_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_mapper_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_MAPPER_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_MAPPER_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_MAPPER_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_MAPPER_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_MAPPER_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_PH2_FF
`define RTLGEN_MBY_PPE_MAPPER_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_MAPPER_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_MAPPER_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_LATCH
`define RTLGEN_MBY_PPE_MAPPER_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_MAPPER_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_MAPPER_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_mapper_map ( //lintra s-2096
    // Clocks


    // Resets



    // Register Inputs
    handcode_reg_rdata_MAP_DOMAIN_ACTION0,
    handcode_reg_rdata_MAP_DOMAIN_ACTION1,
    handcode_reg_rdata_MAP_DOMAIN_POL_CFG,
    handcode_reg_rdata_MAP_DOMAIN_PROFILE,
    handcode_reg_rdata_MAP_DOMAIN_TCAM,
    handcode_reg_rdata_MAP_DSCP_TC,
    handcode_reg_rdata_MAP_EXP_TC,
    handcode_reg_rdata_MAP_IP_CFG,
    handcode_reg_rdata_MAP_IP_HI,
    handcode_reg_rdata_MAP_IP_LO,
    handcode_reg_rdata_MAP_L4_DST,
    handcode_reg_rdata_MAP_L4_SRC,
    handcode_reg_rdata_MAP_MAC,
    handcode_reg_rdata_MAP_PORT,
    handcode_reg_rdata_MAP_PORT_CFG,
    handcode_reg_rdata_MAP_PORT_DEFAULT,
    handcode_reg_rdata_MAP_PROFILE_ACTION,
    handcode_reg_rdata_MAP_PROFILE_KEY0,
    handcode_reg_rdata_MAP_PROFILE_KEY1,
    handcode_reg_rdata_MAP_PROFILE_KEY_INVERT0,
    handcode_reg_rdata_MAP_PROFILE_KEY_INVERT1,
    handcode_reg_rdata_MAP_PROT,
    handcode_reg_rdata_MAP_REWRITE,
    handcode_reg_rdata_MAP_VPRI,
    handcode_reg_rdata_MAP_VPRI_TC,

    handcode_rvalid_MAP_DOMAIN_ACTION0,
    handcode_rvalid_MAP_DOMAIN_ACTION1,
    handcode_rvalid_MAP_DOMAIN_POL_CFG,
    handcode_rvalid_MAP_DOMAIN_PROFILE,
    handcode_rvalid_MAP_DOMAIN_TCAM,
    handcode_rvalid_MAP_DSCP_TC,
    handcode_rvalid_MAP_EXP_TC,
    handcode_rvalid_MAP_IP_CFG,
    handcode_rvalid_MAP_IP_HI,
    handcode_rvalid_MAP_IP_LO,
    handcode_rvalid_MAP_L4_DST,
    handcode_rvalid_MAP_L4_SRC,
    handcode_rvalid_MAP_MAC,
    handcode_rvalid_MAP_PORT,
    handcode_rvalid_MAP_PORT_CFG,
    handcode_rvalid_MAP_PORT_DEFAULT,
    handcode_rvalid_MAP_PROFILE_ACTION,
    handcode_rvalid_MAP_PROFILE_KEY0,
    handcode_rvalid_MAP_PROFILE_KEY1,
    handcode_rvalid_MAP_PROFILE_KEY_INVERT0,
    handcode_rvalid_MAP_PROFILE_KEY_INVERT1,
    handcode_rvalid_MAP_PROT,
    handcode_rvalid_MAP_REWRITE,
    handcode_rvalid_MAP_VPRI,
    handcode_rvalid_MAP_VPRI_TC,

    handcode_wvalid_MAP_DOMAIN_ACTION0,
    handcode_wvalid_MAP_DOMAIN_ACTION1,
    handcode_wvalid_MAP_DOMAIN_POL_CFG,
    handcode_wvalid_MAP_DOMAIN_PROFILE,
    handcode_wvalid_MAP_DOMAIN_TCAM,
    handcode_wvalid_MAP_DSCP_TC,
    handcode_wvalid_MAP_EXP_TC,
    handcode_wvalid_MAP_IP_CFG,
    handcode_wvalid_MAP_IP_HI,
    handcode_wvalid_MAP_IP_LO,
    handcode_wvalid_MAP_L4_DST,
    handcode_wvalid_MAP_L4_SRC,
    handcode_wvalid_MAP_MAC,
    handcode_wvalid_MAP_PORT,
    handcode_wvalid_MAP_PORT_CFG,
    handcode_wvalid_MAP_PORT_DEFAULT,
    handcode_wvalid_MAP_PROFILE_ACTION,
    handcode_wvalid_MAP_PROFILE_KEY0,
    handcode_wvalid_MAP_PROFILE_KEY1,
    handcode_wvalid_MAP_PROFILE_KEY_INVERT0,
    handcode_wvalid_MAP_PROFILE_KEY_INVERT1,
    handcode_wvalid_MAP_PROT,
    handcode_wvalid_MAP_REWRITE,
    handcode_wvalid_MAP_VPRI,
    handcode_wvalid_MAP_VPRI_TC,

    handcode_error_MAP_DOMAIN_ACTION0,
    handcode_error_MAP_DOMAIN_ACTION1,
    handcode_error_MAP_DOMAIN_POL_CFG,
    handcode_error_MAP_DOMAIN_PROFILE,
    handcode_error_MAP_DOMAIN_TCAM,
    handcode_error_MAP_DSCP_TC,
    handcode_error_MAP_EXP_TC,
    handcode_error_MAP_IP_CFG,
    handcode_error_MAP_IP_HI,
    handcode_error_MAP_IP_LO,
    handcode_error_MAP_L4_DST,
    handcode_error_MAP_L4_SRC,
    handcode_error_MAP_MAC,
    handcode_error_MAP_PORT,
    handcode_error_MAP_PORT_CFG,
    handcode_error_MAP_PORT_DEFAULT,
    handcode_error_MAP_PROFILE_ACTION,
    handcode_error_MAP_PROFILE_KEY0,
    handcode_error_MAP_PROFILE_KEY1,
    handcode_error_MAP_PROFILE_KEY_INVERT0,
    handcode_error_MAP_PROFILE_KEY_INVERT1,
    handcode_error_MAP_PROT,
    handcode_error_MAP_REWRITE,
    handcode_error_MAP_VPRI,
    handcode_error_MAP_VPRI_TC,


    // Register Outputs

    // Register signals for HandCoded registers
    handcode_reg_wdata_MAP_DOMAIN_ACTION0,
    handcode_reg_wdata_MAP_DOMAIN_ACTION1,
    handcode_reg_wdata_MAP_DOMAIN_POL_CFG,
    handcode_reg_wdata_MAP_DOMAIN_PROFILE,
    handcode_reg_wdata_MAP_DOMAIN_TCAM,
    handcode_reg_wdata_MAP_DSCP_TC,
    handcode_reg_wdata_MAP_EXP_TC,
    handcode_reg_wdata_MAP_IP_CFG,
    handcode_reg_wdata_MAP_IP_HI,
    handcode_reg_wdata_MAP_IP_LO,
    handcode_reg_wdata_MAP_L4_DST,
    handcode_reg_wdata_MAP_L4_SRC,
    handcode_reg_wdata_MAP_MAC,
    handcode_reg_wdata_MAP_PORT,
    handcode_reg_wdata_MAP_PORT_CFG,
    handcode_reg_wdata_MAP_PORT_DEFAULT,
    handcode_reg_wdata_MAP_PROFILE_ACTION,
    handcode_reg_wdata_MAP_PROFILE_KEY0,
    handcode_reg_wdata_MAP_PROFILE_KEY1,
    handcode_reg_wdata_MAP_PROFILE_KEY_INVERT0,
    handcode_reg_wdata_MAP_PROFILE_KEY_INVERT1,
    handcode_reg_wdata_MAP_PROT,
    handcode_reg_wdata_MAP_REWRITE,
    handcode_reg_wdata_MAP_VPRI,
    handcode_reg_wdata_MAP_VPRI_TC,

    we_MAP_DOMAIN_ACTION0,
    we_MAP_DOMAIN_ACTION1,
    we_MAP_DOMAIN_POL_CFG,
    we_MAP_DOMAIN_PROFILE,
    we_MAP_DOMAIN_TCAM,
    we_MAP_DSCP_TC,
    we_MAP_EXP_TC,
    we_MAP_IP_CFG,
    we_MAP_IP_HI,
    we_MAP_IP_LO,
    we_MAP_L4_DST,
    we_MAP_L4_SRC,
    we_MAP_MAC,
    we_MAP_PORT,
    we_MAP_PORT_CFG,
    we_MAP_PORT_DEFAULT,
    we_MAP_PROFILE_ACTION,
    we_MAP_PROFILE_KEY0,
    we_MAP_PROFILE_KEY1,
    we_MAP_PROFILE_KEY_INVERT0,
    we_MAP_PROFILE_KEY_INVERT1,
    we_MAP_PROT,
    we_MAP_REWRITE,
    we_MAP_VPRI,
    we_MAP_VPRI_TC,

    re_MAP_DOMAIN_ACTION0,
    re_MAP_DOMAIN_ACTION1,
    re_MAP_DOMAIN_POL_CFG,
    re_MAP_DOMAIN_PROFILE,
    re_MAP_DOMAIN_TCAM,
    re_MAP_DSCP_TC,
    re_MAP_EXP_TC,
    re_MAP_IP_CFG,
    re_MAP_IP_HI,
    re_MAP_IP_LO,
    re_MAP_L4_DST,
    re_MAP_L4_SRC,
    re_MAP_MAC,
    re_MAP_PORT,
    re_MAP_PORT_CFG,
    re_MAP_PORT_DEFAULT,
    re_MAP_PROFILE_ACTION,
    re_MAP_PROFILE_KEY0,
    re_MAP_PROFILE_KEY1,
    re_MAP_PROFILE_KEY_INVERT0,
    re_MAP_PROFILE_KEY_INVERT1,
    re_MAP_PROT,
    re_MAP_REWRITE,
    re_MAP_VPRI,
    re_MAP_VPRI_TC,




    // Config Access
    req,
    ack
    

);

import mby_ppe_mapper_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:0] MBY_PPE_MAPPER_MAP_OFFSET = {MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] MAPPER_SB_BAR = 3'b0;
parameter [7:0] MAPPER_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;

    // Clocks


    // Resets



    // Register Inputs
input MAP_DOMAIN_ACTION0_t  handcode_reg_rdata_MAP_DOMAIN_ACTION0;
input MAP_DOMAIN_ACTION1_t  handcode_reg_rdata_MAP_DOMAIN_ACTION1;
input MAP_DOMAIN_POL_CFG_t  handcode_reg_rdata_MAP_DOMAIN_POL_CFG;
input MAP_DOMAIN_PROFILE_t  handcode_reg_rdata_MAP_DOMAIN_PROFILE;
input MAP_DOMAIN_TCAM_t  handcode_reg_rdata_MAP_DOMAIN_TCAM;
input MAP_DSCP_TC_t  handcode_reg_rdata_MAP_DSCP_TC;
input MAP_EXP_TC_t  handcode_reg_rdata_MAP_EXP_TC;
input MAP_IP_CFG_t  handcode_reg_rdata_MAP_IP_CFG;
input MAP_IP_HI_t  handcode_reg_rdata_MAP_IP_HI;
input MAP_IP_LO_t  handcode_reg_rdata_MAP_IP_LO;
input MAP_L4_DST_t  handcode_reg_rdata_MAP_L4_DST;
input MAP_L4_SRC_t  handcode_reg_rdata_MAP_L4_SRC;
input MAP_MAC_t  handcode_reg_rdata_MAP_MAC;
input MAP_PORT_t  handcode_reg_rdata_MAP_PORT;
input MAP_PORT_CFG_t  handcode_reg_rdata_MAP_PORT_CFG;
input MAP_PORT_DEFAULT_t  handcode_reg_rdata_MAP_PORT_DEFAULT;
input MAP_PROFILE_ACTION_t  handcode_reg_rdata_MAP_PROFILE_ACTION;
input MAP_PROFILE_KEY0_t  handcode_reg_rdata_MAP_PROFILE_KEY0;
input MAP_PROFILE_KEY1_t  handcode_reg_rdata_MAP_PROFILE_KEY1;
input MAP_PROFILE_KEY_INVERT0_t  handcode_reg_rdata_MAP_PROFILE_KEY_INVERT0;
input MAP_PROFILE_KEY_INVERT1_t  handcode_reg_rdata_MAP_PROFILE_KEY_INVERT1;
input MAP_PROT_t  handcode_reg_rdata_MAP_PROT;
input MAP_REWRITE_t  handcode_reg_rdata_MAP_REWRITE;
input MAP_VPRI_t  handcode_reg_rdata_MAP_VPRI;
input MAP_VPRI_TC_t  handcode_reg_rdata_MAP_VPRI_TC;

input handcode_rvalid_MAP_DOMAIN_ACTION0_t  handcode_rvalid_MAP_DOMAIN_ACTION0;
input handcode_rvalid_MAP_DOMAIN_ACTION1_t  handcode_rvalid_MAP_DOMAIN_ACTION1;
input handcode_rvalid_MAP_DOMAIN_POL_CFG_t  handcode_rvalid_MAP_DOMAIN_POL_CFG;
input handcode_rvalid_MAP_DOMAIN_PROFILE_t  handcode_rvalid_MAP_DOMAIN_PROFILE;
input handcode_rvalid_MAP_DOMAIN_TCAM_t  handcode_rvalid_MAP_DOMAIN_TCAM;
input handcode_rvalid_MAP_DSCP_TC_t  handcode_rvalid_MAP_DSCP_TC;
input handcode_rvalid_MAP_EXP_TC_t  handcode_rvalid_MAP_EXP_TC;
input handcode_rvalid_MAP_IP_CFG_t  handcode_rvalid_MAP_IP_CFG;
input handcode_rvalid_MAP_IP_HI_t  handcode_rvalid_MAP_IP_HI;
input handcode_rvalid_MAP_IP_LO_t  handcode_rvalid_MAP_IP_LO;
input handcode_rvalid_MAP_L4_DST_t  handcode_rvalid_MAP_L4_DST;
input handcode_rvalid_MAP_L4_SRC_t  handcode_rvalid_MAP_L4_SRC;
input handcode_rvalid_MAP_MAC_t  handcode_rvalid_MAP_MAC;
input handcode_rvalid_MAP_PORT_t  handcode_rvalid_MAP_PORT;
input handcode_rvalid_MAP_PORT_CFG_t  handcode_rvalid_MAP_PORT_CFG;
input handcode_rvalid_MAP_PORT_DEFAULT_t  handcode_rvalid_MAP_PORT_DEFAULT;
input handcode_rvalid_MAP_PROFILE_ACTION_t  handcode_rvalid_MAP_PROFILE_ACTION;
input handcode_rvalid_MAP_PROFILE_KEY0_t  handcode_rvalid_MAP_PROFILE_KEY0;
input handcode_rvalid_MAP_PROFILE_KEY1_t  handcode_rvalid_MAP_PROFILE_KEY1;
input handcode_rvalid_MAP_PROFILE_KEY_INVERT0_t  handcode_rvalid_MAP_PROFILE_KEY_INVERT0;
input handcode_rvalid_MAP_PROFILE_KEY_INVERT1_t  handcode_rvalid_MAP_PROFILE_KEY_INVERT1;
input handcode_rvalid_MAP_PROT_t  handcode_rvalid_MAP_PROT;
input handcode_rvalid_MAP_REWRITE_t  handcode_rvalid_MAP_REWRITE;
input handcode_rvalid_MAP_VPRI_t  handcode_rvalid_MAP_VPRI;
input handcode_rvalid_MAP_VPRI_TC_t  handcode_rvalid_MAP_VPRI_TC;

input handcode_wvalid_MAP_DOMAIN_ACTION0_t  handcode_wvalid_MAP_DOMAIN_ACTION0;
input handcode_wvalid_MAP_DOMAIN_ACTION1_t  handcode_wvalid_MAP_DOMAIN_ACTION1;
input handcode_wvalid_MAP_DOMAIN_POL_CFG_t  handcode_wvalid_MAP_DOMAIN_POL_CFG;
input handcode_wvalid_MAP_DOMAIN_PROFILE_t  handcode_wvalid_MAP_DOMAIN_PROFILE;
input handcode_wvalid_MAP_DOMAIN_TCAM_t  handcode_wvalid_MAP_DOMAIN_TCAM;
input handcode_wvalid_MAP_DSCP_TC_t  handcode_wvalid_MAP_DSCP_TC;
input handcode_wvalid_MAP_EXP_TC_t  handcode_wvalid_MAP_EXP_TC;
input handcode_wvalid_MAP_IP_CFG_t  handcode_wvalid_MAP_IP_CFG;
input handcode_wvalid_MAP_IP_HI_t  handcode_wvalid_MAP_IP_HI;
input handcode_wvalid_MAP_IP_LO_t  handcode_wvalid_MAP_IP_LO;
input handcode_wvalid_MAP_L4_DST_t  handcode_wvalid_MAP_L4_DST;
input handcode_wvalid_MAP_L4_SRC_t  handcode_wvalid_MAP_L4_SRC;
input handcode_wvalid_MAP_MAC_t  handcode_wvalid_MAP_MAC;
input handcode_wvalid_MAP_PORT_t  handcode_wvalid_MAP_PORT;
input handcode_wvalid_MAP_PORT_CFG_t  handcode_wvalid_MAP_PORT_CFG;
input handcode_wvalid_MAP_PORT_DEFAULT_t  handcode_wvalid_MAP_PORT_DEFAULT;
input handcode_wvalid_MAP_PROFILE_ACTION_t  handcode_wvalid_MAP_PROFILE_ACTION;
input handcode_wvalid_MAP_PROFILE_KEY0_t  handcode_wvalid_MAP_PROFILE_KEY0;
input handcode_wvalid_MAP_PROFILE_KEY1_t  handcode_wvalid_MAP_PROFILE_KEY1;
input handcode_wvalid_MAP_PROFILE_KEY_INVERT0_t  handcode_wvalid_MAP_PROFILE_KEY_INVERT0;
input handcode_wvalid_MAP_PROFILE_KEY_INVERT1_t  handcode_wvalid_MAP_PROFILE_KEY_INVERT1;
input handcode_wvalid_MAP_PROT_t  handcode_wvalid_MAP_PROT;
input handcode_wvalid_MAP_REWRITE_t  handcode_wvalid_MAP_REWRITE;
input handcode_wvalid_MAP_VPRI_t  handcode_wvalid_MAP_VPRI;
input handcode_wvalid_MAP_VPRI_TC_t  handcode_wvalid_MAP_VPRI_TC;

input handcode_error_MAP_DOMAIN_ACTION0_t  handcode_error_MAP_DOMAIN_ACTION0;
input handcode_error_MAP_DOMAIN_ACTION1_t  handcode_error_MAP_DOMAIN_ACTION1;
input handcode_error_MAP_DOMAIN_POL_CFG_t  handcode_error_MAP_DOMAIN_POL_CFG;
input handcode_error_MAP_DOMAIN_PROFILE_t  handcode_error_MAP_DOMAIN_PROFILE;
input handcode_error_MAP_DOMAIN_TCAM_t  handcode_error_MAP_DOMAIN_TCAM;
input handcode_error_MAP_DSCP_TC_t  handcode_error_MAP_DSCP_TC;
input handcode_error_MAP_EXP_TC_t  handcode_error_MAP_EXP_TC;
input handcode_error_MAP_IP_CFG_t  handcode_error_MAP_IP_CFG;
input handcode_error_MAP_IP_HI_t  handcode_error_MAP_IP_HI;
input handcode_error_MAP_IP_LO_t  handcode_error_MAP_IP_LO;
input handcode_error_MAP_L4_DST_t  handcode_error_MAP_L4_DST;
input handcode_error_MAP_L4_SRC_t  handcode_error_MAP_L4_SRC;
input handcode_error_MAP_MAC_t  handcode_error_MAP_MAC;
input handcode_error_MAP_PORT_t  handcode_error_MAP_PORT;
input handcode_error_MAP_PORT_CFG_t  handcode_error_MAP_PORT_CFG;
input handcode_error_MAP_PORT_DEFAULT_t  handcode_error_MAP_PORT_DEFAULT;
input handcode_error_MAP_PROFILE_ACTION_t  handcode_error_MAP_PROFILE_ACTION;
input handcode_error_MAP_PROFILE_KEY0_t  handcode_error_MAP_PROFILE_KEY0;
input handcode_error_MAP_PROFILE_KEY1_t  handcode_error_MAP_PROFILE_KEY1;
input handcode_error_MAP_PROFILE_KEY_INVERT0_t  handcode_error_MAP_PROFILE_KEY_INVERT0;
input handcode_error_MAP_PROFILE_KEY_INVERT1_t  handcode_error_MAP_PROFILE_KEY_INVERT1;
input handcode_error_MAP_PROT_t  handcode_error_MAP_PROT;
input handcode_error_MAP_REWRITE_t  handcode_error_MAP_REWRITE;
input handcode_error_MAP_VPRI_t  handcode_error_MAP_VPRI;
input handcode_error_MAP_VPRI_TC_t  handcode_error_MAP_VPRI_TC;


    // Register Outputs

    // Register signals for HandCoded registers
output MAP_DOMAIN_ACTION0_t  handcode_reg_wdata_MAP_DOMAIN_ACTION0;
output MAP_DOMAIN_ACTION1_t  handcode_reg_wdata_MAP_DOMAIN_ACTION1;
output MAP_DOMAIN_POL_CFG_t  handcode_reg_wdata_MAP_DOMAIN_POL_CFG;
output MAP_DOMAIN_PROFILE_t  handcode_reg_wdata_MAP_DOMAIN_PROFILE;
output MAP_DOMAIN_TCAM_t  handcode_reg_wdata_MAP_DOMAIN_TCAM;
output MAP_DSCP_TC_t  handcode_reg_wdata_MAP_DSCP_TC;
output MAP_EXP_TC_t  handcode_reg_wdata_MAP_EXP_TC;
output MAP_IP_CFG_t  handcode_reg_wdata_MAP_IP_CFG;
output MAP_IP_HI_t  handcode_reg_wdata_MAP_IP_HI;
output MAP_IP_LO_t  handcode_reg_wdata_MAP_IP_LO;
output MAP_L4_DST_t  handcode_reg_wdata_MAP_L4_DST;
output MAP_L4_SRC_t  handcode_reg_wdata_MAP_L4_SRC;
output MAP_MAC_t  handcode_reg_wdata_MAP_MAC;
output MAP_PORT_t  handcode_reg_wdata_MAP_PORT;
output MAP_PORT_CFG_t  handcode_reg_wdata_MAP_PORT_CFG;
output MAP_PORT_DEFAULT_t  handcode_reg_wdata_MAP_PORT_DEFAULT;
output MAP_PROFILE_ACTION_t  handcode_reg_wdata_MAP_PROFILE_ACTION;
output MAP_PROFILE_KEY0_t  handcode_reg_wdata_MAP_PROFILE_KEY0;
output MAP_PROFILE_KEY1_t  handcode_reg_wdata_MAP_PROFILE_KEY1;
output MAP_PROFILE_KEY_INVERT0_t  handcode_reg_wdata_MAP_PROFILE_KEY_INVERT0;
output MAP_PROFILE_KEY_INVERT1_t  handcode_reg_wdata_MAP_PROFILE_KEY_INVERT1;
output MAP_PROT_t  handcode_reg_wdata_MAP_PROT;
output MAP_REWRITE_t  handcode_reg_wdata_MAP_REWRITE;
output MAP_VPRI_t  handcode_reg_wdata_MAP_VPRI;
output MAP_VPRI_TC_t  handcode_reg_wdata_MAP_VPRI_TC;

output we_MAP_DOMAIN_ACTION0_t  we_MAP_DOMAIN_ACTION0;
output we_MAP_DOMAIN_ACTION1_t  we_MAP_DOMAIN_ACTION1;
output we_MAP_DOMAIN_POL_CFG_t  we_MAP_DOMAIN_POL_CFG;
output we_MAP_DOMAIN_PROFILE_t  we_MAP_DOMAIN_PROFILE;
output we_MAP_DOMAIN_TCAM_t  we_MAP_DOMAIN_TCAM;
output we_MAP_DSCP_TC_t  we_MAP_DSCP_TC;
output we_MAP_EXP_TC_t  we_MAP_EXP_TC;
output we_MAP_IP_CFG_t  we_MAP_IP_CFG;
output we_MAP_IP_HI_t  we_MAP_IP_HI;
output we_MAP_IP_LO_t  we_MAP_IP_LO;
output we_MAP_L4_DST_t  we_MAP_L4_DST;
output we_MAP_L4_SRC_t  we_MAP_L4_SRC;
output we_MAP_MAC_t  we_MAP_MAC;
output we_MAP_PORT_t  we_MAP_PORT;
output we_MAP_PORT_CFG_t  we_MAP_PORT_CFG;
output we_MAP_PORT_DEFAULT_t  we_MAP_PORT_DEFAULT;
output we_MAP_PROFILE_ACTION_t  we_MAP_PROFILE_ACTION;
output we_MAP_PROFILE_KEY0_t  we_MAP_PROFILE_KEY0;
output we_MAP_PROFILE_KEY1_t  we_MAP_PROFILE_KEY1;
output we_MAP_PROFILE_KEY_INVERT0_t  we_MAP_PROFILE_KEY_INVERT0;
output we_MAP_PROFILE_KEY_INVERT1_t  we_MAP_PROFILE_KEY_INVERT1;
output we_MAP_PROT_t  we_MAP_PROT;
output we_MAP_REWRITE_t  we_MAP_REWRITE;
output we_MAP_VPRI_t  we_MAP_VPRI;
output we_MAP_VPRI_TC_t  we_MAP_VPRI_TC;

output re_MAP_DOMAIN_ACTION0_t  re_MAP_DOMAIN_ACTION0;
output re_MAP_DOMAIN_ACTION1_t  re_MAP_DOMAIN_ACTION1;
output re_MAP_DOMAIN_POL_CFG_t  re_MAP_DOMAIN_POL_CFG;
output re_MAP_DOMAIN_PROFILE_t  re_MAP_DOMAIN_PROFILE;
output re_MAP_DOMAIN_TCAM_t  re_MAP_DOMAIN_TCAM;
output re_MAP_DSCP_TC_t  re_MAP_DSCP_TC;
output re_MAP_EXP_TC_t  re_MAP_EXP_TC;
output re_MAP_IP_CFG_t  re_MAP_IP_CFG;
output re_MAP_IP_HI_t  re_MAP_IP_HI;
output re_MAP_IP_LO_t  re_MAP_IP_LO;
output re_MAP_L4_DST_t  re_MAP_L4_DST;
output re_MAP_L4_SRC_t  re_MAP_L4_SRC;
output re_MAP_MAC_t  re_MAP_MAC;
output re_MAP_PORT_t  re_MAP_PORT;
output re_MAP_PORT_CFG_t  re_MAP_PORT_CFG;
output re_MAP_PORT_DEFAULT_t  re_MAP_PORT_DEFAULT;
output re_MAP_PROFILE_ACTION_t  re_MAP_PROFILE_ACTION;
output re_MAP_PROFILE_KEY0_t  re_MAP_PROFILE_KEY0;
output re_MAP_PROFILE_KEY1_t  re_MAP_PROFILE_KEY1;
output re_MAP_PROFILE_KEY_INVERT0_t  re_MAP_PROFILE_KEY_INVERT0;
output re_MAP_PROFILE_KEY_INVERT1_t  re_MAP_PROFILE_KEY_INVERT1;
output re_MAP_PROT_t  re_MAP_PROT;
output re_MAP_REWRITE_t  re_MAP_REWRITE;
output re_MAP_VPRI_t  re_MAP_VPRI;
output re_MAP_VPRI_TC_t  re_MAP_VPRI_TC;




    // Config Access
input mby_ppe_mapper_map_cr_req_t  req;
output mby_ppe_mapper_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_mapper_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_MAPPER_MAP_MEM;
assign case_req_addr_MBY_PPE_MAPPER_MAP_MEM = req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_mapper;
always_comb begin : sb_fid_cond_mapper_BLOCK
    unique casez (req_fid) 
		MAPPER_SB_FID: sb_fid_cond_mapper = 1;
		default: sb_fid_cond_mapper = 0;
    endcase 
end


logic sb_bar_cond_mapper;
always_comb begin : sb_bar_cond_mapper_BLOCK
    unique casez (req_bar) 
		MAPPER_SB_BAR: sb_bar_cond_mapper = 1;
		default: sb_bar_cond_mapper = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// MAP_PORT_CFG using HANDCODED_REG template.
logic addr_decode_MAP_PORT_CFG;
logic write_req_MAP_PORT_CFG;
logic read_req_MAP_PORT_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'b0???,1'b?},
      {44'h8,1'b?}:
          addr_decode_MAP_PORT_CFG = req.valid;
      default: 
         addr_decode_MAP_PORT_CFG = 1'b0; 
   endcase
end

always_comb write_req_MAP_PORT_CFG = f_IsMEMWr(req_opcode) && addr_decode_MAP_PORT_CFG ;
always_comb read_req_MAP_PORT_CFG  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PORT_CFG ;

always_comb we_MAP_PORT_CFG = {8{write_req_MAP_PORT_CFG}} & be;
always_comb re_MAP_PORT_CFG = {8{read_req_MAP_PORT_CFG}} & be;
always_comb handcode_reg_wdata_MAP_PORT_CFG = write_data;


// ----------------------------------------------------------------------
// MAP_PORT_DEFAULT using HANDCODED_REG template.
logic addr_decode_MAP_PORT_DEFAULT;
logic write_req_MAP_PORT_DEFAULT;
logic read_req_MAP_PORT_DEFAULT;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'b1???0?,1'b?},
      {44'b1???10,1'b?},
      {44'b10???0?,1'b?},
      {44'b10???10,1'b?},
      {40'h6,4'b0?0?,1'b?},
      {40'h6,4'b0?10,1'b?}:
          addr_decode_MAP_PORT_DEFAULT = req.valid;
      default: 
         addr_decode_MAP_PORT_DEFAULT = 1'b0; 
   endcase
end

always_comb write_req_MAP_PORT_DEFAULT = f_IsMEMWr(req_opcode) && addr_decode_MAP_PORT_DEFAULT ;
always_comb read_req_MAP_PORT_DEFAULT  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PORT_DEFAULT ;

always_comb we_MAP_PORT_DEFAULT = {8{write_req_MAP_PORT_DEFAULT}} & be;
always_comb re_MAP_PORT_DEFAULT = {8{read_req_MAP_PORT_DEFAULT}} & be;
always_comb handcode_reg_wdata_MAP_PORT_DEFAULT = write_data;


// ----------------------------------------------------------------------
// MAP_DOMAIN_TCAM using HANDCODED_REG template.
logic addr_decode_MAP_DOMAIN_TCAM;
logic write_req_MAP_DOMAIN_TCAM;
logic read_req_MAP_DOMAIN_TCAM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h1???,1'b0}: 
         addr_decode_MAP_DOMAIN_TCAM = req.valid;
      default: 
         addr_decode_MAP_DOMAIN_TCAM = 1'b0; 
   endcase
end

always_comb write_req_MAP_DOMAIN_TCAM = f_IsMEMWr(req_opcode) && addr_decode_MAP_DOMAIN_TCAM ;
always_comb read_req_MAP_DOMAIN_TCAM  = f_IsMEMRd(req_opcode) && addr_decode_MAP_DOMAIN_TCAM ;

always_comb we_MAP_DOMAIN_TCAM = {16{write_req_MAP_DOMAIN_TCAM}} & req.be[15:0];
always_comb re_MAP_DOMAIN_TCAM = {16{read_req_MAP_DOMAIN_TCAM}} & req.be[15:0];
always_comb handcode_reg_wdata_MAP_DOMAIN_TCAM = req.data[127:0];


// ----------------------------------------------------------------------
// MAP_DOMAIN_ACTION0 using HANDCODED_REG template.
logic addr_decode_MAP_DOMAIN_ACTION0;
logic write_req_MAP_DOMAIN_ACTION0;
logic read_req_MAP_DOMAIN_ACTION0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h2,4'b0???,8'h??,1'b?}: 
         addr_decode_MAP_DOMAIN_ACTION0 = req.valid;
      default: 
         addr_decode_MAP_DOMAIN_ACTION0 = 1'b0; 
   endcase
end

always_comb write_req_MAP_DOMAIN_ACTION0 = f_IsMEMWr(req_opcode) && addr_decode_MAP_DOMAIN_ACTION0 ;
always_comb read_req_MAP_DOMAIN_ACTION0  = f_IsMEMRd(req_opcode) && addr_decode_MAP_DOMAIN_ACTION0 ;

always_comb we_MAP_DOMAIN_ACTION0 = {8{write_req_MAP_DOMAIN_ACTION0}} & be;
always_comb re_MAP_DOMAIN_ACTION0 = {8{read_req_MAP_DOMAIN_ACTION0}} & be;
always_comb handcode_reg_wdata_MAP_DOMAIN_ACTION0 = write_data;


// ----------------------------------------------------------------------
// MAP_DOMAIN_ACTION1 using HANDCODED_REG template.
logic addr_decode_MAP_DOMAIN_ACTION1;
logic write_req_MAP_DOMAIN_ACTION1;
logic read_req_MAP_DOMAIN_ACTION1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h2,4'b1???,8'h??,1'b?}: 
         addr_decode_MAP_DOMAIN_ACTION1 = req.valid;
      default: 
         addr_decode_MAP_DOMAIN_ACTION1 = 1'b0; 
   endcase
end

always_comb write_req_MAP_DOMAIN_ACTION1 = f_IsMEMWr(req_opcode) && addr_decode_MAP_DOMAIN_ACTION1 ;
always_comb read_req_MAP_DOMAIN_ACTION1  = f_IsMEMRd(req_opcode) && addr_decode_MAP_DOMAIN_ACTION1 ;

always_comb we_MAP_DOMAIN_ACTION1 = {8{write_req_MAP_DOMAIN_ACTION1}} & be;
always_comb re_MAP_DOMAIN_ACTION1 = {8{read_req_MAP_DOMAIN_ACTION1}} & be;
always_comb handcode_reg_wdata_MAP_DOMAIN_ACTION1 = write_data;


// ----------------------------------------------------------------------
// MAP_DOMAIN_PROFILE using HANDCODED_REG template.
logic addr_decode_MAP_DOMAIN_PROFILE;
logic write_req_MAP_DOMAIN_PROFILE;
logic read_req_MAP_DOMAIN_PROFILE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h30,4'b0???,4'h?,1'b?}: 
         addr_decode_MAP_DOMAIN_PROFILE = req.valid;
      default: 
         addr_decode_MAP_DOMAIN_PROFILE = 1'b0; 
   endcase
end

always_comb write_req_MAP_DOMAIN_PROFILE = f_IsMEMWr(req_opcode) && addr_decode_MAP_DOMAIN_PROFILE ;
always_comb read_req_MAP_DOMAIN_PROFILE  = f_IsMEMRd(req_opcode) && addr_decode_MAP_DOMAIN_PROFILE ;

always_comb we_MAP_DOMAIN_PROFILE = {8{write_req_MAP_DOMAIN_PROFILE}} & be;
always_comb re_MAP_DOMAIN_PROFILE = {8{read_req_MAP_DOMAIN_PROFILE}} & be;
always_comb handcode_reg_wdata_MAP_DOMAIN_PROFILE = write_data;


// ----------------------------------------------------------------------
// MAP_PORT using HANDCODED_REG template.
logic addr_decode_MAP_PORT;
logic write_req_MAP_PORT;
logic read_req_MAP_PORT;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h310,4'b0???,1'b?},
      {44'h3108,1'b?}:
          addr_decode_MAP_PORT = req.valid;
      default: 
         addr_decode_MAP_PORT = 1'b0; 
   endcase
end

always_comb write_req_MAP_PORT = f_IsMEMWr(req_opcode) && addr_decode_MAP_PORT ;
always_comb read_req_MAP_PORT  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PORT ;

always_comb we_MAP_PORT = {8{write_req_MAP_PORT}} & be;
always_comb re_MAP_PORT = {8{read_req_MAP_PORT}} & be;
always_comb handcode_reg_wdata_MAP_PORT = write_data;


// ----------------------------------------------------------------------
// MAP_MAC using HANDCODED_REG template.
logic addr_decode_MAP_MAC;
logic write_req_MAP_MAC;
logic read_req_MAP_MAC;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h31,4'b10??,4'h?,1'b0},
      {36'h31,4'b110?,4'h?,1'b0}:
          addr_decode_MAP_MAC = req.valid;
      default: 
         addr_decode_MAP_MAC = 1'b0; 
   endcase
end

always_comb write_req_MAP_MAC = f_IsMEMWr(req_opcode) && addr_decode_MAP_MAC ;
always_comb read_req_MAP_MAC  = f_IsMEMRd(req_opcode) && addr_decode_MAP_MAC ;

always_comb we_MAP_MAC = {16{write_req_MAP_MAC}} & req.be[15:0];
always_comb re_MAP_MAC = {16{read_req_MAP_MAC}} & req.be[15:0];
always_comb handcode_reg_wdata_MAP_MAC = req.data[127:0];


// ----------------------------------------------------------------------
// MAP_IP_LO using HANDCODED_REG template.
logic addr_decode_MAP_IP_LO;
logic write_req_MAP_IP_LO;
logic read_req_MAP_IP_LO;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h320,4'b1???,1'b?}: 
         addr_decode_MAP_IP_LO = req.valid;
      default: 
         addr_decode_MAP_IP_LO = 1'b0; 
   endcase
end

always_comb write_req_MAP_IP_LO = f_IsMEMWr(req_opcode) && addr_decode_MAP_IP_LO ;
always_comb read_req_MAP_IP_LO  = f_IsMEMRd(req_opcode) && addr_decode_MAP_IP_LO ;

always_comb we_MAP_IP_LO = {8{write_req_MAP_IP_LO}} & be;
always_comb re_MAP_IP_LO = {8{read_req_MAP_IP_LO}} & be;
always_comb handcode_reg_wdata_MAP_IP_LO = write_data;


// ----------------------------------------------------------------------
// MAP_IP_HI using HANDCODED_REG template.
logic addr_decode_MAP_IP_HI;
logic write_req_MAP_IP_HI;
logic read_req_MAP_IP_HI;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h321,4'b0???,1'b?}: 
         addr_decode_MAP_IP_HI = req.valid;
      default: 
         addr_decode_MAP_IP_HI = 1'b0; 
   endcase
end

always_comb write_req_MAP_IP_HI = f_IsMEMWr(req_opcode) && addr_decode_MAP_IP_HI ;
always_comb read_req_MAP_IP_HI  = f_IsMEMRd(req_opcode) && addr_decode_MAP_IP_HI ;

always_comb we_MAP_IP_HI = {8{write_req_MAP_IP_HI}} & be;
always_comb re_MAP_IP_HI = {8{read_req_MAP_IP_HI}} & be;
always_comb handcode_reg_wdata_MAP_IP_HI = write_data;


// ----------------------------------------------------------------------
// MAP_IP_CFG using HANDCODED_REG template.
logic addr_decode_MAP_IP_CFG;
logic write_req_MAP_IP_CFG;
logic read_req_MAP_IP_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h321,4'b1???,1'b?}: 
         addr_decode_MAP_IP_CFG = req.valid;
      default: 
         addr_decode_MAP_IP_CFG = 1'b0; 
   endcase
end

always_comb write_req_MAP_IP_CFG = f_IsMEMWr(req_opcode) && addr_decode_MAP_IP_CFG ;
always_comb read_req_MAP_IP_CFG  = f_IsMEMRd(req_opcode) && addr_decode_MAP_IP_CFG ;

always_comb we_MAP_IP_CFG = {8{write_req_MAP_IP_CFG}} & be;
always_comb re_MAP_IP_CFG = {8{read_req_MAP_IP_CFG}} & be;
always_comb handcode_reg_wdata_MAP_IP_CFG = write_data;


// ----------------------------------------------------------------------
// MAP_PROT using HANDCODED_REG template.
logic addr_decode_MAP_PROT;
logic write_req_MAP_PROT;
logic read_req_MAP_PROT;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h322,4'b00??,1'b?}: 
         addr_decode_MAP_PROT = req.valid;
      default: 
         addr_decode_MAP_PROT = 1'b0; 
   endcase
end

always_comb write_req_MAP_PROT = f_IsMEMWr(req_opcode) && addr_decode_MAP_PROT ;
always_comb read_req_MAP_PROT  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PROT ;

always_comb we_MAP_PROT = {8{write_req_MAP_PROT}} & be;
always_comb re_MAP_PROT = {8{read_req_MAP_PROT}} & be;
always_comb handcode_reg_wdata_MAP_PROT = write_data;


// ----------------------------------------------------------------------
// MAP_L4_SRC using HANDCODED_REG template.
logic addr_decode_MAP_L4_SRC;
logic write_req_MAP_L4_SRC;
logic read_req_MAP_L4_SRC;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h32,4'b010?,4'h?,1'b?}: 
         addr_decode_MAP_L4_SRC = req.valid;
      default: 
         addr_decode_MAP_L4_SRC = 1'b0; 
   endcase
end

always_comb write_req_MAP_L4_SRC = f_IsMEMWr(req_opcode) && addr_decode_MAP_L4_SRC ;
always_comb read_req_MAP_L4_SRC  = f_IsMEMRd(req_opcode) && addr_decode_MAP_L4_SRC ;

always_comb we_MAP_L4_SRC = {8{write_req_MAP_L4_SRC}} & be;
always_comb re_MAP_L4_SRC = {8{read_req_MAP_L4_SRC}} & be;
always_comb handcode_reg_wdata_MAP_L4_SRC = write_data;


// ----------------------------------------------------------------------
// MAP_L4_DST using HANDCODED_REG template.
logic addr_decode_MAP_L4_DST;
logic write_req_MAP_L4_DST;
logic read_req_MAP_L4_DST;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h32,4'b011?,4'h?,1'b?}: 
         addr_decode_MAP_L4_DST = req.valid;
      default: 
         addr_decode_MAP_L4_DST = 1'b0; 
   endcase
end

always_comb write_req_MAP_L4_DST = f_IsMEMWr(req_opcode) && addr_decode_MAP_L4_DST ;
always_comb read_req_MAP_L4_DST  = f_IsMEMRd(req_opcode) && addr_decode_MAP_L4_DST ;

always_comb we_MAP_L4_DST = {8{write_req_MAP_L4_DST}} & be;
always_comb re_MAP_L4_DST = {8{read_req_MAP_L4_DST}} & be;
always_comb handcode_reg_wdata_MAP_L4_DST = write_data;


// ----------------------------------------------------------------------
// MAP_EXP_TC using HANDCODED_REG template.
logic addr_decode_MAP_EXP_TC;
logic write_req_MAP_EXP_TC;
logic read_req_MAP_EXP_TC;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h328?,1'b?}: 
         addr_decode_MAP_EXP_TC = req.valid;
      default: 
         addr_decode_MAP_EXP_TC = 1'b0; 
   endcase
end

always_comb write_req_MAP_EXP_TC = f_IsMEMWr(req_opcode) && addr_decode_MAP_EXP_TC ;
always_comb read_req_MAP_EXP_TC  = f_IsMEMRd(req_opcode) && addr_decode_MAP_EXP_TC ;

always_comb we_MAP_EXP_TC = {8{write_req_MAP_EXP_TC}} & be;
always_comb re_MAP_EXP_TC = {8{read_req_MAP_EXP_TC}} & be;
always_comb handcode_reg_wdata_MAP_EXP_TC = write_data;


// ----------------------------------------------------------------------
// MAP_DSCP_TC using HANDCODED_REG template.
logic addr_decode_MAP_DSCP_TC;
logic write_req_MAP_DSCP_TC;
logic read_req_MAP_DSCP_TC;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h3,4'b01??,8'h??,1'b?}: 
         addr_decode_MAP_DSCP_TC = req.valid;
      default: 
         addr_decode_MAP_DSCP_TC = 1'b0; 
   endcase
end

always_comb write_req_MAP_DSCP_TC = f_IsMEMWr(req_opcode) && addr_decode_MAP_DSCP_TC ;
always_comb read_req_MAP_DSCP_TC  = f_IsMEMRd(req_opcode) && addr_decode_MAP_DSCP_TC ;

always_comb we_MAP_DSCP_TC = {8{write_req_MAP_DSCP_TC}} & be;
always_comb re_MAP_DSCP_TC = {8{read_req_MAP_DSCP_TC}} & be;
always_comb handcode_reg_wdata_MAP_DSCP_TC = write_data;


// ----------------------------------------------------------------------
// MAP_VPRI_TC using HANDCODED_REG template.
logic addr_decode_MAP_VPRI_TC;
logic write_req_MAP_VPRI_TC;
logic read_req_MAP_VPRI_TC;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h380?,1'b?}: 
         addr_decode_MAP_VPRI_TC = req.valid;
      default: 
         addr_decode_MAP_VPRI_TC = 1'b0; 
   endcase
end

always_comb write_req_MAP_VPRI_TC = f_IsMEMWr(req_opcode) && addr_decode_MAP_VPRI_TC ;
always_comb read_req_MAP_VPRI_TC  = f_IsMEMRd(req_opcode) && addr_decode_MAP_VPRI_TC ;

always_comb we_MAP_VPRI_TC = {8{write_req_MAP_VPRI_TC}} & be;
always_comb re_MAP_VPRI_TC = {8{read_req_MAP_VPRI_TC}} & be;
always_comb handcode_reg_wdata_MAP_VPRI_TC = write_data;


// ----------------------------------------------------------------------
// MAP_VPRI using HANDCODED_REG template.
logic addr_decode_MAP_VPRI;
logic write_req_MAP_VPRI;
logic read_req_MAP_VPRI;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h381?,1'b?}: 
         addr_decode_MAP_VPRI = req.valid;
      default: 
         addr_decode_MAP_VPRI = 1'b0; 
   endcase
end

always_comb write_req_MAP_VPRI = f_IsMEMWr(req_opcode) && addr_decode_MAP_VPRI ;
always_comb read_req_MAP_VPRI  = f_IsMEMRd(req_opcode) && addr_decode_MAP_VPRI ;

always_comb we_MAP_VPRI = {8{write_req_MAP_VPRI}} & be;
always_comb re_MAP_VPRI = {8{read_req_MAP_VPRI}} & be;
always_comb handcode_reg_wdata_MAP_VPRI = write_data;


// ----------------------------------------------------------------------
// MAP_PROFILE_KEY0 using HANDCODED_REG template.
logic addr_decode_MAP_PROFILE_KEY0;
logic write_req_MAP_PROFILE_KEY0;
logic read_req_MAP_PROFILE_KEY0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h38,4'b010?,4'h?,1'b?},
      {44'h386?,1'b?}:
          addr_decode_MAP_PROFILE_KEY0 = req.valid;
      default: 
         addr_decode_MAP_PROFILE_KEY0 = 1'b0; 
   endcase
end

always_comb write_req_MAP_PROFILE_KEY0 = f_IsMEMWr(req_opcode) && addr_decode_MAP_PROFILE_KEY0 ;
always_comb read_req_MAP_PROFILE_KEY0  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PROFILE_KEY0 ;

always_comb we_MAP_PROFILE_KEY0 = {8{write_req_MAP_PROFILE_KEY0}} & be;
always_comb re_MAP_PROFILE_KEY0 = {8{read_req_MAP_PROFILE_KEY0}} & be;
always_comb handcode_reg_wdata_MAP_PROFILE_KEY0 = write_data;


// ----------------------------------------------------------------------
// MAP_PROFILE_KEY_INVERT0 using HANDCODED_REG template.
logic addr_decode_MAP_PROFILE_KEY_INVERT0;
logic write_req_MAP_PROFILE_KEY_INVERT0;
logic read_req_MAP_PROFILE_KEY_INVERT0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h38,4'b100?,4'h?,1'b?},
      {44'h38A?,1'b?}:
          addr_decode_MAP_PROFILE_KEY_INVERT0 = req.valid;
      default: 
         addr_decode_MAP_PROFILE_KEY_INVERT0 = 1'b0; 
   endcase
end

always_comb write_req_MAP_PROFILE_KEY_INVERT0 = f_IsMEMWr(req_opcode) && addr_decode_MAP_PROFILE_KEY_INVERT0 ;
always_comb read_req_MAP_PROFILE_KEY_INVERT0  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PROFILE_KEY_INVERT0 ;

always_comb we_MAP_PROFILE_KEY_INVERT0 = {8{write_req_MAP_PROFILE_KEY_INVERT0}} & be;
always_comb re_MAP_PROFILE_KEY_INVERT0 = {8{read_req_MAP_PROFILE_KEY_INVERT0}} & be;
always_comb handcode_reg_wdata_MAP_PROFILE_KEY_INVERT0 = write_data;


// ----------------------------------------------------------------------
// MAP_PROFILE_KEY1 using HANDCODED_REG template.
logic addr_decode_MAP_PROFILE_KEY1;
logic write_req_MAP_PROFILE_KEY1;
logic read_req_MAP_PROFILE_KEY1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h38,4'b110?,4'h?,1'b?},
      {44'h38E?,1'b?}:
          addr_decode_MAP_PROFILE_KEY1 = req.valid;
      default: 
         addr_decode_MAP_PROFILE_KEY1 = 1'b0; 
   endcase
end

always_comb write_req_MAP_PROFILE_KEY1 = f_IsMEMWr(req_opcode) && addr_decode_MAP_PROFILE_KEY1 ;
always_comb read_req_MAP_PROFILE_KEY1  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PROFILE_KEY1 ;

always_comb we_MAP_PROFILE_KEY1 = {8{write_req_MAP_PROFILE_KEY1}} & be;
always_comb re_MAP_PROFILE_KEY1 = {8{read_req_MAP_PROFILE_KEY1}} & be;
always_comb handcode_reg_wdata_MAP_PROFILE_KEY1 = write_data;


// ----------------------------------------------------------------------
// MAP_PROFILE_KEY_INVERT1 using HANDCODED_REG template.
logic addr_decode_MAP_PROFILE_KEY_INVERT1;
logic write_req_MAP_PROFILE_KEY_INVERT1;
logic read_req_MAP_PROFILE_KEY_INVERT1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h39,4'b000?,4'h?,1'b?},
      {44'h392?,1'b?}:
          addr_decode_MAP_PROFILE_KEY_INVERT1 = req.valid;
      default: 
         addr_decode_MAP_PROFILE_KEY_INVERT1 = 1'b0; 
   endcase
end

always_comb write_req_MAP_PROFILE_KEY_INVERT1 = f_IsMEMWr(req_opcode) && addr_decode_MAP_PROFILE_KEY_INVERT1 ;
always_comb read_req_MAP_PROFILE_KEY_INVERT1  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PROFILE_KEY_INVERT1 ;

always_comb we_MAP_PROFILE_KEY_INVERT1 = {8{write_req_MAP_PROFILE_KEY_INVERT1}} & be;
always_comb re_MAP_PROFILE_KEY_INVERT1 = {8{read_req_MAP_PROFILE_KEY_INVERT1}} & be;
always_comb handcode_reg_wdata_MAP_PROFILE_KEY_INVERT1 = write_data;


// ----------------------------------------------------------------------
// MAP_PROFILE_ACTION using HANDCODED_REG template.
logic addr_decode_MAP_PROFILE_ACTION;
logic write_req_MAP_PROFILE_ACTION;
logic read_req_MAP_PROFILE_ACTION;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h39,4'b010?,4'h?,1'b?},
      {44'h396?,1'b?}:
          addr_decode_MAP_PROFILE_ACTION = req.valid;
      default: 
         addr_decode_MAP_PROFILE_ACTION = 1'b0; 
   endcase
end

always_comb write_req_MAP_PROFILE_ACTION = f_IsMEMWr(req_opcode) && addr_decode_MAP_PROFILE_ACTION ;
always_comb read_req_MAP_PROFILE_ACTION  = f_IsMEMRd(req_opcode) && addr_decode_MAP_PROFILE_ACTION ;

always_comb we_MAP_PROFILE_ACTION = {8{write_req_MAP_PROFILE_ACTION}} & be;
always_comb re_MAP_PROFILE_ACTION = {8{read_req_MAP_PROFILE_ACTION}} & be;
always_comb handcode_reg_wdata_MAP_PROFILE_ACTION = write_data;


// ----------------------------------------------------------------------
// MAP_DOMAIN_POL_CFG using HANDCODED_REG template.
logic addr_decode_MAP_DOMAIN_POL_CFG;
logic write_req_MAP_DOMAIN_POL_CFG;
logic read_req_MAP_DOMAIN_POL_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h3980,1'b0}: 
         addr_decode_MAP_DOMAIN_POL_CFG = req.valid;
      default: 
         addr_decode_MAP_DOMAIN_POL_CFG = 1'b0; 
   endcase
end

always_comb write_req_MAP_DOMAIN_POL_CFG = f_IsMEMWr(req_opcode) && addr_decode_MAP_DOMAIN_POL_CFG ;
always_comb read_req_MAP_DOMAIN_POL_CFG  = f_IsMEMRd(req_opcode) && addr_decode_MAP_DOMAIN_POL_CFG ;

always_comb we_MAP_DOMAIN_POL_CFG = {8{write_req_MAP_DOMAIN_POL_CFG}} & be;
always_comb re_MAP_DOMAIN_POL_CFG = {8{read_req_MAP_DOMAIN_POL_CFG}} & be;
always_comb handcode_reg_wdata_MAP_DOMAIN_POL_CFG = write_data;


// ----------------------------------------------------------------------
// MAP_REWRITE using HANDCODED_REG template.
logic addr_decode_MAP_REWRITE;
logic write_req_MAP_REWRITE;
logic read_req_MAP_REWRITE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MAPPER_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h3A??,1'b?}: 
         addr_decode_MAP_REWRITE = req.valid;
      default: 
         addr_decode_MAP_REWRITE = 1'b0; 
   endcase
end

always_comb write_req_MAP_REWRITE = f_IsMEMWr(req_opcode) && addr_decode_MAP_REWRITE ;
always_comb read_req_MAP_REWRITE  = f_IsMEMRd(req_opcode) && addr_decode_MAP_REWRITE ;

always_comb we_MAP_REWRITE = {8{write_req_MAP_REWRITE}} & be;
always_comb re_MAP_REWRITE = {8{read_req_MAP_REWRITE}} & be;
always_comb handcode_reg_wdata_MAP_REWRITE = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_MAPPER_MAP_MEM) 
           {44'b0???,1'b?},
           {44'h8,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PORT_CFG;
                    ack.read_miss = handcode_error_MAP_PORT_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'b1???0?,1'b?},
           {44'b1???10,1'b?},
           {44'b10???0?,1'b?},
           {44'b10???10,1'b?},
           {40'h6,4'b0?0?,1'b?},
           {40'h6,4'b0?10,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PORT_DEFAULT;
                    ack.read_miss = handcode_error_MAP_PORT_DEFAULT;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h1???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_DOMAIN_TCAM;
                    ack.read_miss = handcode_error_MAP_DOMAIN_TCAM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h2,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_DOMAIN_ACTION0;
                    ack.read_miss = handcode_error_MAP_DOMAIN_ACTION0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h2,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_DOMAIN_ACTION1;
                    ack.read_miss = handcode_error_MAP_DOMAIN_ACTION1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h30,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_DOMAIN_PROFILE;
                    ack.read_miss = handcode_error_MAP_DOMAIN_PROFILE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h310,4'b0???,1'b?},
           {44'h3108,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PORT;
                    ack.read_miss = handcode_error_MAP_PORT;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h31,4'b10??,4'h?,1'b0},
           {36'h31,4'b110?,4'h?,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_MAC;
                    ack.read_miss = handcode_error_MAP_MAC;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h320,4'b1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_IP_LO;
                    ack.read_miss = handcode_error_MAP_IP_LO;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h321,4'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_IP_HI;
                    ack.read_miss = handcode_error_MAP_IP_HI;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h321,4'b1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_IP_CFG;
                    ack.read_miss = handcode_error_MAP_IP_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h322,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PROT;
                    ack.read_miss = handcode_error_MAP_PROT;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h32,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_L4_SRC;
                    ack.read_miss = handcode_error_MAP_L4_SRC;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h32,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_L4_DST;
                    ack.read_miss = handcode_error_MAP_L4_DST;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h328?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_EXP_TC;
                    ack.read_miss = handcode_error_MAP_EXP_TC;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h3,4'b01??,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_DSCP_TC;
                    ack.read_miss = handcode_error_MAP_DSCP_TC;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h380?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_VPRI_TC;
                    ack.read_miss = handcode_error_MAP_VPRI_TC;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h381?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_VPRI;
                    ack.read_miss = handcode_error_MAP_VPRI;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h38,4'b010?,4'h?,1'b?},
           {44'h386?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PROFILE_KEY0;
                    ack.read_miss = handcode_error_MAP_PROFILE_KEY0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h38,4'b100?,4'h?,1'b?},
           {44'h38A?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PROFILE_KEY_INVERT0;
                    ack.read_miss = handcode_error_MAP_PROFILE_KEY_INVERT0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h38,4'b110?,4'h?,1'b?},
           {44'h38E?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PROFILE_KEY1;
                    ack.read_miss = handcode_error_MAP_PROFILE_KEY1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h39,4'b000?,4'h?,1'b?},
           {44'h392?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PROFILE_KEY_INVERT1;
                    ack.read_miss = handcode_error_MAP_PROFILE_KEY_INVERT1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h39,4'b010?,4'h?,1'b?},
           {44'h396?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_PROFILE_ACTION;
                    ack.read_miss = handcode_error_MAP_PROFILE_ACTION;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h3980,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_DOMAIN_POL_CFG;
                    ack.read_miss = handcode_error_MAP_DOMAIN_POL_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h3A??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MAP_REWRITE;
                    ack.read_miss = handcode_error_MAP_REWRITE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_MAPPER_MAP_MEM) 
           {44'b0???,1'b?},
           {44'h8,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PORT_CFG;
                    ack.write_miss = handcode_error_MAP_PORT_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'b1???0?,1'b?},
           {44'b1???10,1'b?},
           {44'b10???0?,1'b?},
           {44'b10???10,1'b?},
           {40'h6,4'b0?0?,1'b?},
           {40'h6,4'b0?10,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PORT_DEFAULT;
                    ack.write_miss = handcode_error_MAP_PORT_DEFAULT;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h1???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_DOMAIN_TCAM;
                    ack.write_miss = handcode_error_MAP_DOMAIN_TCAM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h2,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_DOMAIN_ACTION0;
                    ack.write_miss = handcode_error_MAP_DOMAIN_ACTION0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h2,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_DOMAIN_ACTION1;
                    ack.write_miss = handcode_error_MAP_DOMAIN_ACTION1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h30,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_DOMAIN_PROFILE;
                    ack.write_miss = handcode_error_MAP_DOMAIN_PROFILE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h310,4'b0???,1'b?},
           {44'h3108,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PORT;
                    ack.write_miss = handcode_error_MAP_PORT;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h31,4'b10??,4'h?,1'b0},
           {36'h31,4'b110?,4'h?,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_MAC;
                    ack.write_miss = handcode_error_MAP_MAC;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h320,4'b1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_IP_LO;
                    ack.write_miss = handcode_error_MAP_IP_LO;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h321,4'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_IP_HI;
                    ack.write_miss = handcode_error_MAP_IP_HI;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h321,4'b1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_IP_CFG;
                    ack.write_miss = handcode_error_MAP_IP_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h322,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PROT;
                    ack.write_miss = handcode_error_MAP_PROT;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h32,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_L4_SRC;
                    ack.write_miss = handcode_error_MAP_L4_SRC;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h32,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_L4_DST;
                    ack.write_miss = handcode_error_MAP_L4_DST;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h328?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_EXP_TC;
                    ack.write_miss = handcode_error_MAP_EXP_TC;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h3,4'b01??,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_DSCP_TC;
                    ack.write_miss = handcode_error_MAP_DSCP_TC;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h380?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_VPRI_TC;
                    ack.write_miss = handcode_error_MAP_VPRI_TC;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h381?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_VPRI;
                    ack.write_miss = handcode_error_MAP_VPRI;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h38,4'b010?,4'h?,1'b?},
           {44'h386?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PROFILE_KEY0;
                    ack.write_miss = handcode_error_MAP_PROFILE_KEY0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h38,4'b100?,4'h?,1'b?},
           {44'h38A?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PROFILE_KEY_INVERT0;
                    ack.write_miss = handcode_error_MAP_PROFILE_KEY_INVERT0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h38,4'b110?,4'h?,1'b?},
           {44'h38E?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PROFILE_KEY1;
                    ack.write_miss = handcode_error_MAP_PROFILE_KEY1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h39,4'b000?,4'h?,1'b?},
           {44'h392?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PROFILE_KEY_INVERT1;
                    ack.write_miss = handcode_error_MAP_PROFILE_KEY_INVERT1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h39,4'b010?,4'h?,1'b?},
           {44'h396?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_PROFILE_ACTION;
                    ack.write_miss = handcode_error_MAP_PROFILE_ACTION;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h3980,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_DOMAIN_POL_CFG;
                    ack.write_miss = handcode_error_MAP_DOMAIN_POL_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h3A??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MAP_REWRITE;
                    ack.write_miss = handcode_error_MAP_REWRITE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_MAPPER_MAP_MEM) 
           {44'b0???,1'b?},
           {44'h8,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PORT_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'b1???0?,1'b?},
           {44'b1???10,1'b?},
           {44'b10???0?,1'b?},
           {44'b10???10,1'b?},
           {40'h6,4'b0?0?,1'b?},
           {40'h6,4'b0?10,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PORT_DEFAULT;
                 default: read_data = '0;
              endcase
           end
           {44'h1???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_DOMAIN_TCAM;
                 default: read_data = '0;
              endcase
           end
           {32'h2,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_DOMAIN_ACTION0;
                 default: read_data = '0;
              endcase
           end
           {32'h2,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_DOMAIN_ACTION1;
                 default: read_data = '0;
              endcase
           end
           {36'h30,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_DOMAIN_PROFILE;
                 default: read_data = '0;
              endcase
           end
           {40'h310,4'b0???,1'b?},
           {44'h3108,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PORT;
                 default: read_data = '0;
              endcase
           end
           {36'h31,4'b10??,4'h?,1'b0},
           {36'h31,4'b110?,4'h?,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_MAC;
                 default: read_data = '0;
              endcase
           end
           {40'h320,4'b1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_IP_LO;
                 default: read_data = '0;
              endcase
           end
           {40'h321,4'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_IP_HI;
                 default: read_data = '0;
              endcase
           end
           {40'h321,4'b1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_IP_CFG;
                 default: read_data = '0;
              endcase
           end
           {40'h322,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PROT;
                 default: read_data = '0;
              endcase
           end
           {36'h32,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_L4_SRC;
                 default: read_data = '0;
              endcase
           end
           {36'h32,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_L4_DST;
                 default: read_data = '0;
              endcase
           end
           {44'h328?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_EXP_TC;
                 default: read_data = '0;
              endcase
           end
           {32'h3,4'b01??,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_DSCP_TC;
                 default: read_data = '0;
              endcase
           end
           {44'h380?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_VPRI_TC;
                 default: read_data = '0;
              endcase
           end
           {44'h381?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_VPRI;
                 default: read_data = '0;
              endcase
           end
           {36'h38,4'b010?,4'h?,1'b?},
           {44'h386?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PROFILE_KEY0;
                 default: read_data = '0;
              endcase
           end
           {36'h38,4'b100?,4'h?,1'b?},
           {44'h38A?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PROFILE_KEY_INVERT0;
                 default: read_data = '0;
              endcase
           end
           {36'h38,4'b110?,4'h?,1'b?},
           {44'h38E?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PROFILE_KEY1;
                 default: read_data = '0;
              endcase
           end
           {36'h39,4'b000?,4'h?,1'b?},
           {44'h392?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PROFILE_KEY_INVERT1;
                 default: read_data = '0;
              endcase
           end
           {36'h39,4'b010?,4'h?,1'b?},
           {44'h396?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_PROFILE_ACTION;
                 default: read_data = '0;
              endcase
           end
           {44'h3980,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_DOMAIN_POL_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'h3A??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MAPPER_SB_FID,MAPPER_SB_BAR}: read_data = handcode_reg_rdata_MAP_REWRITE;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {


// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
