// -----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Raghu P Gudla
// Created On   :  09/22/2018
// Description  :  Full-Chip Config stub
// -----------------------------------------------------------------------------

//`include "fc_liblist.svh"
`ifdef AXI_ENV_ENABLE
`include "axi_svt_dut.sv"
`endif
`ifdef APB_ENV_ENABLE
`include "apb_svt_dut.sv"
`endif
`ifdef CHI_ENV_ENABLE
`include "chi_svt_dut.sv"
`endif

//config `HDL_TOP_CFG;
config fc_hdl_top_cfg;

    design `HDL_TOP_LIB.`HDL_TOP;

    `ifdef FC_MODEL
        `include "fc_config_include.svh";
    `endif

    `ifdef MPP_8
        instance `soc.mby_mpp_1 liblist fc_top_lib;
        instance `soc.mby_mpp_2 liblist fc_top_lib;
        instance `soc.mby_mpp_3 liblist fc_top_lib;
        instance `soc.mby_mpp_4 liblist fc_top_lib;
        instance `soc.mby_mpp_5 liblist fc_top_lib;
        instance `soc.mby_mpp_6 liblist fc_top_lib;
        instance `soc.mby_mpp_7 liblist fc_top_lib;
        instance `soc.mby_mpp_8 liblist fc_top_lib;
    `elsif MPP_2
        instance `soc.mby_mpp_1 liblist fc_top_lib;
        instance `soc.mby_mpp_2 liblist fc_top_lib;
        instance `soc.mby_mpp_3 liblist soc_ip_stub_lib;
        instance `soc.mby_mpp_4 liblist soc_ip_stub_lib;
        instance `soc.mby_mpp_5 liblist soc_ip_stub_lib;
        instance `soc.mby_mpp_6 liblist soc_ip_stub_lib; 
        instance `soc.mby_mpp_7 liblist soc_ip_stub_lib;
        instance `soc.mby_mpp_8 liblist soc_ip_stub_lib;
    `endif

    `ifdef EPC_8
        instance `soc.mby_ec_top_1 liblist fc_top_lib;
        instance `soc.mby_ec_top_2 liblist fc_top_lib;
        instance `soc.mby_ec_top_3 liblist fc_top_lib;
        instance `soc.mby_ec_top_4 liblist fc_top_lib;
        instance `soc.mby_ec_top_5 liblist fc_top_lib;
        instance `soc.mby_ec_top_6 liblist fc_top_lib;
        instance `soc.mby_ec_top_7 liblist fc_top_lib;
        instance `soc.mby_ec_top_8 liblist fc_top_lib;
    `elsif EPC_2
        instance `soc.mby_ec_top_1 liblist fc_top_lib;
        instance `soc.mby_ec_top_2 liblist fc_top_lib;
        instance `soc.mby_ec_top_3 liblist soc_ip_stub_lib;
        instance `soc.mby_ec_top_4 liblist soc_ip_stub_lib;
        instance `soc.mby_ec_top_5 liblist soc_ip_stub_lib;
        instance `soc.mby_ec_top_6 liblist soc_ip_stub_lib; 
        instance `soc.mby_ec_top_7 liblist soc_ip_stub_lib;
        instance `soc.mby_ec_top_8 liblist soc_ip_stub_lib;

    `endif

    `ifdef MPP_WITH_SERDES
    `endif

    `ifdef EPC_WITH_SERDES
    `endif

endconfig


