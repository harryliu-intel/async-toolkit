// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

module mby_checker(

                   );

`include "mby_sva_include.sv"

endmodule 
