///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cgrp_a_nested_map.sv                               
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_cgrp_a_nested_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_RSTD


module rtlgen_mby_ppe_cgrp_a_nested_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_cgrp_a_nested_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_PH2_FF
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CGRP_A_NESTED_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_cgrp_a_nested_map ( //lintra s-2096
    // Clocks


    // Resets



    // Register Inputs
    handcode_reg_rdata_EM_HASH_LOOKUP,
    handcode_reg_rdata_LPM_KEY_MASK,
    handcode_reg_rdata_LPM_KEY_SEL0,
    handcode_reg_rdata_LPM_KEY_SEL1,
    handcode_reg_rdata_LPM_KEY_SEL2,
    handcode_reg_rdata_LPM_KEY_SEL3,
    handcode_reg_rdata_LPM_MATCH_ACTION,
    handcode_reg_rdata_LPM_MATCH_TCAM,
    handcode_reg_rdata_LPM_SUBTRIE_APTR,
    handcode_reg_rdata_LPM_SUBTRIE_BITMAPS,
    handcode_reg_rdata_LPM_SUBTRIE_CPTR,

    handcode_rvalid_EM_HASH_LOOKUP,
    handcode_rvalid_LPM_KEY_MASK,
    handcode_rvalid_LPM_KEY_SEL0,
    handcode_rvalid_LPM_KEY_SEL1,
    handcode_rvalid_LPM_KEY_SEL2,
    handcode_rvalid_LPM_KEY_SEL3,
    handcode_rvalid_LPM_MATCH_ACTION,
    handcode_rvalid_LPM_MATCH_TCAM,
    handcode_rvalid_LPM_SUBTRIE_APTR,
    handcode_rvalid_LPM_SUBTRIE_BITMAPS,
    handcode_rvalid_LPM_SUBTRIE_CPTR,

    handcode_wvalid_EM_HASH_LOOKUP,
    handcode_wvalid_LPM_KEY_MASK,
    handcode_wvalid_LPM_KEY_SEL0,
    handcode_wvalid_LPM_KEY_SEL1,
    handcode_wvalid_LPM_KEY_SEL2,
    handcode_wvalid_LPM_KEY_SEL3,
    handcode_wvalid_LPM_MATCH_ACTION,
    handcode_wvalid_LPM_MATCH_TCAM,
    handcode_wvalid_LPM_SUBTRIE_APTR,
    handcode_wvalid_LPM_SUBTRIE_BITMAPS,
    handcode_wvalid_LPM_SUBTRIE_CPTR,

    handcode_error_EM_HASH_LOOKUP,
    handcode_error_LPM_KEY_MASK,
    handcode_error_LPM_KEY_SEL0,
    handcode_error_LPM_KEY_SEL1,
    handcode_error_LPM_KEY_SEL2,
    handcode_error_LPM_KEY_SEL3,
    handcode_error_LPM_MATCH_ACTION,
    handcode_error_LPM_MATCH_TCAM,
    handcode_error_LPM_SUBTRIE_APTR,
    handcode_error_LPM_SUBTRIE_BITMAPS,
    handcode_error_LPM_SUBTRIE_CPTR,


    // Register Outputs

    // Register signals for HandCoded registers
    handcode_reg_wdata_EM_HASH_LOOKUP,
    handcode_reg_wdata_LPM_KEY_MASK,
    handcode_reg_wdata_LPM_KEY_SEL0,
    handcode_reg_wdata_LPM_KEY_SEL1,
    handcode_reg_wdata_LPM_KEY_SEL2,
    handcode_reg_wdata_LPM_KEY_SEL3,
    handcode_reg_wdata_LPM_MATCH_ACTION,
    handcode_reg_wdata_LPM_MATCH_TCAM,
    handcode_reg_wdata_LPM_SUBTRIE_APTR,
    handcode_reg_wdata_LPM_SUBTRIE_BITMAPS,
    handcode_reg_wdata_LPM_SUBTRIE_CPTR,

    we_EM_HASH_LOOKUP,
    we_LPM_KEY_MASK,
    we_LPM_KEY_SEL0,
    we_LPM_KEY_SEL1,
    we_LPM_KEY_SEL2,
    we_LPM_KEY_SEL3,
    we_LPM_MATCH_ACTION,
    we_LPM_MATCH_TCAM,
    we_LPM_SUBTRIE_APTR,
    we_LPM_SUBTRIE_BITMAPS,
    we_LPM_SUBTRIE_CPTR,

    re_EM_HASH_LOOKUP,
    re_LPM_KEY_MASK,
    re_LPM_KEY_SEL0,
    re_LPM_KEY_SEL1,
    re_LPM_KEY_SEL2,
    re_LPM_KEY_SEL3,
    re_LPM_MATCH_ACTION,
    re_LPM_MATCH_TCAM,
    re_LPM_SUBTRIE_APTR,
    re_LPM_SUBTRIE_BITMAPS,
    re_LPM_SUBTRIE_CPTR,




    // Config Access
    req,
    ack
    

);

import mby_ppe_cgrp_a_nested_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:0] MBY_PPE_CGRP_A_NESTED_MAP_OFFSET = {MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] A_SB_BAR = 3'b0;
parameter [7:0] A_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;

    // Clocks


    // Resets



    // Register Inputs
input EM_HASH_LOOKUP_t  handcode_reg_rdata_EM_HASH_LOOKUP;
input LPM_KEY_MASK_t  handcode_reg_rdata_LPM_KEY_MASK;
input LPM_KEY_SEL0_t  handcode_reg_rdata_LPM_KEY_SEL0;
input LPM_KEY_SEL1_t  handcode_reg_rdata_LPM_KEY_SEL1;
input LPM_KEY_SEL2_t  handcode_reg_rdata_LPM_KEY_SEL2;
input LPM_KEY_SEL3_t  handcode_reg_rdata_LPM_KEY_SEL3;
input LPM_MATCH_ACTION_t  handcode_reg_rdata_LPM_MATCH_ACTION;
input LPM_MATCH_TCAM_t  handcode_reg_rdata_LPM_MATCH_TCAM;
input LPM_SUBTRIE_APTR_t  handcode_reg_rdata_LPM_SUBTRIE_APTR;
input LPM_SUBTRIE_BITMAPS_t  handcode_reg_rdata_LPM_SUBTRIE_BITMAPS;
input LPM_SUBTRIE_CPTR_t  handcode_reg_rdata_LPM_SUBTRIE_CPTR;

input handcode_rvalid_EM_HASH_LOOKUP_t  handcode_rvalid_EM_HASH_LOOKUP;
input handcode_rvalid_LPM_KEY_MASK_t  handcode_rvalid_LPM_KEY_MASK;
input handcode_rvalid_LPM_KEY_SEL0_t  handcode_rvalid_LPM_KEY_SEL0;
input handcode_rvalid_LPM_KEY_SEL1_t  handcode_rvalid_LPM_KEY_SEL1;
input handcode_rvalid_LPM_KEY_SEL2_t  handcode_rvalid_LPM_KEY_SEL2;
input handcode_rvalid_LPM_KEY_SEL3_t  handcode_rvalid_LPM_KEY_SEL3;
input handcode_rvalid_LPM_MATCH_ACTION_t  handcode_rvalid_LPM_MATCH_ACTION;
input handcode_rvalid_LPM_MATCH_TCAM_t  handcode_rvalid_LPM_MATCH_TCAM;
input handcode_rvalid_LPM_SUBTRIE_APTR_t  handcode_rvalid_LPM_SUBTRIE_APTR;
input handcode_rvalid_LPM_SUBTRIE_BITMAPS_t  handcode_rvalid_LPM_SUBTRIE_BITMAPS;
input handcode_rvalid_LPM_SUBTRIE_CPTR_t  handcode_rvalid_LPM_SUBTRIE_CPTR;

input handcode_wvalid_EM_HASH_LOOKUP_t  handcode_wvalid_EM_HASH_LOOKUP;
input handcode_wvalid_LPM_KEY_MASK_t  handcode_wvalid_LPM_KEY_MASK;
input handcode_wvalid_LPM_KEY_SEL0_t  handcode_wvalid_LPM_KEY_SEL0;
input handcode_wvalid_LPM_KEY_SEL1_t  handcode_wvalid_LPM_KEY_SEL1;
input handcode_wvalid_LPM_KEY_SEL2_t  handcode_wvalid_LPM_KEY_SEL2;
input handcode_wvalid_LPM_KEY_SEL3_t  handcode_wvalid_LPM_KEY_SEL3;
input handcode_wvalid_LPM_MATCH_ACTION_t  handcode_wvalid_LPM_MATCH_ACTION;
input handcode_wvalid_LPM_MATCH_TCAM_t  handcode_wvalid_LPM_MATCH_TCAM;
input handcode_wvalid_LPM_SUBTRIE_APTR_t  handcode_wvalid_LPM_SUBTRIE_APTR;
input handcode_wvalid_LPM_SUBTRIE_BITMAPS_t  handcode_wvalid_LPM_SUBTRIE_BITMAPS;
input handcode_wvalid_LPM_SUBTRIE_CPTR_t  handcode_wvalid_LPM_SUBTRIE_CPTR;

input handcode_error_EM_HASH_LOOKUP_t  handcode_error_EM_HASH_LOOKUP;
input handcode_error_LPM_KEY_MASK_t  handcode_error_LPM_KEY_MASK;
input handcode_error_LPM_KEY_SEL0_t  handcode_error_LPM_KEY_SEL0;
input handcode_error_LPM_KEY_SEL1_t  handcode_error_LPM_KEY_SEL1;
input handcode_error_LPM_KEY_SEL2_t  handcode_error_LPM_KEY_SEL2;
input handcode_error_LPM_KEY_SEL3_t  handcode_error_LPM_KEY_SEL3;
input handcode_error_LPM_MATCH_ACTION_t  handcode_error_LPM_MATCH_ACTION;
input handcode_error_LPM_MATCH_TCAM_t  handcode_error_LPM_MATCH_TCAM;
input handcode_error_LPM_SUBTRIE_APTR_t  handcode_error_LPM_SUBTRIE_APTR;
input handcode_error_LPM_SUBTRIE_BITMAPS_t  handcode_error_LPM_SUBTRIE_BITMAPS;
input handcode_error_LPM_SUBTRIE_CPTR_t  handcode_error_LPM_SUBTRIE_CPTR;


    // Register Outputs

    // Register signals for HandCoded registers
output EM_HASH_LOOKUP_t  handcode_reg_wdata_EM_HASH_LOOKUP;
output LPM_KEY_MASK_t  handcode_reg_wdata_LPM_KEY_MASK;
output LPM_KEY_SEL0_t  handcode_reg_wdata_LPM_KEY_SEL0;
output LPM_KEY_SEL1_t  handcode_reg_wdata_LPM_KEY_SEL1;
output LPM_KEY_SEL2_t  handcode_reg_wdata_LPM_KEY_SEL2;
output LPM_KEY_SEL3_t  handcode_reg_wdata_LPM_KEY_SEL3;
output LPM_MATCH_ACTION_t  handcode_reg_wdata_LPM_MATCH_ACTION;
output LPM_MATCH_TCAM_t  handcode_reg_wdata_LPM_MATCH_TCAM;
output LPM_SUBTRIE_APTR_t  handcode_reg_wdata_LPM_SUBTRIE_APTR;
output LPM_SUBTRIE_BITMAPS_t  handcode_reg_wdata_LPM_SUBTRIE_BITMAPS;
output LPM_SUBTRIE_CPTR_t  handcode_reg_wdata_LPM_SUBTRIE_CPTR;

output we_EM_HASH_LOOKUP_t  we_EM_HASH_LOOKUP;
output we_LPM_KEY_MASK_t  we_LPM_KEY_MASK;
output we_LPM_KEY_SEL0_t  we_LPM_KEY_SEL0;
output we_LPM_KEY_SEL1_t  we_LPM_KEY_SEL1;
output we_LPM_KEY_SEL2_t  we_LPM_KEY_SEL2;
output we_LPM_KEY_SEL3_t  we_LPM_KEY_SEL3;
output we_LPM_MATCH_ACTION_t  we_LPM_MATCH_ACTION;
output we_LPM_MATCH_TCAM_t  we_LPM_MATCH_TCAM;
output we_LPM_SUBTRIE_APTR_t  we_LPM_SUBTRIE_APTR;
output we_LPM_SUBTRIE_BITMAPS_t  we_LPM_SUBTRIE_BITMAPS;
output we_LPM_SUBTRIE_CPTR_t  we_LPM_SUBTRIE_CPTR;

output re_EM_HASH_LOOKUP_t  re_EM_HASH_LOOKUP;
output re_LPM_KEY_MASK_t  re_LPM_KEY_MASK;
output re_LPM_KEY_SEL0_t  re_LPM_KEY_SEL0;
output re_LPM_KEY_SEL1_t  re_LPM_KEY_SEL1;
output re_LPM_KEY_SEL2_t  re_LPM_KEY_SEL2;
output re_LPM_KEY_SEL3_t  re_LPM_KEY_SEL3;
output re_LPM_MATCH_ACTION_t  re_LPM_MATCH_ACTION;
output re_LPM_MATCH_TCAM_t  re_LPM_MATCH_TCAM;
output re_LPM_SUBTRIE_APTR_t  re_LPM_SUBTRIE_APTR;
output re_LPM_SUBTRIE_BITMAPS_t  re_LPM_SUBTRIE_BITMAPS;
output re_LPM_SUBTRIE_CPTR_t  re_LPM_SUBTRIE_CPTR;




    // Config Access
input mby_ppe_cgrp_a_nested_map_cr_req_t  req;
output mby_ppe_cgrp_a_nested_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_cgrp_a_nested_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_CGRP_A_NESTED_MAP_MEM;
assign case_req_addr_MBY_PPE_CGRP_A_NESTED_MAP_MEM = req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_a;
always_comb begin : sb_fid_cond_a_BLOCK
    unique casez (req_fid) 
		A_SB_FID: sb_fid_cond_a = 1;
		default: sb_fid_cond_a = 0;
    endcase 
end


logic sb_bar_cond_a;
always_comb begin : sb_bar_cond_a_BLOCK
    unique casez (req_bar) 
		A_SB_BAR: sb_bar_cond_a = 1;
		default: sb_bar_cond_a = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// EM_HASH_LOOKUP using HANDCODED_REG template.
logic addr_decode_EM_HASH_LOOKUP;
logic write_req_EM_HASH_LOOKUP;
logic read_req_EM_HASH_LOOKUP;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b0???,12'h???,1'b0}: 
         addr_decode_EM_HASH_LOOKUP = req.valid;
      default: 
         addr_decode_EM_HASH_LOOKUP = 1'b0; 
   endcase
end

always_comb write_req_EM_HASH_LOOKUP = f_IsMEMWr(req_opcode) && addr_decode_EM_HASH_LOOKUP ;
always_comb read_req_EM_HASH_LOOKUP  = f_IsMEMRd(req_opcode) && addr_decode_EM_HASH_LOOKUP ;

always_comb we_EM_HASH_LOOKUP = {16{write_req_EM_HASH_LOOKUP}} & req.be[15:0];
always_comb re_EM_HASH_LOOKUP = {16{read_req_EM_HASH_LOOKUP}} & req.be[15:0];
always_comb handcode_reg_wdata_EM_HASH_LOOKUP = req.data[127:0];


// ----------------------------------------------------------------------
// LPM_SUBTRIE_APTR using HANDCODED_REG template.
logic addr_decode_LPM_SUBTRIE_APTR;
logic write_req_LPM_SUBTRIE_APTR;
logic read_req_LPM_SUBTRIE_APTR;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b100?,12'h???,1'b?},
      {44'hA???,1'b?}:
          addr_decode_LPM_SUBTRIE_APTR = req.valid;
      default: 
         addr_decode_LPM_SUBTRIE_APTR = 1'b0; 
   endcase
end

always_comb write_req_LPM_SUBTRIE_APTR = f_IsMEMWr(req_opcode) && addr_decode_LPM_SUBTRIE_APTR ;
always_comb read_req_LPM_SUBTRIE_APTR  = f_IsMEMRd(req_opcode) && addr_decode_LPM_SUBTRIE_APTR ;

always_comb we_LPM_SUBTRIE_APTR = {8{write_req_LPM_SUBTRIE_APTR}} & be;
always_comb re_LPM_SUBTRIE_APTR = {8{read_req_LPM_SUBTRIE_APTR}} & be;
always_comb handcode_reg_wdata_LPM_SUBTRIE_APTR = write_data;


// ----------------------------------------------------------------------
// LPM_SUBTRIE_CPTR using HANDCODED_REG template.
logic addr_decode_LPM_SUBTRIE_CPTR;
logic write_req_LPM_SUBTRIE_CPTR;
logic read_req_LPM_SUBTRIE_CPTR;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b110?,12'h???,1'b?},
      {44'hE???,1'b?}:
          addr_decode_LPM_SUBTRIE_CPTR = req.valid;
      default: 
         addr_decode_LPM_SUBTRIE_CPTR = 1'b0; 
   endcase
end

always_comb write_req_LPM_SUBTRIE_CPTR = f_IsMEMWr(req_opcode) && addr_decode_LPM_SUBTRIE_CPTR ;
always_comb read_req_LPM_SUBTRIE_CPTR  = f_IsMEMRd(req_opcode) && addr_decode_LPM_SUBTRIE_CPTR ;

always_comb we_LPM_SUBTRIE_CPTR = {8{write_req_LPM_SUBTRIE_CPTR}} & be;
always_comb re_LPM_SUBTRIE_CPTR = {8{read_req_LPM_SUBTRIE_CPTR}} & be;
always_comb handcode_reg_wdata_LPM_SUBTRIE_CPTR = write_data;


// ----------------------------------------------------------------------
// LPM_SUBTRIE_BITMAPS using HANDCODED_REG template.
logic addr_decode_LPM_SUBTRIE_BITMAPS;
logic write_req_LPM_SUBTRIE_BITMAPS;
logic read_req_LPM_SUBTRIE_BITMAPS;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h2????,1'b?},
      {28'h3,4'b0???,12'h???,1'b?}:
          addr_decode_LPM_SUBTRIE_BITMAPS = req.valid;
      default: 
         addr_decode_LPM_SUBTRIE_BITMAPS = 1'b0; 
   endcase
end

always_comb write_req_LPM_SUBTRIE_BITMAPS = f_IsMEMWr(req_opcode) && addr_decode_LPM_SUBTRIE_BITMAPS ;
always_comb read_req_LPM_SUBTRIE_BITMAPS  = f_IsMEMRd(req_opcode) && addr_decode_LPM_SUBTRIE_BITMAPS ;

always_comb we_LPM_SUBTRIE_BITMAPS = {8{write_req_LPM_SUBTRIE_BITMAPS}} & be;
always_comb re_LPM_SUBTRIE_BITMAPS = {8{read_req_LPM_SUBTRIE_BITMAPS}} & be;
always_comb handcode_reg_wdata_LPM_SUBTRIE_BITMAPS = write_data;


// ----------------------------------------------------------------------
// LPM_MATCH_TCAM using HANDCODED_REG template.
logic addr_decode_LPM_MATCH_TCAM;
logic write_req_LPM_MATCH_TCAM;
logic read_req_LPM_MATCH_TCAM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h380??,1'b?}: 
         addr_decode_LPM_MATCH_TCAM = req.valid;
      default: 
         addr_decode_LPM_MATCH_TCAM = 1'b0; 
   endcase
end

always_comb write_req_LPM_MATCH_TCAM = f_IsMEMWr(req_opcode) && addr_decode_LPM_MATCH_TCAM ;
always_comb read_req_LPM_MATCH_TCAM  = f_IsMEMRd(req_opcode) && addr_decode_LPM_MATCH_TCAM ;

always_comb we_LPM_MATCH_TCAM = {8{write_req_LPM_MATCH_TCAM}} & be;
always_comb re_LPM_MATCH_TCAM = {8{read_req_LPM_MATCH_TCAM}} & be;
always_comb handcode_reg_wdata_LPM_MATCH_TCAM = write_data;


// ----------------------------------------------------------------------
// LPM_MATCH_ACTION using HANDCODED_REG template.
logic addr_decode_LPM_MATCH_ACTION;
logic write_req_LPM_MATCH_ACTION;
logic read_req_LPM_MATCH_ACTION;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h381??,1'b?}: 
         addr_decode_LPM_MATCH_ACTION = req.valid;
      default: 
         addr_decode_LPM_MATCH_ACTION = 1'b0; 
   endcase
end

always_comb write_req_LPM_MATCH_ACTION = f_IsMEMWr(req_opcode) && addr_decode_LPM_MATCH_ACTION ;
always_comb read_req_LPM_MATCH_ACTION  = f_IsMEMRd(req_opcode) && addr_decode_LPM_MATCH_ACTION ;

always_comb we_LPM_MATCH_ACTION = {8{write_req_LPM_MATCH_ACTION}} & be;
always_comb re_LPM_MATCH_ACTION = {8{read_req_LPM_MATCH_ACTION}} & be;
always_comb handcode_reg_wdata_LPM_MATCH_ACTION = write_data;


// ----------------------------------------------------------------------
// LPM_KEY_MASK using HANDCODED_REG template.
logic addr_decode_LPM_KEY_MASK;
logic write_req_LPM_KEY_MASK;
logic read_req_LPM_KEY_MASK;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h38,4'b01??,4'h?,4'b0???,1'b?},
      {32'h38,4'b01??,4'h?,4'b100?,1'b?}:
          addr_decode_LPM_KEY_MASK = req.valid;
      default: 
         addr_decode_LPM_KEY_MASK = 1'b0; 
   endcase
end

always_comb write_req_LPM_KEY_MASK = f_IsMEMWr(req_opcode) && addr_decode_LPM_KEY_MASK ;
always_comb read_req_LPM_KEY_MASK  = f_IsMEMRd(req_opcode) && addr_decode_LPM_KEY_MASK ;

always_comb we_LPM_KEY_MASK = {8{write_req_LPM_KEY_MASK}} & be;
always_comb re_LPM_KEY_MASK = {8{read_req_LPM_KEY_MASK}} & be;
always_comb handcode_reg_wdata_LPM_KEY_MASK = write_data;


// ----------------------------------------------------------------------
// LPM_KEY_SEL0 using HANDCODED_REG template.
logic addr_decode_LPM_KEY_SEL0;
logic write_req_LPM_KEY_SEL0;
logic read_req_LPM_KEY_SEL0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h388,4'b000?,4'h?,1'b?}: 
         addr_decode_LPM_KEY_SEL0 = req.valid;
      default: 
         addr_decode_LPM_KEY_SEL0 = 1'b0; 
   endcase
end

always_comb write_req_LPM_KEY_SEL0 = f_IsMEMWr(req_opcode) && addr_decode_LPM_KEY_SEL0 ;
always_comb read_req_LPM_KEY_SEL0  = f_IsMEMRd(req_opcode) && addr_decode_LPM_KEY_SEL0 ;

always_comb we_LPM_KEY_SEL0 = {8{write_req_LPM_KEY_SEL0}} & be;
always_comb re_LPM_KEY_SEL0 = {8{read_req_LPM_KEY_SEL0}} & be;
always_comb handcode_reg_wdata_LPM_KEY_SEL0 = write_data;


// ----------------------------------------------------------------------
// LPM_KEY_SEL1 using HANDCODED_REG template.
logic addr_decode_LPM_KEY_SEL1;
logic write_req_LPM_KEY_SEL1;
logic read_req_LPM_KEY_SEL1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h388,4'b001?,4'h?,1'b?}: 
         addr_decode_LPM_KEY_SEL1 = req.valid;
      default: 
         addr_decode_LPM_KEY_SEL1 = 1'b0; 
   endcase
end

always_comb write_req_LPM_KEY_SEL1 = f_IsMEMWr(req_opcode) && addr_decode_LPM_KEY_SEL1 ;
always_comb read_req_LPM_KEY_SEL1  = f_IsMEMRd(req_opcode) && addr_decode_LPM_KEY_SEL1 ;

always_comb we_LPM_KEY_SEL1 = {8{write_req_LPM_KEY_SEL1}} & be;
always_comb re_LPM_KEY_SEL1 = {8{read_req_LPM_KEY_SEL1}} & be;
always_comb handcode_reg_wdata_LPM_KEY_SEL1 = write_data;


// ----------------------------------------------------------------------
// LPM_KEY_SEL2 using HANDCODED_REG template.
logic addr_decode_LPM_KEY_SEL2;
logic write_req_LPM_KEY_SEL2;
logic read_req_LPM_KEY_SEL2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h388,4'b010?,4'h?,1'b?}: 
         addr_decode_LPM_KEY_SEL2 = req.valid;
      default: 
         addr_decode_LPM_KEY_SEL2 = 1'b0; 
   endcase
end

always_comb write_req_LPM_KEY_SEL2 = f_IsMEMWr(req_opcode) && addr_decode_LPM_KEY_SEL2 ;
always_comb read_req_LPM_KEY_SEL2  = f_IsMEMRd(req_opcode) && addr_decode_LPM_KEY_SEL2 ;

always_comb we_LPM_KEY_SEL2 = {8{write_req_LPM_KEY_SEL2}} & be;
always_comb re_LPM_KEY_SEL2 = {8{read_req_LPM_KEY_SEL2}} & be;
always_comb handcode_reg_wdata_LPM_KEY_SEL2 = write_data;


// ----------------------------------------------------------------------
// LPM_KEY_SEL3 using HANDCODED_REG template.
logic addr_decode_LPM_KEY_SEL3;
logic write_req_LPM_KEY_SEL3;
logic read_req_LPM_KEY_SEL3;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_A_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h388,4'b011?,4'h?,1'b?}: 
         addr_decode_LPM_KEY_SEL3 = req.valid;
      default: 
         addr_decode_LPM_KEY_SEL3 = 1'b0; 
   endcase
end

always_comb write_req_LPM_KEY_SEL3 = f_IsMEMWr(req_opcode) && addr_decode_LPM_KEY_SEL3 ;
always_comb read_req_LPM_KEY_SEL3  = f_IsMEMRd(req_opcode) && addr_decode_LPM_KEY_SEL3 ;

always_comb we_LPM_KEY_SEL3 = {8{write_req_LPM_KEY_SEL3}} & be;
always_comb re_LPM_KEY_SEL3 = {8{read_req_LPM_KEY_SEL3}} & be;
always_comb handcode_reg_wdata_LPM_KEY_SEL3 = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_CGRP_A_NESTED_MAP_MEM) 
           {32'b0???,12'h???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_EM_HASH_LOOKUP;
                    ack.read_miss = handcode_error_EM_HASH_LOOKUP;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b100?,12'h???,1'b?},
           {44'hA???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_SUBTRIE_APTR;
                    ack.read_miss = handcode_error_LPM_SUBTRIE_APTR;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b110?,12'h???,1'b?},
           {44'hE???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_SUBTRIE_CPTR;
                    ack.read_miss = handcode_error_LPM_SUBTRIE_CPTR;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h2????,1'b?},
           {28'h3,4'b0???,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_SUBTRIE_BITMAPS;
                    ack.read_miss = handcode_error_LPM_SUBTRIE_BITMAPS;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h380??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_MATCH_TCAM;
                    ack.read_miss = handcode_error_LPM_MATCH_TCAM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h381??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_MATCH_ACTION;
                    ack.read_miss = handcode_error_LPM_MATCH_ACTION;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h38,4'b01??,4'h?,4'b0???,1'b?},
           {32'h38,4'b01??,4'h?,4'b100?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_KEY_MASK;
                    ack.read_miss = handcode_error_LPM_KEY_MASK;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h388,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_KEY_SEL0;
                    ack.read_miss = handcode_error_LPM_KEY_SEL0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h388,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_KEY_SEL1;
                    ack.read_miss = handcode_error_LPM_KEY_SEL1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h388,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_KEY_SEL2;
                    ack.read_miss = handcode_error_LPM_KEY_SEL2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h388,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_LPM_KEY_SEL3;
                    ack.read_miss = handcode_error_LPM_KEY_SEL3;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_CGRP_A_NESTED_MAP_MEM) 
           {32'b0???,12'h???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_EM_HASH_LOOKUP;
                    ack.write_miss = handcode_error_EM_HASH_LOOKUP;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b100?,12'h???,1'b?},
           {44'hA???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_SUBTRIE_APTR;
                    ack.write_miss = handcode_error_LPM_SUBTRIE_APTR;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b110?,12'h???,1'b?},
           {44'hE???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_SUBTRIE_CPTR;
                    ack.write_miss = handcode_error_LPM_SUBTRIE_CPTR;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h2????,1'b?},
           {28'h3,4'b0???,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_SUBTRIE_BITMAPS;
                    ack.write_miss = handcode_error_LPM_SUBTRIE_BITMAPS;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h380??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_MATCH_TCAM;
                    ack.write_miss = handcode_error_LPM_MATCH_TCAM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h381??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_MATCH_ACTION;
                    ack.write_miss = handcode_error_LPM_MATCH_ACTION;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h38,4'b01??,4'h?,4'b0???,1'b?},
           {32'h38,4'b01??,4'h?,4'b100?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_KEY_MASK;
                    ack.write_miss = handcode_error_LPM_KEY_MASK;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h388,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_KEY_SEL0;
                    ack.write_miss = handcode_error_LPM_KEY_SEL0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h388,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_KEY_SEL1;
                    ack.write_miss = handcode_error_LPM_KEY_SEL1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h388,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_KEY_SEL2;
                    ack.write_miss = handcode_error_LPM_KEY_SEL2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h388,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_LPM_KEY_SEL3;
                    ack.write_miss = handcode_error_LPM_KEY_SEL3;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_CGRP_A_NESTED_MAP_MEM) 
           {32'b0???,12'h???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_EM_HASH_LOOKUP;
                 default: read_data = '0;
              endcase
           end
           {32'b100?,12'h???,1'b?},
           {44'hA???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_SUBTRIE_APTR;
                 default: read_data = '0;
              endcase
           end
           {32'b110?,12'h???,1'b?},
           {44'hE???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_SUBTRIE_CPTR;
                 default: read_data = '0;
              endcase
           end
           {44'h2????,1'b?},
           {28'h3,4'b0???,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_SUBTRIE_BITMAPS;
                 default: read_data = '0;
              endcase
           end
           {44'h380??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_MATCH_TCAM;
                 default: read_data = '0;
              endcase
           end
           {44'h381??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_MATCH_ACTION;
                 default: read_data = '0;
              endcase
           end
           {32'h38,4'b01??,4'h?,4'b0???,1'b?},
           {32'h38,4'b01??,4'h?,4'b100?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_KEY_MASK;
                 default: read_data = '0;
              endcase
           end
           {36'h388,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_KEY_SEL0;
                 default: read_data = '0;
              endcase
           end
           {36'h388,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_KEY_SEL1;
                 default: read_data = '0;
              endcase
           end
           {36'h388,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_KEY_SEL2;
                 default: read_data = '0;
              endcase
           end
           {36'h388,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {A_SB_FID,A_SB_BAR}: read_data = handcode_reg_rdata_LPM_KEY_SEL3;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {


// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
