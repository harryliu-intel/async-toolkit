///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_rx_voq_map.sv                                          
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_rx_voq_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_RX_VOQ_MAP_FF
`define RTLGEN_MBY_RX_VOQ_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_RX_VOQ_MAP_FF

`ifndef RTLGEN_MBY_RX_VOQ_MAP_EN_FF
`define RTLGEN_MBY_RX_VOQ_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_RX_VOQ_MAP_EN_FF

`ifndef RTLGEN_MBY_RX_VOQ_MAP_FF_RSTD
`define RTLGEN_MBY_RX_VOQ_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_RX_VOQ_MAP_FF_RSTD


module rtlgen_mby_rx_voq_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_RX_VOQ_MAP_EN_FF_RSTD
`define RTLGEN_MBY_RX_VOQ_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_rx_voq_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_RX_VOQ_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_RX_VOQ_MAP_FF_SYNCRST
`define RTLGEN_MBY_RX_VOQ_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_RX_VOQ_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_RX_VOQ_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_RX_VOQ_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_RX_VOQ_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_RX_VOQ_MAP_FF_BOTHRST
// `define RTLGEN_MBY_RX_VOQ_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_RX_VOQ_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_RX_VOQ_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_RX_VOQ_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_RX_VOQ_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_RX_VOQ_MAP_LATCH_LOW
`define RTLGEN_MBY_RX_VOQ_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_RX_VOQ_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_RX_VOQ_MAP_PH2_FF
`define RTLGEN_MBY_RX_VOQ_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_RX_VOQ_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_RX_VOQ_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_RX_VOQ_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_RX_VOQ_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_RX_VOQ_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_RX_VOQ_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_RX_VOQ_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_RX_VOQ_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_RX_VOQ_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_RX_VOQ_MAP_LATCH
`define RTLGEN_MBY_RX_VOQ_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_RX_VOQ_MAP_LATCH

`ifndef RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH
`define RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH

`ifndef RTLGEN_MBY_RX_VOQ_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_RX_VOQ_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_RX_VOQ_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_RX_VOQ_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_RX_VOQ_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_RX_VOQ_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_RX_VOQ_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_rx_voq_map ( //lintra s-2096
    // Clocks


    // Resets



    // Register Inputs
    handcode_reg_rdata_RX_VOQ_PORT_CFG,
    handcode_reg_rdata_SAF_EGRESS_SPEED,
    handcode_reg_rdata_SAF_INGRESS_SPEED,
    handcode_reg_rdata_SAF_TC,

    handcode_rvalid_RX_VOQ_PORT_CFG,
    handcode_rvalid_SAF_EGRESS_SPEED,
    handcode_rvalid_SAF_INGRESS_SPEED,
    handcode_rvalid_SAF_TC,

    handcode_wvalid_RX_VOQ_PORT_CFG,
    handcode_wvalid_SAF_EGRESS_SPEED,
    handcode_wvalid_SAF_INGRESS_SPEED,
    handcode_wvalid_SAF_TC,

    handcode_error_RX_VOQ_PORT_CFG,
    handcode_error_SAF_EGRESS_SPEED,
    handcode_error_SAF_INGRESS_SPEED,
    handcode_error_SAF_TC,


    // Register Outputs

    // Register signals for HandCoded registers
    handcode_reg_wdata_RX_VOQ_PORT_CFG,
    handcode_reg_wdata_SAF_EGRESS_SPEED,
    handcode_reg_wdata_SAF_INGRESS_SPEED,
    handcode_reg_wdata_SAF_TC,

    we_RX_VOQ_PORT_CFG,
    we_SAF_EGRESS_SPEED,
    we_SAF_INGRESS_SPEED,
    we_SAF_TC,

    re_RX_VOQ_PORT_CFG,
    re_SAF_EGRESS_SPEED,
    re_SAF_INGRESS_SPEED,
    re_SAF_TC,




    // Config Access
    req,
    ack
    

);

import mby_rx_voq_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_RX_VOQ_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_RX_VOQ_MAP_MEM_ADDR_MSB:0] MBY_RX_VOQ_MAP_OFFSET = {MBY_RX_VOQ_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] RX_VOQ_SB_BAR = 3'b0;
parameter [7:0] RX_VOQ_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;

    // Clocks


    // Resets



    // Register Inputs
input RX_VOQ_PORT_CFG_t  handcode_reg_rdata_RX_VOQ_PORT_CFG;
input SAF_EGRESS_SPEED_t  handcode_reg_rdata_SAF_EGRESS_SPEED;
input SAF_INGRESS_SPEED_t  handcode_reg_rdata_SAF_INGRESS_SPEED;
input SAF_TC_t  handcode_reg_rdata_SAF_TC;

input handcode_rvalid_RX_VOQ_PORT_CFG_t  handcode_rvalid_RX_VOQ_PORT_CFG;
input handcode_rvalid_SAF_EGRESS_SPEED_t  handcode_rvalid_SAF_EGRESS_SPEED;
input handcode_rvalid_SAF_INGRESS_SPEED_t  handcode_rvalid_SAF_INGRESS_SPEED;
input handcode_rvalid_SAF_TC_t  handcode_rvalid_SAF_TC;

input handcode_wvalid_RX_VOQ_PORT_CFG_t  handcode_wvalid_RX_VOQ_PORT_CFG;
input handcode_wvalid_SAF_EGRESS_SPEED_t  handcode_wvalid_SAF_EGRESS_SPEED;
input handcode_wvalid_SAF_INGRESS_SPEED_t  handcode_wvalid_SAF_INGRESS_SPEED;
input handcode_wvalid_SAF_TC_t  handcode_wvalid_SAF_TC;

input handcode_error_RX_VOQ_PORT_CFG_t  handcode_error_RX_VOQ_PORT_CFG;
input handcode_error_SAF_EGRESS_SPEED_t  handcode_error_SAF_EGRESS_SPEED;
input handcode_error_SAF_INGRESS_SPEED_t  handcode_error_SAF_INGRESS_SPEED;
input handcode_error_SAF_TC_t  handcode_error_SAF_TC;


    // Register Outputs

    // Register signals for HandCoded registers
output RX_VOQ_PORT_CFG_t  handcode_reg_wdata_RX_VOQ_PORT_CFG;
output SAF_EGRESS_SPEED_t  handcode_reg_wdata_SAF_EGRESS_SPEED;
output SAF_INGRESS_SPEED_t  handcode_reg_wdata_SAF_INGRESS_SPEED;
output SAF_TC_t  handcode_reg_wdata_SAF_TC;

output we_RX_VOQ_PORT_CFG_t  we_RX_VOQ_PORT_CFG;
output we_SAF_EGRESS_SPEED_t  we_SAF_EGRESS_SPEED;
output we_SAF_INGRESS_SPEED_t  we_SAF_INGRESS_SPEED;
output we_SAF_TC_t  we_SAF_TC;

output re_RX_VOQ_PORT_CFG_t  re_RX_VOQ_PORT_CFG;
output re_SAF_EGRESS_SPEED_t  re_SAF_EGRESS_SPEED;
output re_SAF_INGRESS_SPEED_t  re_SAF_INGRESS_SPEED;
output re_SAF_TC_t  re_SAF_TC;




    // Config Access
input mby_rx_voq_map_cr_req_t  req;
output mby_rx_voq_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_rx_voq_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_RX_VOQ_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_RX_VOQ_MAP_MEM;
assign case_req_addr_MBY_RX_VOQ_MAP_MEM = req_addr[MBY_RX_VOQ_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_rx_voq;
always_comb begin : sb_fid_cond_rx_voq_BLOCK
    unique casez (req_fid) 
		RX_VOQ_SB_FID: sb_fid_cond_rx_voq = 1;
		default: sb_fid_cond_rx_voq = 0;
    endcase 
end


logic sb_bar_cond_rx_voq;
always_comb begin : sb_bar_cond_rx_voq_BLOCK
    unique casez (req_bar) 
		RX_VOQ_SB_BAR: sb_bar_cond_rx_voq = 1;
		default: sb_bar_cond_rx_voq = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// RX_VOQ_PORT_CFG using HANDCODED_REG template.
logic addr_decode_RX_VOQ_PORT_CFG;
logic write_req_RX_VOQ_PORT_CFG;
logic read_req_RX_VOQ_PORT_CFG;

always_comb begin 
   unique casez (req_addr[MBY_RX_VOQ_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h0,1'b0}: 
         addr_decode_RX_VOQ_PORT_CFG = req.valid;
      default: 
         addr_decode_RX_VOQ_PORT_CFG = 1'b0; 
   endcase
end

always_comb write_req_RX_VOQ_PORT_CFG = f_IsMEMWr(req_opcode) && addr_decode_RX_VOQ_PORT_CFG ;
always_comb read_req_RX_VOQ_PORT_CFG  = f_IsMEMRd(req_opcode) && addr_decode_RX_VOQ_PORT_CFG ;

always_comb we_RX_VOQ_PORT_CFG = {8{write_req_RX_VOQ_PORT_CFG}} & be;
always_comb re_RX_VOQ_PORT_CFG = {8{read_req_RX_VOQ_PORT_CFG}} & be;
always_comb handcode_reg_wdata_RX_VOQ_PORT_CFG = write_data;


// ----------------------------------------------------------------------
// SAF_INGRESS_SPEED using HANDCODED_REG template.
logic addr_decode_SAF_INGRESS_SPEED;
logic write_req_SAF_INGRESS_SPEED;
logic read_req_SAF_INGRESS_SPEED;

always_comb begin 
   unique casez (req_addr[MBY_RX_VOQ_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h0,1'b1}: 
         addr_decode_SAF_INGRESS_SPEED = req.valid;
      default: 
         addr_decode_SAF_INGRESS_SPEED = 1'b0; 
   endcase
end

always_comb write_req_SAF_INGRESS_SPEED = f_IsMEMWr(req_opcode) && addr_decode_SAF_INGRESS_SPEED ;
always_comb read_req_SAF_INGRESS_SPEED  = f_IsMEMRd(req_opcode) && addr_decode_SAF_INGRESS_SPEED ;

always_comb we_SAF_INGRESS_SPEED = {8{write_req_SAF_INGRESS_SPEED}} & be;
always_comb re_SAF_INGRESS_SPEED = {8{read_req_SAF_INGRESS_SPEED}} & be;
always_comb handcode_reg_wdata_SAF_INGRESS_SPEED = write_data;


// ----------------------------------------------------------------------
// SAF_EGRESS_SPEED using HANDCODED_REG template.
logic addr_decode_SAF_EGRESS_SPEED;
logic write_req_SAF_EGRESS_SPEED;
logic read_req_SAF_EGRESS_SPEED;

always_comb begin 
   unique casez (req_addr[MBY_RX_VOQ_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b1???,4'h?,1'b?}: 
         addr_decode_SAF_EGRESS_SPEED = req.valid;
      default: 
         addr_decode_SAF_EGRESS_SPEED = 1'b0; 
   endcase
end

always_comb write_req_SAF_EGRESS_SPEED = f_IsMEMWr(req_opcode) && addr_decode_SAF_EGRESS_SPEED ;
always_comb read_req_SAF_EGRESS_SPEED  = f_IsMEMRd(req_opcode) && addr_decode_SAF_EGRESS_SPEED ;

always_comb we_SAF_EGRESS_SPEED = {8{write_req_SAF_EGRESS_SPEED}} & be;
always_comb re_SAF_EGRESS_SPEED = {8{read_req_SAF_EGRESS_SPEED}} & be;
always_comb handcode_reg_wdata_SAF_EGRESS_SPEED = write_data;


// ----------------------------------------------------------------------
// SAF_TC using HANDCODED_REG template.
logic addr_decode_SAF_TC;
logic write_req_SAF_TC;
logic read_req_SAF_TC;

always_comb begin 
   unique casez (req_addr[MBY_RX_VOQ_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h10,4'b0???,1'b?}: 
         addr_decode_SAF_TC = req.valid;
      default: 
         addr_decode_SAF_TC = 1'b0; 
   endcase
end

always_comb write_req_SAF_TC = f_IsMEMWr(req_opcode) && addr_decode_SAF_TC ;
always_comb read_req_SAF_TC  = f_IsMEMRd(req_opcode) && addr_decode_SAF_TC ;

always_comb we_SAF_TC = {8{write_req_SAF_TC}} & be;
always_comb re_SAF_TC = {8{read_req_SAF_TC}} & be;
always_comb handcode_reg_wdata_SAF_TC = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_RX_VOQ_MAP_MEM) 
           {44'h0,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_RX_VOQ_PORT_CFG;
                    ack.read_miss = handcode_error_RX_VOQ_PORT_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h0,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_SAF_INGRESS_SPEED;
                    ack.read_miss = handcode_error_SAF_INGRESS_SPEED;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'b1???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_SAF_EGRESS_SPEED;
                    ack.read_miss = handcode_error_SAF_EGRESS_SPEED;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h10,4'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_SAF_TC;
                    ack.read_miss = handcode_error_SAF_TC;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_RX_VOQ_MAP_MEM) 
           {44'h0,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_RX_VOQ_PORT_CFG;
                    ack.write_miss = handcode_error_RX_VOQ_PORT_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h0,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_SAF_INGRESS_SPEED;
                    ack.write_miss = handcode_error_SAF_INGRESS_SPEED;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'b1???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_SAF_EGRESS_SPEED;
                    ack.write_miss = handcode_error_SAF_EGRESS_SPEED;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h10,4'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_SAF_TC;
                    ack.write_miss = handcode_error_SAF_TC;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_RX_VOQ_MAP_MEM) 
           {44'h0,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: read_data = handcode_reg_rdata_RX_VOQ_PORT_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'h0,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: read_data = handcode_reg_rdata_SAF_INGRESS_SPEED;
                 default: read_data = '0;
              endcase
           end
           {40'b1???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: read_data = handcode_reg_rdata_SAF_EGRESS_SPEED;
                 default: read_data = '0;
              endcase
           end
           {40'h10,4'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {RX_VOQ_SB_FID,RX_VOQ_SB_BAR}: read_data = handcode_reg_rdata_SAF_TC;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {


// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
