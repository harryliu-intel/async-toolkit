magic
tech scmos
timestamp 970031125
<< ndiffusion >>
rect -24 81 -8 82
rect -24 73 -8 78
rect -24 65 -8 70
rect -24 57 -8 62
rect -24 49 -8 54
rect -24 41 -8 46
rect -24 37 -8 38
rect -24 28 -8 29
<< pdiffusion >>
rect 14 91 40 92
rect 14 87 40 88
rect 28 79 40 87
rect 14 78 40 79
rect 14 74 40 75
rect 14 65 40 66
rect 14 61 40 62
rect 28 53 40 61
rect 14 52 40 53
rect 14 48 40 49
rect 14 39 40 40
rect 14 35 40 36
rect 14 24 30 27
rect 14 20 30 21
<< ntransistor >>
rect -24 78 -8 81
rect -24 70 -8 73
rect -24 62 -8 65
rect -24 54 -8 57
rect -24 46 -8 49
rect -24 38 -8 41
<< ptransistor >>
rect 14 88 40 91
rect 14 75 40 78
rect 14 62 40 65
rect 14 49 40 52
rect 14 36 40 39
rect 14 21 30 24
<< polysilicon >>
rect -6 88 14 91
rect 40 88 44 91
rect -6 81 -3 88
rect -28 78 -24 81
rect -8 78 -3 81
rect 9 75 14 78
rect 40 75 44 78
rect 9 73 12 75
rect -28 70 -24 73
rect -8 70 12 73
rect -28 62 -24 65
rect -8 62 14 65
rect 40 62 44 65
rect -28 54 -24 57
rect -8 54 12 57
rect 9 52 12 54
rect 9 49 14 52
rect 40 49 44 52
rect -33 46 -24 49
rect -8 46 4 49
rect -31 38 -24 41
rect -8 38 -4 41
rect 1 39 4 46
rect -31 20 -28 38
rect 1 36 14 39
rect 40 36 44 39
rect 10 21 14 24
rect 30 21 37 24
rect 34 20 37 21
<< ndcontact >>
rect -24 82 -8 90
rect -24 29 -8 37
<< pdcontact >>
rect 14 92 40 100
rect 14 79 28 87
rect 14 66 40 74
rect 14 53 28 61
rect 14 40 40 48
rect 14 27 40 35
rect 14 12 30 20
<< psubstratepcontact >>
rect -24 20 -8 28
<< nsubstratencontact >>
rect 49 88 57 96
<< polycontact >>
rect -36 78 -28 86
rect 44 73 52 81
rect -41 46 -33 54
rect 44 60 52 68
rect 44 47 52 55
rect -36 12 -28 20
rect 34 12 42 20
<< metal1 >>
rect 21 96 40 100
rect 14 92 57 96
rect -36 78 -28 84
rect -24 87 7 90
rect 32 88 57 92
rect -24 82 28 87
rect -1 79 28 82
rect -1 61 7 79
rect 32 74 40 88
rect 14 66 40 74
rect 44 78 52 81
rect -41 42 -33 54
rect -1 53 28 61
rect -24 20 -8 37
rect -1 35 7 53
rect 32 48 40 66
rect 44 66 52 68
rect 14 40 40 48
rect 44 54 52 55
rect 44 47 52 48
rect -1 30 40 35
rect 7 27 40 30
rect -36 18 -28 20
rect -21 18 -8 20
rect 14 18 30 20
rect 21 12 30 18
rect 34 18 42 20
<< m2contact >>
rect 3 96 21 102
rect -36 84 -28 90
rect 44 72 52 78
rect -41 36 -33 42
rect 44 60 52 66
rect 44 48 52 54
rect -1 24 7 30
rect -36 12 -28 18
rect -21 12 -3 18
rect 3 12 21 18
rect 34 12 42 18
<< metal2 >>
rect -36 84 0 90
rect 0 72 52 78
rect 0 60 52 66
rect 0 48 52 54
rect -41 36 0 42
rect -3 24 9 30
rect -37 12 -26 18
rect 31 12 42 18
<< m3contact >>
rect 3 96 21 102
rect -21 12 -3 18
rect 3 12 21 18
<< metal3 >>
rect -21 9 -3 105
rect 3 9 21 105
<< labels >>
rlabel polysilicon 31 22 31 22 1 _PReset!
rlabel metal1 18 31 18 31 1 x
rlabel metal1 18 44 18 44 5 Vdd!
rlabel metal1 18 57 18 57 5 x
rlabel metal1 18 70 18 70 1 Vdd!
rlabel metal1 18 83 18 83 1 x
rlabel metal1 18 96 18 96 5 Vdd!
rlabel metal1 -12 33 -12 33 1 GND!
rlabel metal1 -12 86 -12 86 1 x
rlabel polysilicon 41 37 41 37 3 a
rlabel polysilicon 41 50 41 50 3 b
rlabel polysilicon 41 63 41 63 3 c
rlabel polysilicon 41 76 41 76 3 d
rlabel polysilicon 41 89 41 89 3 e
rlabel metal2 38 15 38 15 1 _PReset!
rlabel polysilicon -25 47 -25 47 3 a
rlabel polysilicon -25 79 -25 79 3 e
rlabel polysilicon -25 71 -25 71 3 d
rlabel polysilicon -25 63 -25 63 3 c
rlabel polysilicon -25 55 -25 55 3 b
rlabel polysilicon -25 39 -25 39 3 _SReset!
rlabel m2contact 15 16 15 16 1 Vdd!
rlabel metal2 -32 15 -32 15 3 _SReset!
rlabel metal2 -26 12 -26 18 3 ^n
rlabel metal2 0 24 0 30 1 x
rlabel metal2 0 36 0 42 7 a
rlabel metal2 0 48 0 54 3 b
rlabel metal2 0 60 0 66 3 c
rlabel metal2 0 72 0 78 3 d
rlabel metal2 0 84 0 90 3 e
rlabel space -42 11 -24 91 7 ^n
rlabel metal1 53 92 53 92 7 Vdd!
rlabel space 28 31 58 101 3 ^p
rlabel metal2 -32 87 -32 87 1 e
rlabel metal2 -37 39 -37 39 3 a
rlabel metal2 48 51 48 51 1 b
rlabel metal2 48 63 48 63 1 c
rlabel metal2 48 75 48 75 1 d
<< end >>
