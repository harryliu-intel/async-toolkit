magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect -211 -724 -203 -723
rect -211 -732 -203 -727
rect -211 -740 -203 -735
rect -211 -748 -203 -743
rect -211 -756 -203 -751
rect -211 -760 -203 -759
rect -211 -769 -203 -768
rect -211 -777 -203 -772
rect -211 -785 -203 -780
rect -211 -793 -203 -788
rect -211 -801 -203 -796
rect -211 -805 -203 -804
<< pdiffusion >>
rect -181 -704 -157 -703
rect -181 -708 -157 -707
rect -173 -713 -157 -708
rect -181 -717 -173 -716
rect -181 -721 -173 -720
rect -181 -730 -173 -729
rect -181 -734 -173 -733
rect -181 -743 -173 -742
rect -181 -747 -173 -746
rect -181 -756 -173 -755
rect -181 -760 -173 -759
rect -181 -769 -173 -768
rect -181 -773 -173 -772
rect -181 -782 -173 -781
rect -181 -786 -173 -785
rect -181 -795 -173 -794
rect -181 -799 -173 -798
rect -181 -808 -173 -807
rect -181 -812 -173 -811
<< ntransistor >>
rect -211 -727 -203 -724
rect -211 -735 -203 -732
rect -211 -743 -203 -740
rect -211 -751 -203 -748
rect -211 -759 -203 -756
rect -211 -772 -203 -769
rect -211 -780 -203 -777
rect -211 -788 -203 -785
rect -211 -796 -203 -793
rect -211 -804 -203 -801
<< ptransistor >>
rect -181 -707 -157 -704
rect -181 -720 -173 -717
rect -181 -733 -173 -730
rect -181 -746 -173 -743
rect -181 -759 -173 -756
rect -181 -772 -173 -769
rect -181 -785 -173 -782
rect -181 -798 -173 -795
rect -181 -811 -173 -808
<< polysilicon >>
rect -185 -707 -181 -704
rect -157 -707 -153 -704
rect -186 -720 -181 -717
rect -173 -720 -169 -717
rect -215 -727 -211 -724
rect -203 -727 -199 -724
rect -186 -730 -183 -720
rect -186 -732 -181 -730
rect -215 -735 -211 -732
rect -203 -733 -181 -732
rect -173 -733 -169 -730
rect -203 -735 -183 -733
rect -215 -743 -211 -740
rect -203 -743 -183 -740
rect -186 -746 -181 -743
rect -173 -746 -169 -743
rect -215 -751 -211 -748
rect -203 -751 -191 -748
rect -194 -756 -191 -751
rect -215 -759 -211 -756
rect -203 -759 -199 -756
rect -194 -759 -181 -756
rect -173 -759 -169 -756
rect -215 -772 -211 -769
rect -203 -772 -199 -769
rect -194 -772 -181 -769
rect -173 -772 -169 -769
rect -194 -777 -191 -772
rect -215 -780 -211 -777
rect -203 -780 -191 -777
rect -186 -785 -181 -782
rect -173 -785 -169 -782
rect -215 -788 -211 -785
rect -203 -788 -183 -785
rect -215 -796 -211 -793
rect -203 -795 -183 -793
rect -203 -796 -181 -795
rect -186 -798 -181 -796
rect -173 -798 -169 -795
rect -215 -804 -211 -801
rect -203 -804 -199 -801
rect -186 -808 -183 -798
rect -186 -811 -181 -808
rect -173 -811 -169 -808
<< ndcontact >>
rect -211 -723 -203 -715
rect -211 -768 -203 -760
rect -211 -813 -203 -805
<< pdcontact >>
rect -181 -703 -157 -695
rect -181 -716 -173 -708
rect -181 -729 -173 -721
rect -181 -742 -173 -734
rect -181 -755 -173 -747
rect -181 -768 -173 -760
rect -181 -781 -173 -773
rect -181 -794 -173 -786
rect -181 -807 -173 -799
rect -181 -820 -173 -812
<< metal1 >>
rect -193 -703 -157 -695
rect -211 -723 -203 -715
rect -193 -721 -185 -703
rect -181 -716 -173 -708
rect -193 -729 -173 -721
rect -193 -747 -185 -729
rect -181 -742 -173 -734
rect -193 -755 -173 -747
rect -193 -760 -185 -755
rect -211 -768 -185 -760
rect -181 -768 -173 -760
rect -193 -773 -185 -768
rect -193 -781 -173 -773
rect -193 -799 -185 -781
rect -181 -794 -173 -786
rect -211 -813 -203 -805
rect -193 -807 -173 -799
rect -181 -820 -173 -812
<< labels >>
rlabel metal1 -177 -750 -177 -750 1 x
rlabel metal1 -177 -816 -177 -816 1 Vdd!
rlabel metal1 -177 -725 -177 -725 5 x
rlabel polysilicon -172 -810 -172 -810 7 a
rlabel polysilicon -172 -719 -172 -719 7 d
rlabel metal1 -177 -738 -177 -738 5 Vdd!
rlabel metal1 -177 -764 -177 -764 5 Vdd!
rlabel metal1 -177 -790 -177 -790 1 Vdd!
rlabel metal1 -177 -803 -177 -803 1 x
rlabel metal1 -177 -777 -177 -777 5 x
rlabel metal1 -177 -712 -177 -712 1 Vdd!
rlabel polysilicon -172 -784 -172 -784 7 b
rlabel polysilicon -172 -732 -172 -732 7 d
rlabel polysilicon -172 -797 -172 -797 7 a
rlabel polysilicon -172 -771 -172 -771 7 c
rlabel polysilicon -172 -758 -172 -758 7 b
rlabel polysilicon -172 -745 -172 -745 7 c
rlabel metal1 -177 -699 -177 -699 5 x
rlabel space -173 -820 -168 -715 3 ^p
rlabel polysilicon -156 -706 -156 -706 7 _PReset!
rlabel polysilicon -212 -758 -212 -758 3 a
rlabel polysilicon -212 -750 -212 -750 3 b
rlabel polysilicon -212 -742 -212 -742 3 c
rlabel metal1 -207 -764 -207 -764 5 x
rlabel polysilicon -212 -734 -212 -734 1 d
rlabel polysilicon -212 -787 -212 -787 3 b
rlabel polysilicon -212 -795 -212 -795 3 a
rlabel polysilicon -212 -779 -212 -779 1 c
rlabel polysilicon -212 -726 -212 -726 1 _SReset!
rlabel metal1 -207 -719 -207 -719 5 GND!
rlabel metal1 -207 -809 -207 -809 1 GND!
rlabel polysilicon -212 -803 -212 -803 1 _SReset!
rlabel polysilicon -212 -771 -212 -771 1 d
rlabel space -216 -813 -211 -715 7 ^n
<< end >>
