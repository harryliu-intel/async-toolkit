magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 192 642 202 643
rect 192 639 202 640
rect 192 635 194 639
rect 192 634 202 635
rect 192 631 202 632
rect 196 627 202 631
rect 192 626 202 627
rect 192 623 202 624
rect 192 619 194 623
rect 192 618 202 619
rect 192 615 202 616
rect 196 611 202 615
rect 192 610 202 611
rect 192 607 202 608
rect 192 603 194 607
rect 192 602 202 603
rect 192 599 202 600
rect 196 595 202 599
rect 192 594 202 595
rect 192 591 202 592
rect 192 587 194 591
rect 192 586 202 587
rect 192 583 202 584
<< pdiffusion >>
rect 214 638 220 639
rect 214 632 220 636
rect 214 629 220 630
rect 218 625 220 629
rect 214 624 220 625
rect 214 618 220 622
rect 214 615 220 616
rect 214 610 220 611
rect 214 604 220 608
rect 214 601 220 602
rect 218 597 220 601
rect 214 596 220 597
rect 214 590 220 594
rect 214 587 220 588
<< ntransistor >>
rect 192 640 202 642
rect 192 632 202 634
rect 192 624 202 626
rect 192 616 202 618
rect 192 608 202 610
rect 192 600 202 602
rect 192 592 202 594
rect 192 584 202 586
<< ptransistor >>
rect 214 636 220 638
rect 214 630 220 632
rect 214 622 220 624
rect 214 616 220 618
rect 214 608 220 610
rect 214 602 220 604
rect 214 594 220 596
rect 214 588 220 590
<< polysilicon >>
rect 189 640 192 642
rect 202 640 212 642
rect 210 638 212 640
rect 210 636 214 638
rect 220 636 223 638
rect 189 632 192 634
rect 202 632 206 634
rect 204 630 214 632
rect 220 630 223 632
rect 189 624 192 626
rect 202 624 206 626
rect 204 622 214 624
rect 220 622 223 624
rect 189 616 192 618
rect 202 616 214 618
rect 220 616 223 618
rect 189 608 192 610
rect 202 608 214 610
rect 220 608 223 610
rect 204 602 214 604
rect 220 602 223 604
rect 189 600 192 602
rect 202 600 206 602
rect 204 594 214 596
rect 220 594 223 596
rect 189 592 192 594
rect 202 592 206 594
rect 210 588 214 590
rect 220 588 223 590
rect 210 586 212 588
rect 189 584 192 586
rect 202 584 212 586
<< ndcontact >>
rect 192 643 202 647
rect 194 635 202 639
rect 192 627 196 631
rect 194 619 202 623
rect 192 611 196 615
rect 194 603 202 607
rect 192 595 196 599
rect 194 587 202 591
rect 192 579 202 583
<< pdcontact >>
rect 214 639 220 643
rect 214 625 218 629
rect 214 611 220 615
rect 214 597 218 601
rect 214 583 220 587
<< metal1 >>
rect 192 643 202 647
rect 214 639 220 643
rect 194 635 202 639
rect 192 627 196 631
rect 199 629 202 635
rect 199 625 218 629
rect 199 623 202 625
rect 194 619 202 623
rect 192 611 196 615
rect 199 607 202 619
rect 214 611 220 615
rect 194 603 202 607
rect 199 601 202 603
rect 192 595 196 599
rect 199 597 218 601
rect 199 591 202 597
rect 194 587 202 591
rect 214 583 220 587
rect 192 579 202 583
<< labels >>
rlabel polysilicon 221 603 221 603 7 a
rlabel polysilicon 221 609 221 609 7 b
rlabel polysilicon 221 589 221 589 7 a
rlabel polysilicon 221 595 221 595 7 b
rlabel polysilicon 221 623 221 623 7 b
rlabel polysilicon 221 617 221 617 7 a
rlabel polysilicon 221 637 221 637 7 b
rlabel polysilicon 221 631 221 631 7 a
rlabel polysilicon 191 641 191 641 7 b
rlabel polysilicon 191 625 191 625 7 b
rlabel polysilicon 191 609 191 609 7 b
rlabel polysilicon 191 593 191 593 7 b
rlabel polysilicon 191 585 191 585 7 a
rlabel polysilicon 191 601 191 601 7 a
rlabel polysilicon 191 617 191 617 7 a
rlabel polysilicon 191 633 191 633 7 a
rlabel space 188 579 192 647 7 ^n
rlabel space 220 583 224 643 3 ^p
rlabel pdcontact 216 627 216 627 1 x
rlabel pdcontact 216 599 216 599 1 x
rlabel ndcontact 200 589 200 589 1 x
rlabel ndcontact 200 605 200 605 1 x
rlabel ndcontact 200 621 200 621 1 x
rlabel ndcontact 200 637 200 637 1 x
rlabel ndcontact 197 581 197 581 1 GND!
rlabel ndcontact 194 597 194 597 3 GND!
rlabel ndcontact 194 613 194 613 3 GND!
rlabel ndcontact 194 629 194 629 3 GND!
rlabel ndcontact 197 645 197 645 5 GND!
rlabel pdcontact 216 641 216 641 1 Vdd!
rlabel pdcontact 216 613 216 613 1 Vdd!
rlabel pdcontact 216 585 216 585 1 Vdd!
<< end >>
