// This file created only for purposes of satisfying sla_pkg dependency when creating subsystem corekits.  Is NOT used during model compile/elab
// Should be removed once sla_pkg dependency is removed
`ifndef _SLA_PKG_
`define _SLA_PKG_
package sla_pkg;
endpackage: sla_pkg
`endif

