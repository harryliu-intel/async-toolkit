// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
// ---------------------------------------------------------------------------------------------------------------------
// -- Author : Edward C. Ross <edward.c.ross@intel.com>
// -- Project Name : Madison Bay (MBY)
// -- Description  : PB data memory interface 
// ---------------------------------------------------------------------------------------------------------------------

// This is a connectivity only interface and thus is just a named bundle of nets that can be passed around as a group 
// to save typing.  Anywhere an interface is defined, individual nets in the interface can be referenced as follows:    
//
//      <interface name>.<net name>
//


interface mby_igr_pb_d_if ();

    logic                                   wr_en;
    logic                                   rd_en;
    logic[mby_igr_pkg::PB_BANK_ADRS-1:0]    adr;
    logic[mby_igr_pkg::PB_SHELL_DATA_W-1:0] wr_data;
    logic                                   rd_valid;
    logic[mby_igr_pkg::PB_SHELL_DATA_W-1:0] rd_data;

    modport mem (
       input  wr_en,
       input  rd_en,
       input  adr,
       input  wr_data,
       output rd_valid,
       output rd_data
    );

    modport rtl (
       output wr_en,
       output rd_en,
       output adr,
       output wr_data,
       input  rd_valid,
       input  rd_data
    );

endinterface // mby_igr_pb_d_if
