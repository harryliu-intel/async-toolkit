magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect -205 -739 -197 -738
rect -205 -747 -197 -742
rect -205 -755 -197 -750
rect -205 -763 -197 -758
rect -205 -771 -197 -766
rect -205 -779 -197 -774
rect -205 -783 -197 -782
rect -205 -792 -197 -791
rect -205 -800 -197 -795
rect -205 -808 -197 -803
rect -205 -816 -197 -811
rect -205 -824 -197 -819
rect -205 -832 -197 -827
rect -205 -836 -197 -835
<< pdiffusion >>
rect -174 -714 -150 -713
rect -174 -718 -150 -717
rect -166 -723 -150 -718
rect -174 -727 -166 -726
rect -174 -731 -166 -730
rect -174 -740 -166 -739
rect -174 -744 -166 -743
rect -174 -753 -166 -752
rect -174 -757 -166 -756
rect -174 -766 -166 -765
rect -174 -770 -166 -769
rect -174 -779 -166 -778
rect -174 -783 -166 -782
rect -174 -792 -166 -791
rect -174 -796 -166 -795
rect -174 -805 -166 -804
rect -174 -809 -166 -808
rect -174 -818 -166 -817
rect -174 -822 -166 -821
rect -174 -831 -166 -830
rect -174 -835 -166 -834
rect -174 -844 -166 -843
rect -174 -848 -166 -847
<< ntransistor >>
rect -205 -742 -197 -739
rect -205 -750 -197 -747
rect -205 -758 -197 -755
rect -205 -766 -197 -763
rect -205 -774 -197 -771
rect -205 -782 -197 -779
rect -205 -795 -197 -792
rect -205 -803 -197 -800
rect -205 -811 -197 -808
rect -205 -819 -197 -816
rect -205 -827 -197 -824
rect -205 -835 -197 -832
<< ptransistor >>
rect -174 -717 -150 -714
rect -174 -730 -166 -727
rect -174 -743 -166 -740
rect -174 -756 -166 -753
rect -174 -769 -166 -766
rect -174 -782 -166 -779
rect -174 -795 -166 -792
rect -174 -808 -166 -805
rect -174 -821 -166 -818
rect -174 -834 -166 -831
rect -174 -847 -166 -844
<< polysilicon >>
rect -178 -717 -174 -714
rect -150 -717 -146 -714
rect -188 -730 -174 -727
rect -166 -730 -162 -727
rect -209 -742 -205 -739
rect -197 -742 -193 -739
rect -188 -747 -185 -730
rect -209 -750 -205 -747
rect -197 -750 -185 -747
rect -179 -743 -174 -740
rect -166 -743 -162 -740
rect -179 -753 -176 -743
rect -179 -755 -174 -753
rect -209 -758 -205 -755
rect -197 -756 -174 -755
rect -166 -756 -162 -753
rect -197 -758 -176 -756
rect -209 -766 -205 -763
rect -197 -766 -176 -763
rect -179 -769 -174 -766
rect -166 -769 -162 -766
rect -209 -774 -205 -771
rect -197 -774 -193 -771
rect -209 -782 -205 -779
rect -197 -782 -174 -779
rect -166 -782 -162 -779
rect -209 -795 -205 -792
rect -197 -795 -174 -792
rect -166 -795 -162 -792
rect -209 -803 -205 -800
rect -197 -803 -193 -800
rect -179 -808 -174 -805
rect -166 -808 -162 -805
rect -209 -811 -205 -808
rect -197 -811 -176 -808
rect -209 -819 -205 -816
rect -197 -818 -176 -816
rect -197 -819 -174 -818
rect -179 -821 -174 -819
rect -166 -821 -162 -818
rect -209 -827 -205 -824
rect -197 -827 -185 -824
rect -209 -835 -205 -832
rect -197 -835 -193 -832
rect -188 -844 -185 -827
rect -179 -831 -176 -821
rect -179 -834 -174 -831
rect -166 -834 -162 -831
rect -188 -847 -174 -844
rect -166 -847 -162 -844
<< ndcontact >>
rect -205 -738 -197 -730
rect -205 -791 -197 -783
rect -205 -844 -197 -836
<< pdcontact >>
rect -174 -713 -150 -705
rect -174 -726 -166 -718
rect -174 -739 -166 -731
rect -174 -752 -166 -744
rect -174 -765 -166 -757
rect -174 -778 -166 -770
rect -174 -791 -166 -783
rect -174 -804 -166 -796
rect -174 -817 -166 -809
rect -174 -830 -166 -822
rect -174 -843 -166 -835
rect -174 -856 -166 -848
<< metal1 >>
rect -186 -713 -150 -705
rect -205 -738 -197 -730
rect -186 -731 -178 -713
rect -174 -726 -166 -718
rect -186 -739 -166 -731
rect -186 -757 -178 -739
rect -174 -752 -166 -744
rect -186 -765 -166 -757
rect -186 -783 -178 -765
rect -174 -778 -166 -770
rect -205 -791 -166 -783
rect -186 -809 -178 -791
rect -174 -804 -166 -796
rect -186 -817 -166 -809
rect -186 -835 -178 -817
rect -174 -830 -166 -822
rect -205 -844 -197 -836
rect -186 -843 -166 -835
rect -174 -856 -166 -848
<< labels >>
rlabel metal1 -170 -773 -170 -773 5 Vdd!
rlabel metal1 -170 -799 -170 -799 5 Vdd!
rlabel metal1 -170 -852 -170 -852 1 Vdd!
rlabel metal1 -170 -761 -170 -761 5 x
rlabel metal1 -170 -723 -170 -723 1 Vdd!
rlabel metal1 -170 -735 -170 -735 5 x
rlabel metal1 -170 -748 -170 -748 1 Vdd!
rlabel metal1 -170 -787 -170 -787 1 x
rlabel metal1 -170 -813 -170 -813 5 x
rlabel metal1 -170 -839 -170 -839 1 x
rlabel metal1 -170 -826 -170 -826 1 Vdd!
rlabel polysilicon -165 -729 -165 -729 7 e
rlabel polysilicon -165 -794 -165 -794 7 e
rlabel polysilicon -165 -846 -165 -846 7 a
rlabel polysilicon -165 -781 -165 -781 7 a
rlabel polysilicon -165 -768 -165 -768 7 c
rlabel polysilicon -165 -807 -165 -807 7 c
rlabel polysilicon -165 -833 -165 -833 7 b
rlabel polysilicon -165 -820 -165 -820 7 b
rlabel polysilicon -165 -755 -165 -755 7 d
rlabel polysilicon -165 -742 -165 -742 7 d
rlabel metal1 -170 -709 -170 -709 5 x
rlabel polysilicon -206 -781 -206 -781 3 a
rlabel polysilicon -206 -773 -206 -773 3 b
rlabel polysilicon -206 -765 -206 -765 3 c
rlabel metal1 -201 -787 -201 -787 5 x
rlabel polysilicon -206 -757 -206 -757 1 d
rlabel polysilicon -206 -810 -206 -810 3 c
rlabel polysilicon -206 -818 -206 -818 3 b
rlabel polysilicon -206 -826 -206 -826 3 a
rlabel polysilicon -206 -802 -206 -802 1 d
rlabel polysilicon -206 -794 -206 -794 3 e
rlabel polysilicon -206 -749 -206 -749 3 e
rlabel metal1 -201 -733 -201 -733 5 GND!
rlabel polysilicon -207 -741 -207 -741 1 _SReset!
rlabel polysilicon -206 -834 -206 -834 1 _SReset!
rlabel metal1 -201 -840 -201 -840 1 GND!
rlabel space -210 -844 -205 -730 7 ^n
rlabel space -166 -856 -161 -725 3 ^p
rlabel polysilicon -149 -716 -149 -716 7 _PReset!
<< end >>
