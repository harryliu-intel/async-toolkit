magic
tech scmos
timestamp 965153727
<< ndiffusion >>
rect 57 77 83 78
rect 57 73 83 74
rect 57 65 69 73
rect 57 64 83 65
rect 57 60 83 61
rect 71 52 83 60
rect 57 51 83 52
rect 57 47 83 48
rect 57 39 69 47
rect 57 38 83 39
rect 57 34 83 35
rect 71 26 83 34
rect 57 25 83 26
rect 57 21 83 22
rect 57 13 69 21
rect 57 12 83 13
rect 57 8 83 9
<< pdiffusion >>
rect 99 77 125 78
rect 99 73 125 74
rect 113 65 125 73
rect 99 64 125 65
rect 99 60 125 61
rect 99 52 111 60
rect 99 51 125 52
rect 99 47 125 48
rect 113 39 125 47
rect 99 38 125 39
rect 99 34 125 35
rect 99 26 111 34
rect 99 25 125 26
rect 99 21 125 22
rect 113 13 125 21
rect 99 12 125 13
rect 99 8 125 9
<< ntransistor >>
rect 57 74 83 77
rect 57 61 83 64
rect 57 48 83 51
rect 57 35 83 38
rect 57 22 83 25
rect 57 9 83 12
<< ptransistor >>
rect 99 74 125 77
rect 99 61 125 64
rect 99 48 125 51
rect 99 35 125 38
rect 99 22 125 25
rect 99 9 125 12
<< polysilicon >>
rect 53 74 57 77
rect 83 74 99 77
rect 125 74 129 77
rect 87 64 95 74
rect 53 61 57 64
rect 83 61 99 64
rect 125 61 129 64
rect 87 51 95 61
rect 53 48 57 51
rect 83 49 99 51
rect 83 48 87 49
rect 53 35 57 38
rect 83 35 87 38
rect 53 22 57 25
rect 83 22 87 25
rect 53 9 57 12
rect 83 9 87 12
rect 95 48 99 49
rect 125 48 129 51
rect 95 35 99 38
rect 125 35 129 38
rect 95 22 99 25
rect 125 22 129 25
rect 95 9 99 12
rect 125 9 129 12
<< ndcontact >>
rect 57 78 83 86
rect 69 65 83 73
rect 57 52 71 60
rect 69 39 83 47
rect 57 26 71 34
rect 69 13 83 21
rect 57 0 83 8
<< pdcontact >>
rect 99 78 125 86
rect 99 65 113 73
rect 111 52 125 60
rect 99 39 113 47
rect 111 26 125 34
rect 99 13 113 21
rect 99 0 125 8
<< polycontact >>
rect 87 9 95 49
<< metal1 >>
rect 57 78 83 86
rect 99 78 125 86
rect 57 60 65 78
rect 69 65 113 73
rect 57 52 71 60
rect 75 53 107 65
rect 117 60 125 78
rect 57 34 65 52
rect 75 47 83 53
rect 69 39 83 47
rect 57 26 71 34
rect 57 8 65 26
rect 75 21 83 39
rect 69 13 83 21
rect 87 9 95 49
rect 99 47 107 53
rect 111 52 125 60
rect 99 39 113 47
rect 99 21 107 39
rect 117 34 125 52
rect 111 26 125 34
rect 99 13 113 21
rect 117 8 125 26
rect 57 0 83 8
rect 99 0 125 8
<< labels >>
rlabel ndcontact 75 43 75 43 1 x
rlabel ndcontact 75 17 75 17 1 x
rlabel ndcontact 75 69 75 69 1 x
rlabel ndcontact 65 30 65 30 5 GND!
rlabel ndcontact 65 56 65 56 5 GND!
rlabel ndcontact 65 82 65 82 5 GND!
rlabel ndcontact 65 4 65 4 1 GND!
rlabel space 52 -1 70 87 7 ^n
rlabel pdcontact 107 43 107 43 1 x
rlabel pdcontact 107 17 107 17 1 x
rlabel pdcontact 107 69 107 69 1 x
rlabel pdcontact 117 4 117 4 1 Vdd!
rlabel pdcontact 117 30 117 30 5 Vdd!
rlabel pdcontact 117 56 117 56 5 Vdd!
rlabel pdcontact 117 82 117 82 5 Vdd!
rlabel space 112 -1 130 87 3 ^p
rlabel metal1 91 29 91 29 1 a
<< end >>
