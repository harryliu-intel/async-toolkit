magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect -15 90 -7 91
rect -15 82 -7 87
rect -15 74 -7 79
rect -15 66 -7 71
rect -15 58 -7 63
rect -15 50 -7 55
rect -15 46 -7 47
<< pdiffusion >>
rect 15 100 23 101
rect 15 96 23 97
rect 15 87 23 88
rect 15 83 23 84
rect 15 74 23 75
rect 15 70 23 71
rect 15 61 23 62
rect 15 57 23 58
rect 15 48 23 49
rect 15 44 23 45
rect 23 36 31 41
rect 15 35 31 36
rect 15 31 31 32
<< ntransistor >>
rect -15 87 -7 90
rect -15 79 -7 82
rect -15 71 -7 74
rect -15 63 -7 66
rect -15 55 -7 58
rect -15 47 -7 50
<< ptransistor >>
rect 15 97 23 100
rect 15 84 23 87
rect 15 71 23 74
rect 15 58 23 61
rect 15 45 23 48
rect 15 32 31 35
<< polysilicon >>
rect -5 97 15 100
rect 23 97 27 100
rect -5 90 -2 97
rect -19 87 -15 90
rect -7 87 -2 90
rect 10 84 15 87
rect 23 84 27 87
rect 10 82 13 84
rect -19 79 -15 82
rect -7 79 13 82
rect -19 71 -15 74
rect -7 71 15 74
rect 23 71 27 74
rect -19 63 -15 66
rect -7 63 13 66
rect 10 61 13 63
rect 10 58 15 61
rect 23 58 27 61
rect -19 55 -15 58
rect -7 55 5 58
rect -19 47 -15 50
rect -7 47 -3 50
rect 2 48 5 55
rect 2 45 15 48
rect 23 45 27 48
rect 11 32 15 35
rect 31 32 35 35
<< ndcontact >>
rect -15 91 -7 99
rect -15 38 -7 46
<< pdcontact >>
rect 15 101 23 109
rect 15 88 23 96
rect 15 75 23 83
rect 15 62 23 70
rect 15 49 23 57
rect 15 36 23 44
rect 15 23 31 31
<< metal1 >>
rect 15 101 23 109
rect -15 96 11 99
rect -15 91 23 96
rect 3 88 23 91
rect 3 70 11 88
rect 15 75 23 83
rect 3 62 23 70
rect -15 38 -7 46
rect 3 44 11 62
rect 15 49 23 57
rect 3 36 23 44
rect 15 23 31 31
<< labels >>
rlabel metal1 19 40 19 40 1 x
rlabel metal1 19 53 19 53 5 Vdd!
rlabel metal1 19 66 19 66 5 x
rlabel metal1 19 79 19 79 1 Vdd!
rlabel metal1 19 92 19 92 1 x
rlabel metal1 19 105 19 105 5 Vdd!
rlabel polysilicon 24 46 24 46 3 a
rlabel polysilicon 24 59 24 59 3 b
rlabel polysilicon 24 72 24 72 3 c
rlabel polysilicon 24 85 24 85 3 d
rlabel polysilicon 24 98 24 98 3 e
rlabel metal1 19 27 19 27 1 Vdd!
rlabel metal1 -11 42 -11 42 1 GND!
rlabel metal1 -11 95 -11 95 1 x
rlabel polysilicon -16 48 -16 48 3 _SReset!
rlabel polysilicon -16 64 -16 64 3 b
rlabel polysilicon -16 72 -16 72 3 c
rlabel polysilicon -16 80 -16 80 3 d
rlabel polysilicon -16 88 -16 88 3 e
rlabel polysilicon -16 56 -16 56 3 a
rlabel space -20 38 -15 99 7 ^n
rlabel polysilicon 32 33 32 33 1 _PReset!
rlabel space 23 43 28 109 3 ^p
<< end >>
