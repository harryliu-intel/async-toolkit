// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Raghu P Gudla
// Created On   :  09/22/2018
// Description  :  CHI request node directed basic sequence. provides initiator 
//                 scenario information to the RN agent present in the system env.
//                 this class defines a sequence in which a CHI WRITENOSNPFULL seq
//                 is generated by assigning values to the transactions rather than 
//                 randomization, and then transmitted using `uvm_send.
// -------------------------------------------------------------------------------------------------------------

class fc_chi_rn_basic_seq extends svt_chi_rn_transaction_base_sequence;

  /** node configuration obtained from the sequencer */
  svt_chi_node_configuration cfg;

  /** parameter that controls the number of transactions that will be generated */
  rand int unsigned sequence_length;

  /** constrain the sequence length to a reasonable value*/ 
  constraint reasonable_sequence_length {
    sequence_length inside {1};
  }

  /** UVM object utility macro */
  `uvm_object_utils(fc_chi_rn_basic_seq)

    /** class constructor */
  function new(string name="fc_chi_rn_basic_seq");
    super.new(name);
  endfunction

  virtual task body();
    svt_chi_rn_transaction write_tran, read_tran;
    svt_configuration get_cfg;
    bit status;
    int txn_id = 0;

    `uvm_info("body", "entered ...", UVM_LOW)
    
    p_sequencer.get_cfg(get_cfg);
    if (!$cast(cfg, get_cfg)) begin
      `uvm_fatal("body", "unable to $cast the configuration to a svt_chi_port_configuration class");
    end
    /** 
     * this method is defined in the svt_chi_rn_transaction_base_sequence.
     * it obtains the virtual sequencer rn_virt_seqr of type svt_chi_rn_virtual_sequencer 
     * from the configuration database and sets up the shared resources obtained from it: the response_request_port.
     * 
     **/
    get_rn_virt_seqr();

    super.body();

    /** gets the user provided sequence_length. */
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
    `uvm_info("body", $sformatf("sequence_length is %0d as a result of %0s.", sequence_length, status ? "config DB" : "randomization"), UVM_LOW);
    
    for(int i=0; i<sequence_length; i++) begin
      
      /** set up the write transaction */
      `uvm_create(write_tran)
      write_tran.cfg = this.cfg;
      write_tran.txn_id = txn_id++;
      write_tran.data_size = svt_chi_rn_transaction::SIZE_64BYTE;
      write_tran.addr         = 64'h0001_0000_0100_0010;
      
      if (i%2) begin
        write_tran.xact_type    = svt_chi_rn_transaction::WRITENOSNPFULL;
      end
      else begin
        write_tran.xact_type = svt_chi_rn_transaction::WRITENOSNPPTL;
      end
      
      for (int j=0; j<8; j++)
        write_tran.data[64*j+:64] = 64'hdead_beef_feed_beef;

      if(write_tran.xact_type  == svt_chi_rn_transaction::WRITENOSNPFULL) 
        write_tran.byte_enable = {`SVT_CHI_MAX_BE_WIDTH{1'b1}};
      else 
        write_tran.byte_enable = $urandom_range((write_tran.power_of_2(`SVT_CHI_DAT_FLIT_MAX_BE_WIDTH)-1), 1);
      
      write_tran.exp_comp_ack = 1'b0;
      write_tran.is_likely_shared = 1'b0;
      write_tran.snp_attr_is_snoopable = 1'b0;
      write_tran.snp_attr_snp_domain_type = svt_chi_transaction::INNER;
      write_tran.mem_attr_is_early_wr_ack_allowed = 1'b1;
      write_tran.mem_attr_mem_type = svt_chi_transaction::NORMAL;

      // construct dat_rsvdc to accomodate for the number of tx DAT
      // flits associated to this transaction and then setup the values.
      write_tran.dat_rsvdc = new[write_tran.compute_num_dat_flits()];
      foreach (write_tran.dat_rsvdc[idx])
        write_tran.dat_rsvdc[idx] = (idx+1);

      // adjust byte_enable field to make sure that the generated byte_enable
      // doesn't violate the protocol.
      write_tran.post_randomize();
      
      `uvm_info("body", $sformatf("sending CHI WRITE transaction %0s", `SVT_CHI_PRINT_PREFIX(write_tran)), UVM_LOW);      
      /** send the write transaction */
      `uvm_send(write_tran);
      /** wait for the write transaction to complete */
      get_response(rsp);
      `uvm_info("body", $sformatf("sending CHI WRITE transaction %0s completed", `SVT_CHI_PRINT_PREFIX(write_tran)), UVM_LOW)

       /** set up the read transaction */
      `uvm_create(read_tran)
      read_tran.cfg = this.cfg;
      read_tran.txn_id = txn_id++;
      read_tran.data_size = svt_chi_transaction::SIZE_64BYTE;
      read_tran.xact_type    = svt_chi_transaction::READNOSNP;
      read_tran.addr         = write_tran.addr; // 44'h001_0000_0100 | ('h100 << i)
      read_tran.byte_enable = write_tran.byte_enable;
      read_tran.exp_comp_ack = 1'b1;
      read_tran.is_likely_shared = 1'b0;
      read_tran.snp_attr_is_snoopable = 1'b0;
      read_tran.snp_attr_snp_domain_type = svt_chi_transaction::INNER;
      read_tran.mem_attr_is_early_wr_ack_allowed = 1'b1;
      read_tran.mem_attr_mem_type = svt_chi_transaction::NORMAL;

     `uvm_info("body", $sformatf("sending CHI READ transaction %0s", `SVT_CHI_PRINT_PREFIX(read_tran)), UVM_LOW);
      /** send the read transaction */
      `uvm_send(read_tran)
      /** wait for the read transaction to complete */
      get_response(rsp);
      `uvm_info("body", $sformatf("CHI READ transaction %0s completed", `SVT_CHI_PRINT_PREFIX(read_tran)), UVM_LOW);
    end

    `uvm_info("body", "exiting...", UVM_LOW)
  endtask: body

endclass: fc_chi_rn_basic_seq

