magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -220 -719 -214 -718
rect -220 -725 -214 -721
rect -220 -731 -214 -727
rect -220 -737 -214 -733
rect -220 -743 -214 -739
rect -220 -746 -214 -745
rect -220 -750 -218 -746
rect -220 -751 -214 -750
rect -220 -757 -214 -753
rect -220 -763 -214 -759
rect -220 -769 -214 -765
rect -220 -775 -214 -771
rect -220 -778 -214 -777
<< pdiffusion >>
rect -199 -711 -189 -710
rect -199 -714 -189 -713
rect -191 -718 -189 -714
rect -199 -719 -189 -718
rect -199 -722 -189 -721
rect -199 -726 -193 -722
rect -199 -727 -189 -726
rect -199 -730 -189 -729
rect -191 -734 -189 -730
rect -199 -735 -189 -734
rect -199 -738 -189 -737
rect -199 -742 -193 -738
rect -199 -743 -189 -742
rect -199 -746 -189 -745
rect -191 -750 -189 -746
rect -199 -751 -189 -750
rect -199 -754 -189 -753
rect -199 -758 -193 -754
rect -199 -759 -189 -758
rect -199 -762 -189 -761
rect -191 -766 -189 -762
rect -199 -767 -189 -766
rect -199 -770 -189 -769
rect -199 -774 -193 -770
rect -199 -775 -189 -774
rect -199 -778 -189 -777
rect -191 -782 -189 -778
rect -199 -783 -189 -782
rect -199 -786 -189 -785
<< ntransistor >>
rect -220 -721 -214 -719
rect -220 -727 -214 -725
rect -220 -733 -214 -731
rect -220 -739 -214 -737
rect -220 -745 -214 -743
rect -220 -753 -214 -751
rect -220 -759 -214 -757
rect -220 -765 -214 -763
rect -220 -771 -214 -769
rect -220 -777 -214 -775
<< ptransistor >>
rect -199 -713 -189 -711
rect -199 -721 -189 -719
rect -199 -729 -189 -727
rect -199 -737 -189 -735
rect -199 -745 -189 -743
rect -199 -753 -189 -751
rect -199 -761 -189 -759
rect -199 -769 -189 -767
rect -199 -777 -189 -775
rect -199 -785 -189 -783
<< polysilicon >>
rect -208 -713 -199 -711
rect -189 -713 -186 -711
rect -208 -719 -206 -713
rect -223 -721 -220 -719
rect -214 -721 -206 -719
rect -203 -721 -199 -719
rect -189 -721 -186 -719
rect -203 -725 -201 -721
rect -223 -727 -220 -725
rect -214 -727 -201 -725
rect -203 -729 -199 -727
rect -189 -729 -186 -727
rect -223 -733 -220 -731
rect -214 -733 -206 -731
rect -208 -735 -206 -733
rect -208 -737 -199 -735
rect -189 -737 -186 -735
rect -223 -739 -220 -737
rect -214 -739 -211 -737
rect -223 -745 -220 -743
rect -214 -745 -199 -743
rect -189 -745 -186 -743
rect -223 -753 -220 -751
rect -214 -753 -199 -751
rect -189 -753 -186 -751
rect -223 -759 -220 -757
rect -214 -759 -211 -757
rect -208 -761 -199 -759
rect -189 -761 -186 -759
rect -208 -763 -206 -761
rect -223 -765 -220 -763
rect -214 -765 -206 -763
rect -203 -769 -199 -767
rect -189 -769 -186 -767
rect -223 -771 -220 -769
rect -214 -771 -201 -769
rect -203 -775 -201 -771
rect -223 -777 -220 -775
rect -214 -777 -206 -775
rect -203 -777 -199 -775
rect -189 -777 -186 -775
rect -208 -783 -206 -777
rect -208 -785 -199 -783
rect -189 -785 -186 -783
<< ndcontact >>
rect -220 -718 -214 -714
rect -218 -750 -214 -746
rect -220 -782 -214 -778
<< pdcontact >>
rect -199 -710 -189 -706
rect -199 -718 -191 -714
rect -193 -726 -189 -722
rect -199 -734 -191 -730
rect -193 -742 -189 -738
rect -199 -750 -191 -746
rect -193 -758 -189 -754
rect -199 -766 -191 -762
rect -193 -774 -189 -770
rect -199 -782 -191 -778
rect -199 -790 -189 -786
<< metal1 >>
rect -199 -710 -189 -706
rect -220 -718 -214 -714
rect -199 -718 -191 -714
rect -199 -730 -196 -718
rect -193 -726 -189 -722
rect -199 -734 -191 -730
rect -199 -746 -196 -734
rect -193 -742 -189 -738
rect -218 -750 -191 -746
rect -199 -762 -196 -750
rect -193 -758 -189 -754
rect -199 -766 -191 -762
rect -199 -778 -196 -766
rect -193 -774 -189 -770
rect -220 -782 -214 -778
rect -199 -782 -191 -778
rect -199 -790 -189 -786
<< labels >>
rlabel polysilicon -188 -712 -188 -712 3 e
rlabel polysilicon -188 -720 -188 -720 3 d
rlabel polysilicon -188 -728 -188 -728 3 d
rlabel polysilicon -188 -736 -188 -736 3 c
rlabel polysilicon -188 -744 -188 -744 3 a
rlabel polysilicon -188 -752 -188 -752 3 e
rlabel polysilicon -188 -760 -188 -760 3 c
rlabel polysilicon -188 -768 -188 -768 3 b
rlabel polysilicon -188 -776 -188 -776 3 b
rlabel polysilicon -188 -784 -188 -784 3 a
rlabel space -192 -791 -186 -705 3 ^p
rlabel polysilicon -221 -776 -221 -776 3 a
rlabel polysilicon -221 -770 -221 -770 3 b
rlabel polysilicon -221 -764 -221 -764 3 c
rlabel polysilicon -221 -758 -221 -758 3 d
rlabel polysilicon -221 -744 -221 -744 3 a
rlabel polysilicon -221 -738 -221 -738 3 b
rlabel polysilicon -221 -732 -221 -732 3 c
rlabel polysilicon -221 -726 -221 -726 3 d
rlabel polysilicon -221 -720 -221 -720 3 e
rlabel polysilicon -221 -752 -221 -752 3 e
rlabel space -223 -783 -217 -713 7 ^n
rlabel pdcontact -191 -740 -191 -740 1 Vdd!
rlabel pdcontact -191 -724 -191 -724 1 Vdd!
rlabel pdcontact -191 -756 -191 -756 1 Vdd!
rlabel pdcontact -191 -772 -191 -772 1 Vdd!
rlabel pdcontact -191 -788 -191 -788 1 Vdd!
rlabel pdcontact -191 -708 -191 -708 1 Vdd!
rlabel pdcontact -197 -716 -197 -716 1 x
rlabel pdcontact -197 -732 -197 -732 1 x
rlabel pdcontact -197 -748 -197 -748 1 x
rlabel pdcontact -197 -764 -197 -764 1 x
rlabel pdcontact -197 -780 -197 -780 1 x
rlabel ndcontact -216 -748 -216 -748 1 x
rlabel ndcontact -216 -716 -216 -716 5 GND!
rlabel ndcontact -216 -780 -216 -780 1 GND!
<< end >>
