magic
tech scmos
timestamp 962798985
<< ndiffusion >>
rect -85 1 -77 2
rect -63 -2 -55 -1
rect -85 -7 -77 -2
rect -85 -15 -77 -10
rect -63 -6 -55 -5
rect -63 -15 -55 -14
rect -85 -19 -77 -18
rect -63 -19 -55 -18
<< pdiffusion >>
rect -138 14 -130 19
rect -138 13 -122 14
rect -138 7 -122 10
rect -138 4 -132 7
rect -124 4 -122 7
rect -132 -2 -124 -1
rect -132 -6 -124 -5
rect -39 -2 -31 -1
rect -111 -12 -107 -9
rect -132 -15 -124 -14
rect -132 -19 -124 -18
rect -111 -19 -107 -16
rect -39 -6 -31 -5
rect -39 -15 -31 -14
rect -39 -19 -31 -18
<< ntransistor >>
rect -85 -2 -77 1
rect -63 -5 -55 -2
rect -85 -10 -77 -7
rect -85 -18 -77 -15
rect -63 -18 -55 -15
<< ptransistor >>
rect -138 10 -122 13
rect -132 -5 -124 -2
rect -39 -5 -31 -2
rect -132 -18 -124 -15
rect -111 -16 -107 -12
rect -39 -18 -31 -15
<< polysilicon >>
rect -142 10 -138 13
rect -122 10 -118 13
rect -120 1 -87 4
rect -67 6 -65 9
rect -120 -2 -117 1
rect -137 -5 -132 -2
rect -124 -5 -117 -2
rect -137 -15 -134 -5
rect -90 -2 -85 1
rect -77 -2 -73 1
rect -68 -2 -65 6
rect -68 -5 -63 -2
rect -55 -5 -39 -2
rect -31 -5 -27 -2
rect -98 -10 -85 -7
rect -77 -10 -73 -7
rect -137 -18 -132 -15
rect -124 -18 -120 -15
rect -115 -16 -111 -12
rect -107 -16 -103 -12
rect -68 -15 -65 -5
rect -89 -18 -85 -15
rect -77 -18 -73 -15
rect -68 -18 -63 -15
rect -55 -18 -39 -15
rect -31 -18 -27 -15
<< ndcontact >>
rect -85 2 -77 10
rect -63 -1 -55 7
rect -63 -14 -55 -6
rect -85 -27 -77 -19
rect -63 -27 -55 -19
<< pdcontact >>
rect -130 14 -122 22
rect -132 -1 -124 7
rect -132 -14 -124 -6
rect -115 -9 -107 -1
rect -39 -1 -31 7
rect -39 -14 -31 -6
rect -132 -27 -124 -19
rect -115 -27 -107 -19
rect -39 -27 -31 -19
<< polycontact >>
rect -75 6 -67 14
rect -103 -18 -95 -10
<< metal1 >>
rect -130 18 -122 22
rect -130 14 -116 18
rect -132 -1 -124 7
rect -120 -1 -116 14
rect -75 10 -67 14
rect -85 5 -67 10
rect -85 2 -77 5
rect -85 -1 -80 2
rect -63 -1 -55 7
rect -39 -1 -31 7
rect -120 -6 -80 -1
rect -132 -9 -107 -6
rect -132 -11 -116 -9
rect -63 -10 -31 -6
rect -132 -14 -124 -11
rect -103 -14 -31 -10
rect -103 -18 -95 -14
rect -132 -27 -107 -19
rect -85 -27 -55 -19
rect -39 -27 -31 -19
<< labels >>
rlabel metal1 -111 -23 -111 -23 1 Vdd!
rlabel polysilicon -112 -15 -112 -15 1 x
rlabel metal1 -111 -5 -111 -5 1 _x
rlabel polysilicon -133 -4 -133 -4 1 a
rlabel polysilicon -133 -17 -133 -17 1 a
rlabel metal1 -128 3 -128 3 5 Vdd!
rlabel metal1 -128 -23 -128 -23 1 Vdd!
rlabel metal1 -128 -10 -128 -10 1 _x
rlabel metal1 -126 18 -126 18 1 _x
rlabel polysilicon -139 11 -139 11 3 _PReset!
rlabel space -138 -27 -132 1 7 ^p1
rlabel metal1 -81 6 -81 6 1 _x
rlabel polysilicon -86 -17 -86 -17 1 _SReset!
rlabel polysilicon -86 -9 -86 -9 1 x
rlabel polysilicon -86 -1 -86 -1 1 a
rlabel metal1 -81 -23 -81 -23 1 GND!
rlabel polysilicon -64 -4 -64 -4 3 _x
rlabel polysilicon -64 -17 -64 -17 3 _x
rlabel ndcontact -59 3 -59 3 5 GND!
rlabel ndcontact -59 -23 -59 -23 1 GND!
rlabel ndcontact -59 -10 -59 -10 1 x
rlabel polysilicon -30 -17 -30 -17 1 _x
rlabel polysilicon -30 -4 -30 -4 1 _x
rlabel pdcontact -35 3 -35 3 5 Vdd!
rlabel pdcontact -35 -10 -35 -10 1 x
rlabel pdcontact -35 -23 -35 -23 1 Vdd!
rlabel space -31 -27 -26 7 3 ^p2
rlabel space -55 -28 -25 8 3 ^n2
<< end >>
