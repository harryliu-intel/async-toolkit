magic
tech scmos
timestamp 970030488
<< ndiffusion >>
rect -24 104 -8 105
rect -24 96 -8 101
rect -24 88 -8 93
rect -24 84 -8 85
<< pdiffusion >>
rect 8 109 34 110
rect 8 105 34 106
rect 22 97 34 105
rect 8 96 34 97
rect 8 92 34 93
rect 8 81 34 84
rect 8 77 34 78
rect 16 72 34 77
<< ntransistor >>
rect -24 101 -8 104
rect -24 93 -8 96
rect -24 85 -8 88
<< ptransistor >>
rect 8 106 34 109
rect 8 93 34 96
rect 8 78 34 81
<< polysilicon >>
rect -4 106 8 109
rect 34 106 38 109
rect -4 104 -1 106
rect -28 101 -24 104
rect -8 101 -1 104
rect -28 93 -24 96
rect -8 93 8 96
rect 34 93 38 96
rect -31 85 -24 88
rect -8 85 -4 88
rect -31 77 -28 85
rect 4 78 8 81
rect 34 78 41 81
rect 38 77 41 78
<< ndcontact >>
rect -24 105 -8 113
rect -24 76 -8 84
<< pdcontact >>
rect 8 110 34 118
rect 8 97 22 105
rect 8 84 34 92
rect 8 69 16 77
<< psubstratepcontact >>
rect -41 84 -33 92
<< nsubstratencontact >>
rect 43 110 51 118
<< polycontact >>
rect -36 101 -28 109
rect 38 93 46 101
rect -36 69 -28 77
rect 38 69 46 77
<< metal1 >>
rect 21 117 51 118
rect -24 105 -8 113
rect 8 110 51 117
rect -36 101 -28 105
rect -14 103 -8 105
rect 8 103 22 105
rect -14 97 22 103
rect -41 84 -16 92
rect -4 87 4 97
rect 26 92 34 110
rect 38 99 46 101
rect -36 75 -28 77
rect -24 76 -8 84
rect -21 75 -8 76
rect 8 84 34 92
rect -4 77 4 81
rect -4 69 16 77
rect 38 75 46 77
<< m2contact >>
rect 3 117 21 123
rect -36 105 -28 111
rect 38 93 46 99
rect -36 69 -28 75
rect -21 69 -8 75
rect -4 81 4 87
rect 38 69 46 75
<< metal2 >>
rect -36 105 0 111
rect 0 93 46 99
rect -6 81 6 87
rect -37 69 -26 75
rect 27 69 46 75
<< m3contact >>
rect 3 117 21 123
rect -21 69 -8 75
<< metal3 >>
rect -21 66 -3 126
rect 3 66 21 126
<< labels >>
rlabel polysilicon -25 86 -25 86 3 _SReset!
rlabel polysilicon -25 102 -25 102 3 b
rlabel polysilicon -25 94 -25 94 3 a
rlabel metal1 12 101 12 101 1 x
rlabel metal1 12 114 12 114 5 Vdd!
rlabel metal1 12 88 12 88 1 Vdd!
rlabel metal1 -12 80 -12 80 1 GND!
rlabel metal1 -12 109 -12 109 1 x
rlabel metal1 12 73 12 73 1 x
rlabel polysilicon 35 107 35 107 1 b
rlabel polysilicon 35 94 35 94 1 a
rlabel polysilicon 35 79 35 79 1 _PReset!
rlabel metal2 0 93 0 99 3 a
rlabel metal2 0 105 0 111 7 b
rlabel metal2 42 72 42 72 1 _PReset!
rlabel metal2 -31 72 -31 72 1 _SReset!
rlabel metal2 -26 69 -26 75 3 ^n
rlabel metal2 0 81 0 87 1 x
rlabel metal1 47 114 47 114 7 Vdd!
rlabel space 22 88 52 119 3 ^p
rlabel metal1 -37 88 -37 88 3 GND!
rlabel space -42 68 -23 114 7 ^n
rlabel metal2 -32 108 -32 108 1 b
rlabel metal2 42 96 42 96 1 a
<< end >>
