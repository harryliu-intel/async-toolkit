magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 6 96 10 97
rect 43 100 46 102
rect 43 94 46 98
rect 6 90 10 94
rect 6 87 10 88
rect 43 87 46 89
rect 42 82 46 83
rect 42 79 46 80
<< pdiffusion >>
rect 60 100 63 102
rect 22 96 26 97
rect 60 96 63 98
rect 22 90 26 94
rect 58 91 66 92
rect 22 87 26 88
rect 58 88 66 89
rect 58 85 60 88
rect 64 85 66 88
rect 60 82 64 83
rect 60 79 64 80
<< ntransistor >>
rect 43 98 46 100
rect 6 94 10 96
rect 6 88 10 90
rect 43 89 46 94
rect 42 80 46 82
<< ptransistor >>
rect 60 98 63 100
rect 22 94 26 96
rect 22 88 26 90
rect 58 89 66 91
rect 60 80 64 82
<< polysilicon >>
rect 40 98 43 100
rect 46 98 60 100
rect 63 98 74 100
rect 3 94 6 96
rect 10 94 22 96
rect 26 94 29 96
rect 3 88 6 90
rect 10 88 22 90
rect 26 88 29 90
rect 40 89 43 94
rect 46 91 49 94
rect 46 89 58 91
rect 66 89 69 91
rect 39 80 42 82
rect 46 81 52 82
rect 56 81 60 82
rect 46 80 60 81
rect 64 80 67 82
rect 72 79 74 98
<< ndcontact >>
rect 42 102 46 106
rect 6 97 10 101
rect 6 83 10 87
rect 42 83 46 87
rect 42 75 46 79
<< pdcontact >>
rect 22 97 26 101
rect 60 102 64 106
rect 58 92 66 96
rect 22 83 26 87
rect 60 83 64 88
rect 60 75 64 79
<< polycontact >>
rect 52 81 56 85
rect 71 75 75 79
<< metal1 >>
rect 42 105 46 106
rect 42 102 56 105
rect 60 102 64 106
rect 6 97 26 101
rect 53 96 56 102
rect 53 92 66 96
rect 6 83 10 87
rect 22 83 26 87
rect 42 83 46 87
rect 53 85 56 92
rect 52 81 56 85
rect 60 83 64 88
rect 42 78 46 79
rect 60 78 64 79
rect 71 78 75 79
rect 42 75 75 78
<< labels >>
rlabel polysilicon 5 89 5 89 3 a
rlabel polysilicon 5 95 5 95 3 b
rlabel space 2 82 6 102 7 ^n
rlabel space 26 82 30 102 3 ^p
rlabel polysilicon 27 89 27 89 3 a
rlabel polysilicon 27 95 27 95 3 b
rlabel polysilicon 42 90 42 90 1 _PReset!
rlabel ndcontact 8 99 8 99 1 x
rlabel ndcontact 8 85 8 85 1 GND!
rlabel pdcontact 24 99 24 99 1 x
rlabel pdcontact 24 85 24 85 1 Vdd!
rlabel pdcontact 62 85 62 85 1 Vdd!
rlabel ndcontact 44 85 44 85 1 GND!
rlabel pdcontact 62 94 62 94 1 x
rlabel pdcontact 62 104 62 104 1 Vdd!
rlabel ndcontact 44 104 44 104 5 x
<< end >>
