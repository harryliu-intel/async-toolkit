magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 10 45 14 46
rect 10 39 14 43
rect 10 33 14 37
rect 10 27 14 31
rect 10 21 14 25
rect 10 18 14 19
<< pdiffusion >>
rect 34 50 36 54
rect 26 49 36 50
rect 26 46 36 47
rect 26 42 32 46
rect 26 41 36 42
rect 26 38 36 39
rect 34 34 36 38
rect 26 33 36 34
rect 26 30 36 31
rect 26 26 32 30
rect 26 25 36 26
rect 26 22 36 23
rect 34 18 36 22
rect 26 17 36 18
rect 26 14 36 15
<< ntransistor >>
rect 10 43 14 45
rect 10 37 14 39
rect 10 31 14 33
rect 10 25 14 27
rect 10 19 14 21
<< ptransistor >>
rect 26 47 36 49
rect 26 39 36 41
rect 26 31 36 33
rect 26 23 36 25
rect 26 15 36 17
<< polysilicon >>
rect 16 47 26 49
rect 36 47 39 49
rect 16 45 18 47
rect 7 43 10 45
rect 14 43 18 45
rect 22 39 26 41
rect 36 39 39 41
rect 7 37 10 39
rect 14 37 24 39
rect 7 31 10 33
rect 14 31 26 33
rect 36 31 39 33
rect 7 25 10 27
rect 14 25 24 27
rect 22 23 26 25
rect 36 23 39 25
rect 7 19 10 21
rect 14 19 18 21
rect 16 17 18 19
rect 16 15 26 17
rect 36 15 39 17
<< ndcontact >>
rect 10 46 14 50
rect 10 14 14 18
<< pdcontact >>
rect 26 50 34 54
rect 32 42 36 46
rect 26 34 34 38
rect 32 26 36 30
rect 26 18 34 22
rect 26 10 36 14
<< metal1 >>
rect 26 50 34 54
rect 10 46 29 50
rect 26 38 29 46
rect 32 42 36 46
rect 26 34 34 38
rect 26 22 29 34
rect 32 26 36 30
rect 26 18 34 22
rect 10 14 14 18
rect 26 10 36 14
<< labels >>
rlabel polysilicon 9 38 9 38 3 d
rlabel polysilicon 9 32 9 32 3 c
rlabel polysilicon 9 26 9 26 3 b
rlabel polysilicon 9 20 9 20 3 a
rlabel polysilicon 9 44 9 44 3 e
rlabel space 33 9 39 55 3 ^p
rlabel polysilicon 37 48 37 48 7 e
rlabel polysilicon 37 40 37 40 3 d
rlabel polysilicon 37 16 37 16 3 a
rlabel polysilicon 37 24 37 24 3 b
rlabel polysilicon 37 32 37 32 3 c
rlabel space 7 14 10 50 7 ^n
rlabel ndcontact 12 48 12 48 4 x
rlabel ndcontact 12 16 12 16 5 GND!
rlabel pdcontact 34 28 34 28 1 Vdd!
rlabel pdcontact 34 44 34 44 5 Vdd!
rlabel pdcontact 30 36 30 36 5 x
rlabel pdcontact 30 20 30 20 5 x
rlabel pdcontact 30 52 30 52 5 x
rlabel pdcontact 34 12 34 12 1 Vdd!
<< end >>
