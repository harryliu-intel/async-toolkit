// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

///
///  INTEL CONFIDENTIAL
///
///  Copyright 2019 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_tx_pb_pkg.vh                                           
// Creator:         ggomezde                                                   
// Time:            Wednesday Jan 30, 2019 [10:29:56 am]                       
//                                                                             
// Path:            /tmp/ggomezde/nebulon_run/2289325233_2019-01-30.10:29:27   
// Arguments:       -I                                                         
//                  /nfs/site/disks/sc_mby_00088/ggomezde/mby/work_root/models/mby_ww05_ral_TI/tools/srdl
//                  -sv_no_sai_checks -sverilog -crif -expand_handcoded_arrays 
//                  -maximize_crif -input mby_tx_pb_map.rdl -timeout 60000     
//                  -out_dir /tmp/tmp.0b1MJL16ua -log_file                     
//                  /nfs/site/disks/sc_mby_00088/ggomezde/mby/work_root/models/mby_ww05_ral_TI/target/GenRTL/regflow/mby/subblock/mby_tx_pb_map_crif.xml.log
//                                                                             
// MRE:             5.2018.3.p1                                                
// Machine:         sccj004303                                                 
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww52.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2019 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtlgen_pkg_template

`ifndef MBY_TX_PB_PKG_VH
`define MBY_TX_PB_PKG_VH

`include "rtlgen_include_mby_tx_pb_map.vh"
`include "rtlgen_pkg_mby_tx_pb_map.vh"

package mby_tx_pb_pkg;

import rtlgen_pkg_mby_tx_pb_map::*;

typedef cfg_req_64bit_t mby_tx_pb_cr_req_t;
typedef cfg_ack_64bit_t mby_tx_pb_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_tx_pb_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [31:0] PORT;  // RW
} TX_PB_PORT_CFG_t;

localparam TX_PB_PORT_CFG_REG_STRIDE = 48'h8;
localparam TX_PB_PORT_CFG_REG_ENTRIES = 1;
localparam TX_PB_PORT_CFG_CR_ADDR = 48'h0;
localparam TX_PB_PORT_CFG_SIZE = 64;
localparam TX_PB_PORT_CFG_PORT_LO = 0;
localparam TX_PB_PORT_CFG_PORT_HI = 31;
localparam TX_PB_PORT_CFG_PORT_RESET = 'h0;
localparam TX_PB_PORT_CFG_USEMASK = 64'hFFFFFFFF;
localparam TX_PB_PORT_CFG_RO_MASK = 64'h0;
localparam TX_PB_PORT_CFG_WO_MASK = 64'h0;
localparam TX_PB_PORT_CFG_RESET = 64'h0;

typedef struct packed {
    logic [55:0] reserved0;  // RSVD
    logic  [7:0] BUF_SIZE;  // RW
} TX_PB_PREFETCH_t;

localparam TX_PB_PREFETCH_REG_STRIDE = 48'h8;
localparam TX_PB_PREFETCH_REG_ENTRIES = 16;
localparam TX_PB_PREFETCH_CR_ADDR = 48'h80;
localparam TX_PB_PREFETCH_SIZE = 64;
localparam TX_PB_PREFETCH_BUF_SIZE_LO = 0;
localparam TX_PB_PREFETCH_BUF_SIZE_HI = 7;
localparam TX_PB_PREFETCH_BUF_SIZE_RESET = 'h0;
localparam TX_PB_PREFETCH_USEMASK = 64'hFF;
localparam TX_PB_PREFETCH_RO_MASK = 64'h0;
localparam TX_PB_PREFETCH_WO_MASK = 64'h0;
localparam TX_PB_PREFETCH_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_TX_PB_PORT_CFG_t;

typedef logic [7:0] we_TX_PB_PREFETCH_t;

typedef struct packed {
    we_TX_PB_PORT_CFG_t TX_PB_PORT_CFG;
    we_TX_PB_PREFETCH_t TX_PB_PREFETCH;
} mby_tx_pb_handcoded_t;

typedef logic [7:0] re_TX_PB_PORT_CFG_t;

typedef logic [7:0] re_TX_PB_PREFETCH_t;

typedef struct packed {
    re_TX_PB_PORT_CFG_t TX_PB_PORT_CFG;
    re_TX_PB_PREFETCH_t TX_PB_PREFETCH;
} mby_tx_pb_hc_re_t;

typedef logic handcode_rvalid_TX_PB_PORT_CFG_t;

typedef logic handcode_rvalid_TX_PB_PREFETCH_t;

typedef struct packed {
    handcode_rvalid_TX_PB_PORT_CFG_t TX_PB_PORT_CFG;
    handcode_rvalid_TX_PB_PREFETCH_t TX_PB_PREFETCH;
} mby_tx_pb_hc_rvalid_t;

typedef logic handcode_wvalid_TX_PB_PORT_CFG_t;

typedef logic handcode_wvalid_TX_PB_PREFETCH_t;

typedef struct packed {
    handcode_wvalid_TX_PB_PORT_CFG_t TX_PB_PORT_CFG;
    handcode_wvalid_TX_PB_PREFETCH_t TX_PB_PREFETCH;
} mby_tx_pb_hc_wvalid_t;

typedef logic handcode_error_TX_PB_PORT_CFG_t;

typedef logic handcode_error_TX_PB_PREFETCH_t;

typedef struct packed {
    handcode_error_TX_PB_PORT_CFG_t TX_PB_PORT_CFG;
    handcode_error_TX_PB_PREFETCH_t TX_PB_PREFETCH;
} mby_tx_pb_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    TX_PB_PORT_CFG_t TX_PB_PORT_CFG;
    TX_PB_PREFETCH_t TX_PB_PREFETCH;
} mby_tx_pb_hc_reg_read_t;

typedef struct packed {
    TX_PB_PORT_CFG_t TX_PB_PORT_CFG;
    TX_PB_PREFETCH_t TX_PB_PREFETCH;
} mby_tx_pb_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Parity Bit Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_tx_pb_pkg

`endif // MBY_TX_PB_PKG_VH
