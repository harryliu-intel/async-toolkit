// vim: noai : ts=3 : sw=3 : expandtab : ft=systemverilog

//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors.  The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//   Author        : Nathan Mai
//                 : Lewis Sternberg
//   Project       : Madison Bay
//------------------------------------------------------------------------------

//   Defines : types useful to mby_rx_ppe testbench
//

`ifndef __MBY_RX_PPE_DEFINES_GUARD
`define __MBY_RX_PPE_DEFINES_GUARD

//FIXME:  LNS: `defines are global and should be avoided whenever possible. 
////            When it's not to avoid `defines, their name should be made unambiguously unique by using the prefix MBY_RX_PPE
`define NUM_VPS_PER_IGR   1
`define NUM_PORTS_PER_VP  8
`define NUM_EPLS_PER_RX_PPE 1
`define NUM_PORTS_PER_EPL 16

`ifndef __INSIDE_MBY_RX_PPE_ENV_PKG
`error "Attempt to include file outside of mby_rx_ppe_env_pkg."
`endif


`endif // __MBY_RX_PPE_DEFINES_GUARD
