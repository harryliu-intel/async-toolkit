///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_parser_map_pkg.vh                                  
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_PARSER_MAP_PKG_VH
`define MBY_PPE_PARSER_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_parser_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_parser_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_parser_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_parser_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic  [7:0] INITIAL_W0_OFFSET;  // RW
    logic  [7:0] INITIAL_W1_OFFSET;  // RW
    logic  [7:0] INITIAL_W2_OFFSET;  // RW
    logic  [7:0] INITIAL_PTR;  // RW
    logic [15:0] INITIAL_STATE;  // RW
    logic [11:0] INITIAL_OP_MASK;  // RW
    logic  [3:0] INITIAL_OP_ROT;  // RW
} PARSER_PORT_CFG_t;

localparam PARSER_PORT_CFG_REG_STRIDE = 48'h8;
localparam PARSER_PORT_CFG_REG_ENTRIES = 16;
localparam PARSER_PORT_CFG_CR_ADDR = 48'h0;
localparam PARSER_PORT_CFG_SIZE = 64;
localparam PARSER_PORT_CFG_INITIAL_W0_OFFSET_LO = 56;
localparam PARSER_PORT_CFG_INITIAL_W0_OFFSET_HI = 63;
localparam PARSER_PORT_CFG_INITIAL_W0_OFFSET_RESET = 8'h0;
localparam PARSER_PORT_CFG_INITIAL_W1_OFFSET_LO = 48;
localparam PARSER_PORT_CFG_INITIAL_W1_OFFSET_HI = 55;
localparam PARSER_PORT_CFG_INITIAL_W1_OFFSET_RESET = 8'h0;
localparam PARSER_PORT_CFG_INITIAL_W2_OFFSET_LO = 40;
localparam PARSER_PORT_CFG_INITIAL_W2_OFFSET_HI = 47;
localparam PARSER_PORT_CFG_INITIAL_W2_OFFSET_RESET = 8'h0;
localparam PARSER_PORT_CFG_INITIAL_PTR_LO = 32;
localparam PARSER_PORT_CFG_INITIAL_PTR_HI = 39;
localparam PARSER_PORT_CFG_INITIAL_PTR_RESET = 8'h0;
localparam PARSER_PORT_CFG_INITIAL_STATE_LO = 16;
localparam PARSER_PORT_CFG_INITIAL_STATE_HI = 31;
localparam PARSER_PORT_CFG_INITIAL_STATE_RESET = 16'h0;
localparam PARSER_PORT_CFG_INITIAL_OP_MASK_LO = 4;
localparam PARSER_PORT_CFG_INITIAL_OP_MASK_HI = 15;
localparam PARSER_PORT_CFG_INITIAL_OP_MASK_RESET = 12'h0;
localparam PARSER_PORT_CFG_INITIAL_OP_ROT_LO = 0;
localparam PARSER_PORT_CFG_INITIAL_OP_ROT_HI = 3;
localparam PARSER_PORT_CFG_INITIAL_OP_ROT_RESET = 4'h0;
localparam PARSER_PORT_CFG_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam PARSER_PORT_CFG_RO_MASK = 64'h0;
localparam PARSER_PORT_CFG_WO_MASK = 64'h0;
localparam PARSER_PORT_CFG_RESET = 64'h0;

typedef struct packed {
    logic [53:0] reserved0;  // RSVD
    logic  [0:0] VALIDATE_IPV4_HDR_CSUM;  // RW
    logic  [0:0] VALIDATE_IPV4_HDR_TRUNCATION;  // RW
    logic  [0:0] VALIDATE_IPV4_HDR_LENGTH;  // RW
    logic  [0:0] VALIDATE_IPV4_LENGTH;  // RW
    logic  [1:0] VALIDATE_L4_CSUM;  // RW
    logic  [0:0] STORE_L4_PARTIAL_CSUM;  // RW
    logic  [0:0] COMPUTE_L4_CSUM;  // RW
    logic  [1:0] VALIDATE_L3_LENGTH;  // RW
} PARSER_CSUM_CFG_t;

localparam PARSER_CSUM_CFG_REG_STRIDE = 48'h8;
localparam PARSER_CSUM_CFG_REG_ENTRIES = 16;
localparam PARSER_CSUM_CFG_CR_ADDR = 48'h80;
localparam PARSER_CSUM_CFG_SIZE = 64;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_CSUM_LO = 9;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_CSUM_HI = 9;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_CSUM_RESET = 1'h0;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_TRUNCATION_LO = 8;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_TRUNCATION_HI = 8;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_TRUNCATION_RESET = 1'h0;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_LENGTH_LO = 7;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_LENGTH_HI = 7;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_HDR_LENGTH_RESET = 1'h0;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_LENGTH_LO = 6;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_LENGTH_HI = 6;
localparam PARSER_CSUM_CFG_VALIDATE_IPV4_LENGTH_RESET = 1'h0;
localparam PARSER_CSUM_CFG_VALIDATE_L4_CSUM_LO = 4;
localparam PARSER_CSUM_CFG_VALIDATE_L4_CSUM_HI = 5;
localparam PARSER_CSUM_CFG_VALIDATE_L4_CSUM_RESET = 2'h0;
localparam PARSER_CSUM_CFG_STORE_L4_PARTIAL_CSUM_LO = 3;
localparam PARSER_CSUM_CFG_STORE_L4_PARTIAL_CSUM_HI = 3;
localparam PARSER_CSUM_CFG_STORE_L4_PARTIAL_CSUM_RESET = 1'h0;
localparam PARSER_CSUM_CFG_COMPUTE_L4_CSUM_LO = 2;
localparam PARSER_CSUM_CFG_COMPUTE_L4_CSUM_HI = 2;
localparam PARSER_CSUM_CFG_COMPUTE_L4_CSUM_RESET = 1'h0;
localparam PARSER_CSUM_CFG_VALIDATE_L3_LENGTH_LO = 0;
localparam PARSER_CSUM_CFG_VALIDATE_L3_LENGTH_HI = 1;
localparam PARSER_CSUM_CFG_VALIDATE_L3_LENGTH_RESET = 2'h0;
localparam PARSER_CSUM_CFG_USEMASK = 64'h3FF;
localparam PARSER_CSUM_CFG_RO_MASK = 64'h0;
localparam PARSER_CSUM_CFG_WO_MASK = 64'h0;
localparam PARSER_CSUM_CFG_RESET = 64'h0;

typedef struct packed {
    logic [62:0] reserved0;  // RSVD
    logic  [0:0] MEM_ERROR;  // RW/1C/V
} PARSER_IP_t;

localparam PARSER_IP_REG_STRIDE = 48'h8;
localparam PARSER_IP_REG_ENTRIES = 1;
localparam PARSER_IP_CR_ADDR = 48'h100;
localparam PARSER_IP_SIZE = 64;
localparam PARSER_IP_MEM_ERROR_LO = 0;
localparam PARSER_IP_MEM_ERROR_HI = 0;
localparam PARSER_IP_MEM_ERROR_RESET = 1'h0;
localparam PARSER_IP_USEMASK = 64'h1;
localparam PARSER_IP_RO_MASK = 64'h0;
localparam PARSER_IP_WO_MASK = 64'h0;
localparam PARSER_IP_RESET = 64'h0;

typedef struct packed {
    logic [62:0] reserved0;  // RSVD
    logic  [0:0] MEM_ERROR;  // RW
} PARSER_IM_t;

localparam PARSER_IM_REG_STRIDE = 48'h8;
localparam PARSER_IM_REG_ENTRIES = 1;
localparam PARSER_IM_CR_ADDR = 48'h108;
localparam PARSER_IM_SIZE = 64;
localparam PARSER_IM_MEM_ERROR_LO = 0;
localparam PARSER_IM_MEM_ERROR_HI = 0;
localparam PARSER_IM_MEM_ERROR_RESET = 1'h1;
localparam PARSER_IM_USEMASK = 64'h1;
localparam PARSER_IM_RO_MASK = 64'h0;
localparam PARSER_IM_WO_MASK = 64'h0;
localparam PARSER_IM_RESET = 64'h1;

typedef struct packed {
    logic [15:0] W1_VALUE;  // RW
    logic [15:0] W1_MASK;  // RW
    logic [15:0] W0_VALUE;  // RW
    logic [15:0] W0_MASK;  // RW
} PARSER_KEY_W_t;

localparam PARSER_KEY_W_REG_STRIDE = 48'h8;
localparam PARSER_KEY_W_REG_ENTRIES = 16;
localparam PARSER_KEY_W_REGFILE_STRIDE = 48'h80;
localparam PARSER_KEY_W_REGFILE_ENTRIES = 32;
localparam PARSER_KEY_W_CR_ADDR = 48'h1000;
localparam PARSER_KEY_W_SIZE = 64;
localparam PARSER_KEY_W_W1_VALUE_LO = 48;
localparam PARSER_KEY_W_W1_VALUE_HI = 63;
localparam PARSER_KEY_W_W1_VALUE_RESET = 16'hffff;
localparam PARSER_KEY_W_W1_MASK_LO = 32;
localparam PARSER_KEY_W_W1_MASK_HI = 47;
localparam PARSER_KEY_W_W1_MASK_RESET = 16'h0;
localparam PARSER_KEY_W_W0_VALUE_LO = 16;
localparam PARSER_KEY_W_W0_VALUE_HI = 31;
localparam PARSER_KEY_W_W0_VALUE_RESET = 16'hffff;
localparam PARSER_KEY_W_W0_MASK_LO = 0;
localparam PARSER_KEY_W_W0_MASK_HI = 15;
localparam PARSER_KEY_W_W0_MASK_RESET = 16'h0;
localparam PARSER_KEY_W_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam PARSER_KEY_W_RO_MASK = 64'h0;
localparam PARSER_KEY_W_WO_MASK = 64'h0;
localparam PARSER_KEY_W_RESET = 64'hFFFF0000FFFF0000;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [15:0] STATE_VALUE;  // RW
    logic [15:0] STATE_MASK;  // RW
} PARSER_KEY_S_t;

localparam PARSER_KEY_S_REG_STRIDE = 48'h8;
localparam PARSER_KEY_S_REG_ENTRIES = 16;
localparam PARSER_KEY_S_REGFILE_STRIDE = 48'h80;
localparam PARSER_KEY_S_REGFILE_ENTRIES = 32;
localparam PARSER_KEY_S_CR_ADDR = 48'h2000;
localparam PARSER_KEY_S_SIZE = 64;
localparam PARSER_KEY_S_STATE_VALUE_LO = 16;
localparam PARSER_KEY_S_STATE_VALUE_HI = 31;
localparam PARSER_KEY_S_STATE_VALUE_RESET = 16'hffff;
localparam PARSER_KEY_S_STATE_MASK_LO = 0;
localparam PARSER_KEY_S_STATE_MASK_HI = 15;
localparam PARSER_KEY_S_STATE_MASK_RESET = 16'h0;
localparam PARSER_KEY_S_USEMASK = 64'hFFFFFFFF;
localparam PARSER_KEY_S_RO_MASK = 64'h0;
localparam PARSER_KEY_S_WO_MASK = 64'h0;
localparam PARSER_KEY_S_RESET = 64'hFFFF0000;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic  [7:0] NEXT_W0_OFFSET;  // RW
    logic  [7:0] NEXT_W1_OFFSET;  // RW
    logic  [7:0] NEXT_W2_OFFSET;  // RW
    logic  [7:0] SKIP;  // RW
} PARSER_ANA_W_t;

localparam PARSER_ANA_W_REG_STRIDE = 48'h8;
localparam PARSER_ANA_W_REG_ENTRIES = 16;
localparam PARSER_ANA_W_REGFILE_STRIDE = 48'h80;
localparam PARSER_ANA_W_REGFILE_ENTRIES = 32;
localparam PARSER_ANA_W_CR_ADDR = 48'h3000;
localparam PARSER_ANA_W_SIZE = 64;
localparam PARSER_ANA_W_NEXT_W0_OFFSET_LO = 24;
localparam PARSER_ANA_W_NEXT_W0_OFFSET_HI = 31;
localparam PARSER_ANA_W_NEXT_W0_OFFSET_RESET = 8'h0;
localparam PARSER_ANA_W_NEXT_W1_OFFSET_LO = 16;
localparam PARSER_ANA_W_NEXT_W1_OFFSET_HI = 23;
localparam PARSER_ANA_W_NEXT_W1_OFFSET_RESET = 8'h0;
localparam PARSER_ANA_W_NEXT_W2_OFFSET_LO = 8;
localparam PARSER_ANA_W_NEXT_W2_OFFSET_HI = 15;
localparam PARSER_ANA_W_NEXT_W2_OFFSET_RESET = 8'h0;
localparam PARSER_ANA_W_SKIP_LO = 0;
localparam PARSER_ANA_W_SKIP_HI = 7;
localparam PARSER_ANA_W_SKIP_RESET = 8'h0;
localparam PARSER_ANA_W_USEMASK = 64'hFFFFFFFF;
localparam PARSER_ANA_W_RO_MASK = 64'h0;
localparam PARSER_ANA_W_WO_MASK = 64'h0;
localparam PARSER_ANA_W_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [15:0] NEXT_STATE;  // RW
    logic [15:0] NEXT_STATE_MASK;  // RW
    logic [15:0] NEXT_OP;  // RW
} PARSER_ANA_S_t;

localparam PARSER_ANA_S_REG_STRIDE = 48'h8;
localparam PARSER_ANA_S_REG_ENTRIES = 16;
localparam PARSER_ANA_S_REGFILE_STRIDE = 48'h80;
localparam PARSER_ANA_S_REGFILE_ENTRIES = 32;
localparam PARSER_ANA_S_CR_ADDR = 48'h4000;
localparam PARSER_ANA_S_SIZE = 64;
localparam PARSER_ANA_S_NEXT_STATE_LO = 32;
localparam PARSER_ANA_S_NEXT_STATE_HI = 47;
localparam PARSER_ANA_S_NEXT_STATE_RESET = 16'h0;
localparam PARSER_ANA_S_NEXT_STATE_MASK_LO = 16;
localparam PARSER_ANA_S_NEXT_STATE_MASK_HI = 31;
localparam PARSER_ANA_S_NEXT_STATE_MASK_RESET = 16'h0;
localparam PARSER_ANA_S_NEXT_OP_LO = 0;
localparam PARSER_ANA_S_NEXT_OP_HI = 15;
localparam PARSER_ANA_S_NEXT_OP_RESET = 16'h0;
localparam PARSER_ANA_S_USEMASK = 64'hFFFFFFFFFFFF;
localparam PARSER_ANA_S_RO_MASK = 64'h0;
localparam PARSER_ANA_S_WO_MASK = 64'h0;
localparam PARSER_ANA_S_RESET = 64'h0;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [7:0] EX_OFFSET;  // RW
    logic  [0:0] PARSING_DONE;  // RW
} PARSER_EXC_t;

localparam PARSER_EXC_REG_STRIDE = 48'h8;
localparam PARSER_EXC_REG_ENTRIES = 16;
localparam PARSER_EXC_REGFILE_STRIDE = 48'h80;
localparam PARSER_EXC_REGFILE_ENTRIES = 32;
localparam PARSER_EXC_CR_ADDR = 48'h5000;
localparam PARSER_EXC_SIZE = 64;
localparam PARSER_EXC_EX_OFFSET_LO = 1;
localparam PARSER_EXC_EX_OFFSET_HI = 8;
localparam PARSER_EXC_EX_OFFSET_RESET = 8'h0;
localparam PARSER_EXC_PARSING_DONE_LO = 0;
localparam PARSER_EXC_PARSING_DONE_HI = 0;
localparam PARSER_EXC_PARSING_DONE_RESET = 1'h0;
localparam PARSER_EXC_USEMASK = 64'h1FF;
localparam PARSER_EXC_RO_MASK = 64'h0;
localparam PARSER_EXC_WO_MASK = 64'h0;
localparam PARSER_EXC_RESET = 64'h0;

typedef struct packed {
    logic [37:0] reserved0;  // RSVD
    logic  [7:0] PROTOCOL_ID;  // RW
    logic  [7:0] OFFSET;  // RW
    logic  [5:0] FLAG_NUM;  // RW
    logic  [0:0] FLAG_VALUE;  // RW
    logic  [2:0] PTR_NUM;  // RW
} PARSER_EXT_t;

localparam PARSER_EXT_REG_STRIDE = 48'h8;
localparam PARSER_EXT_REG_ENTRIES = 32;
localparam PARSER_EXT_REGFILE_STRIDE = 48'h100;
localparam PARSER_EXT_REGFILE_ENTRIES = 32;
localparam PARSER_EXT_CR_ADDR = 48'h6000;
localparam PARSER_EXT_SIZE = 64;
localparam PARSER_EXT_PROTOCOL_ID_LO = 18;
localparam PARSER_EXT_PROTOCOL_ID_HI = 25;
localparam PARSER_EXT_PROTOCOL_ID_RESET = 8'hff;
localparam PARSER_EXT_OFFSET_LO = 10;
localparam PARSER_EXT_OFFSET_HI = 17;
localparam PARSER_EXT_OFFSET_RESET = 8'h0;
localparam PARSER_EXT_FLAG_NUM_LO = 4;
localparam PARSER_EXT_FLAG_NUM_HI = 9;
localparam PARSER_EXT_FLAG_NUM_RESET = 6'h0;
localparam PARSER_EXT_FLAG_VALUE_LO = 3;
localparam PARSER_EXT_FLAG_VALUE_HI = 3;
localparam PARSER_EXT_FLAG_VALUE_RESET = 1'h0;
localparam PARSER_EXT_PTR_NUM_LO = 0;
localparam PARSER_EXT_PTR_NUM_HI = 2;
localparam PARSER_EXT_PTR_NUM_RESET = 3'h0;
localparam PARSER_EXT_USEMASK = 64'h3FFFFFF;
localparam PARSER_EXT_RO_MASK = 64'h0;
localparam PARSER_EXT_WO_MASK = 64'h0;
localparam PARSER_EXT_RESET = 64'h3FC0000;

typedef struct packed {
    logic [31:0] KEY_INVERT;  // RW
    logic [31:0] KEY;  // RW
} PARSER_PTYPE_TCAM_t;

localparam PARSER_PTYPE_TCAM_REG_STRIDE = 48'h8;
localparam PARSER_PTYPE_TCAM_REG_ENTRIES = 64;
localparam PARSER_PTYPE_TCAM_REGFILE_STRIDE = 48'h200;
localparam PARSER_PTYPE_TCAM_REGFILE_ENTRIES = 2;
localparam PARSER_PTYPE_TCAM_CR_ADDR = 48'h8000;
localparam PARSER_PTYPE_TCAM_SIZE = 64;
localparam PARSER_PTYPE_TCAM_KEY_INVERT_LO = 32;
localparam PARSER_PTYPE_TCAM_KEY_INVERT_HI = 63;
localparam PARSER_PTYPE_TCAM_KEY_INVERT_RESET = 32'h0;
localparam PARSER_PTYPE_TCAM_KEY_LO = 0;
localparam PARSER_PTYPE_TCAM_KEY_HI = 31;
localparam PARSER_PTYPE_TCAM_KEY_RESET = 32'h0;
localparam PARSER_PTYPE_TCAM_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam PARSER_PTYPE_TCAM_RO_MASK = 64'h0;
localparam PARSER_PTYPE_TCAM_WO_MASK = 64'h0;
localparam PARSER_PTYPE_TCAM_RESET = 64'h0;

typedef struct packed {
    logic [49:0] reserved0;  // RSVD
    logic  [3:0] EXTRACT_IDX;  // RW
    logic  [9:0] PTYPE;  // RW
} PARSER_PTYPE_RAM_t;

localparam PARSER_PTYPE_RAM_REG_STRIDE = 48'h8;
localparam PARSER_PTYPE_RAM_REG_ENTRIES = 64;
localparam PARSER_PTYPE_RAM_REGFILE_STRIDE = 48'h200;
localparam PARSER_PTYPE_RAM_REGFILE_ENTRIES = 2;
localparam PARSER_PTYPE_RAM_CR_ADDR = 48'h8400;
localparam PARSER_PTYPE_RAM_SIZE = 64;
localparam PARSER_PTYPE_RAM_EXTRACT_IDX_LO = 10;
localparam PARSER_PTYPE_RAM_EXTRACT_IDX_HI = 13;
localparam PARSER_PTYPE_RAM_EXTRACT_IDX_RESET = 4'h0;
localparam PARSER_PTYPE_RAM_PTYPE_LO = 0;
localparam PARSER_PTYPE_RAM_PTYPE_HI = 9;
localparam PARSER_PTYPE_RAM_PTYPE_RESET = 10'h0;
localparam PARSER_PTYPE_RAM_USEMASK = 64'h3FFF;
localparam PARSER_PTYPE_RAM_RO_MASK = 64'h0;
localparam PARSER_PTYPE_RAM_WO_MASK = 64'h0;
localparam PARSER_PTYPE_RAM_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic  [7:0] OFFSET;  // RW
    logic  [7:0] PROTOCOL_ID;  // RW
} PARSER_EXTRACT_CFG_t;

localparam PARSER_EXTRACT_CFG_REG_STRIDE = 48'h8;
localparam PARSER_EXTRACT_CFG_REG_ENTRIES = 80;
localparam PARSER_EXTRACT_CFG_REGFILE_STRIDE = 48'h400;
localparam PARSER_EXTRACT_CFG_REGFILE_ENTRIES = 16;
localparam PARSER_EXTRACT_CFG_CR_ADDR = 48'hC000;
localparam PARSER_EXTRACT_CFG_SIZE = 64;
localparam PARSER_EXTRACT_CFG_OFFSET_LO = 8;
localparam PARSER_EXTRACT_CFG_OFFSET_HI = 15;
localparam PARSER_EXTRACT_CFG_OFFSET_RESET = 8'h0;
localparam PARSER_EXTRACT_CFG_PROTOCOL_ID_LO = 0;
localparam PARSER_EXTRACT_CFG_PROTOCOL_ID_HI = 7;
localparam PARSER_EXTRACT_CFG_PROTOCOL_ID_RESET = 8'hff;
localparam PARSER_EXTRACT_CFG_USEMASK = 64'hFFFF;
localparam PARSER_EXTRACT_CFG_RO_MASK = 64'h0;
localparam PARSER_EXTRACT_CFG_WO_MASK = 64'h0;
localparam PARSER_EXTRACT_CFG_RESET = 64'hFF;

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic  [7:0] EXT_DUP_PROTID;  // RW/1C/V
    logic  [7:0] EXT_UNKNOWN_PROTID;  // RW/1C/V
    logic  [7:0] EXT_SEG_BOUNDARY;  // RW/1C/V
} PARSER_COUNTERS_t;

localparam PARSER_COUNTERS_REG_STRIDE = 48'h8;
localparam PARSER_COUNTERS_REG_ENTRIES = 1;
localparam PARSER_COUNTERS_CR_ADDR = 48'h10000;
localparam PARSER_COUNTERS_SIZE = 64;
localparam PARSER_COUNTERS_EXT_DUP_PROTID_LO = 16;
localparam PARSER_COUNTERS_EXT_DUP_PROTID_HI = 23;
localparam PARSER_COUNTERS_EXT_DUP_PROTID_RESET = 8'h0;
localparam PARSER_COUNTERS_EXT_UNKNOWN_PROTID_LO = 8;
localparam PARSER_COUNTERS_EXT_UNKNOWN_PROTID_HI = 15;
localparam PARSER_COUNTERS_EXT_UNKNOWN_PROTID_RESET = 8'h0;
localparam PARSER_COUNTERS_EXT_SEG_BOUNDARY_LO = 0;
localparam PARSER_COUNTERS_EXT_SEG_BOUNDARY_HI = 7;
localparam PARSER_COUNTERS_EXT_SEG_BOUNDARY_RESET = 8'h0;
localparam PARSER_COUNTERS_USEMASK = 64'hFFFFFF;
localparam PARSER_COUNTERS_RO_MASK = 64'h0;
localparam PARSER_COUNTERS_WO_MASK = 64'h0;
localparam PARSER_COUNTERS_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_PARSER_PORT_CFG_t;

typedef logic [7:0] we_PARSER_CSUM_CFG_t;

typedef logic [7:0] we_PARSER_IP_t;

typedef logic [7:0] we_PARSER_IM_t;

typedef logic [7:0] we_PARSER_KEY_W_t;

typedef logic [7:0] we_PARSER_KEY_S_t;

typedef logic [7:0] we_PARSER_ANA_W_t;

typedef logic [7:0] we_PARSER_ANA_S_t;

typedef logic [7:0] we_PARSER_EXC_t;

typedef logic [7:0] we_PARSER_EXT_t;

typedef logic [7:0] we_PARSER_PTYPE_TCAM_t;

typedef logic [7:0] we_PARSER_PTYPE_RAM_t;

typedef logic [7:0] we_PARSER_EXTRACT_CFG_t;

typedef logic [7:0] we_PARSER_COUNTERS_t;

typedef struct packed {
    we_PARSER_PORT_CFG_t PARSER_PORT_CFG;
    we_PARSER_CSUM_CFG_t PARSER_CSUM_CFG;
    we_PARSER_IP_t PARSER_IP;
    we_PARSER_IM_t PARSER_IM;
    we_PARSER_KEY_W_t PARSER_KEY_W;
    we_PARSER_KEY_S_t PARSER_KEY_S;
    we_PARSER_ANA_W_t PARSER_ANA_W;
    we_PARSER_ANA_S_t PARSER_ANA_S;
    we_PARSER_EXC_t PARSER_EXC;
    we_PARSER_EXT_t PARSER_EXT;
    we_PARSER_PTYPE_TCAM_t PARSER_PTYPE_TCAM;
    we_PARSER_PTYPE_RAM_t PARSER_PTYPE_RAM;
    we_PARSER_EXTRACT_CFG_t PARSER_EXTRACT_CFG;
    we_PARSER_COUNTERS_t PARSER_COUNTERS;
} mby_ppe_parser_map_handcoded_t;

typedef logic [7:0] re_PARSER_PORT_CFG_t;

typedef logic [7:0] re_PARSER_CSUM_CFG_t;

typedef logic [7:0] re_PARSER_IP_t;

typedef logic [7:0] re_PARSER_IM_t;

typedef logic [7:0] re_PARSER_KEY_W_t;

typedef logic [7:0] re_PARSER_KEY_S_t;

typedef logic [7:0] re_PARSER_ANA_W_t;

typedef logic [7:0] re_PARSER_ANA_S_t;

typedef logic [7:0] re_PARSER_EXC_t;

typedef logic [7:0] re_PARSER_EXT_t;

typedef logic [7:0] re_PARSER_PTYPE_TCAM_t;

typedef logic [7:0] re_PARSER_PTYPE_RAM_t;

typedef logic [7:0] re_PARSER_EXTRACT_CFG_t;

typedef logic [7:0] re_PARSER_COUNTERS_t;

typedef struct packed {
    re_PARSER_PORT_CFG_t PARSER_PORT_CFG;
    re_PARSER_CSUM_CFG_t PARSER_CSUM_CFG;
    re_PARSER_IP_t PARSER_IP;
    re_PARSER_IM_t PARSER_IM;
    re_PARSER_KEY_W_t PARSER_KEY_W;
    re_PARSER_KEY_S_t PARSER_KEY_S;
    re_PARSER_ANA_W_t PARSER_ANA_W;
    re_PARSER_ANA_S_t PARSER_ANA_S;
    re_PARSER_EXC_t PARSER_EXC;
    re_PARSER_EXT_t PARSER_EXT;
    re_PARSER_PTYPE_TCAM_t PARSER_PTYPE_TCAM;
    re_PARSER_PTYPE_RAM_t PARSER_PTYPE_RAM;
    re_PARSER_EXTRACT_CFG_t PARSER_EXTRACT_CFG;
    re_PARSER_COUNTERS_t PARSER_COUNTERS;
} mby_ppe_parser_map_hc_re_t;

typedef logic handcode_rvalid_PARSER_PORT_CFG_t;

typedef logic handcode_rvalid_PARSER_CSUM_CFG_t;

typedef logic handcode_rvalid_PARSER_IP_t;

typedef logic handcode_rvalid_PARSER_IM_t;

typedef logic handcode_rvalid_PARSER_KEY_W_t;

typedef logic handcode_rvalid_PARSER_KEY_S_t;

typedef logic handcode_rvalid_PARSER_ANA_W_t;

typedef logic handcode_rvalid_PARSER_ANA_S_t;

typedef logic handcode_rvalid_PARSER_EXC_t;

typedef logic handcode_rvalid_PARSER_EXT_t;

typedef logic handcode_rvalid_PARSER_PTYPE_TCAM_t;

typedef logic handcode_rvalid_PARSER_PTYPE_RAM_t;

typedef logic handcode_rvalid_PARSER_EXTRACT_CFG_t;

typedef logic handcode_rvalid_PARSER_COUNTERS_t;

typedef struct packed {
    handcode_rvalid_PARSER_PORT_CFG_t PARSER_PORT_CFG;
    handcode_rvalid_PARSER_CSUM_CFG_t PARSER_CSUM_CFG;
    handcode_rvalid_PARSER_IP_t PARSER_IP;
    handcode_rvalid_PARSER_IM_t PARSER_IM;
    handcode_rvalid_PARSER_KEY_W_t PARSER_KEY_W;
    handcode_rvalid_PARSER_KEY_S_t PARSER_KEY_S;
    handcode_rvalid_PARSER_ANA_W_t PARSER_ANA_W;
    handcode_rvalid_PARSER_ANA_S_t PARSER_ANA_S;
    handcode_rvalid_PARSER_EXC_t PARSER_EXC;
    handcode_rvalid_PARSER_EXT_t PARSER_EXT;
    handcode_rvalid_PARSER_PTYPE_TCAM_t PARSER_PTYPE_TCAM;
    handcode_rvalid_PARSER_PTYPE_RAM_t PARSER_PTYPE_RAM;
    handcode_rvalid_PARSER_EXTRACT_CFG_t PARSER_EXTRACT_CFG;
    handcode_rvalid_PARSER_COUNTERS_t PARSER_COUNTERS;
} mby_ppe_parser_map_hc_rvalid_t;

typedef logic handcode_wvalid_PARSER_PORT_CFG_t;

typedef logic handcode_wvalid_PARSER_CSUM_CFG_t;

typedef logic handcode_wvalid_PARSER_IP_t;

typedef logic handcode_wvalid_PARSER_IM_t;

typedef logic handcode_wvalid_PARSER_KEY_W_t;

typedef logic handcode_wvalid_PARSER_KEY_S_t;

typedef logic handcode_wvalid_PARSER_ANA_W_t;

typedef logic handcode_wvalid_PARSER_ANA_S_t;

typedef logic handcode_wvalid_PARSER_EXC_t;

typedef logic handcode_wvalid_PARSER_EXT_t;

typedef logic handcode_wvalid_PARSER_PTYPE_TCAM_t;

typedef logic handcode_wvalid_PARSER_PTYPE_RAM_t;

typedef logic handcode_wvalid_PARSER_EXTRACT_CFG_t;

typedef logic handcode_wvalid_PARSER_COUNTERS_t;

typedef struct packed {
    handcode_wvalid_PARSER_PORT_CFG_t PARSER_PORT_CFG;
    handcode_wvalid_PARSER_CSUM_CFG_t PARSER_CSUM_CFG;
    handcode_wvalid_PARSER_IP_t PARSER_IP;
    handcode_wvalid_PARSER_IM_t PARSER_IM;
    handcode_wvalid_PARSER_KEY_W_t PARSER_KEY_W;
    handcode_wvalid_PARSER_KEY_S_t PARSER_KEY_S;
    handcode_wvalid_PARSER_ANA_W_t PARSER_ANA_W;
    handcode_wvalid_PARSER_ANA_S_t PARSER_ANA_S;
    handcode_wvalid_PARSER_EXC_t PARSER_EXC;
    handcode_wvalid_PARSER_EXT_t PARSER_EXT;
    handcode_wvalid_PARSER_PTYPE_TCAM_t PARSER_PTYPE_TCAM;
    handcode_wvalid_PARSER_PTYPE_RAM_t PARSER_PTYPE_RAM;
    handcode_wvalid_PARSER_EXTRACT_CFG_t PARSER_EXTRACT_CFG;
    handcode_wvalid_PARSER_COUNTERS_t PARSER_COUNTERS;
} mby_ppe_parser_map_hc_wvalid_t;

typedef logic handcode_error_PARSER_PORT_CFG_t;

typedef logic handcode_error_PARSER_CSUM_CFG_t;

typedef logic handcode_error_PARSER_IP_t;

typedef logic handcode_error_PARSER_IM_t;

typedef logic handcode_error_PARSER_KEY_W_t;

typedef logic handcode_error_PARSER_KEY_S_t;

typedef logic handcode_error_PARSER_ANA_W_t;

typedef logic handcode_error_PARSER_ANA_S_t;

typedef logic handcode_error_PARSER_EXC_t;

typedef logic handcode_error_PARSER_EXT_t;

typedef logic handcode_error_PARSER_PTYPE_TCAM_t;

typedef logic handcode_error_PARSER_PTYPE_RAM_t;

typedef logic handcode_error_PARSER_EXTRACT_CFG_t;

typedef logic handcode_error_PARSER_COUNTERS_t;

typedef struct packed {
    handcode_error_PARSER_PORT_CFG_t PARSER_PORT_CFG;
    handcode_error_PARSER_CSUM_CFG_t PARSER_CSUM_CFG;
    handcode_error_PARSER_IP_t PARSER_IP;
    handcode_error_PARSER_IM_t PARSER_IM;
    handcode_error_PARSER_KEY_W_t PARSER_KEY_W;
    handcode_error_PARSER_KEY_S_t PARSER_KEY_S;
    handcode_error_PARSER_ANA_W_t PARSER_ANA_W;
    handcode_error_PARSER_ANA_S_t PARSER_ANA_S;
    handcode_error_PARSER_EXC_t PARSER_EXC;
    handcode_error_PARSER_EXT_t PARSER_EXT;
    handcode_error_PARSER_PTYPE_TCAM_t PARSER_PTYPE_TCAM;
    handcode_error_PARSER_PTYPE_RAM_t PARSER_PTYPE_RAM;
    handcode_error_PARSER_EXTRACT_CFG_t PARSER_EXTRACT_CFG;
    handcode_error_PARSER_COUNTERS_t PARSER_COUNTERS;
} mby_ppe_parser_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    PARSER_PORT_CFG_t PARSER_PORT_CFG;
    PARSER_CSUM_CFG_t PARSER_CSUM_CFG;
    PARSER_IP_t PARSER_IP;
    PARSER_IM_t PARSER_IM;
    PARSER_KEY_W_t PARSER_KEY_W;
    PARSER_KEY_S_t PARSER_KEY_S;
    PARSER_ANA_W_t PARSER_ANA_W;
    PARSER_ANA_S_t PARSER_ANA_S;
    PARSER_EXC_t PARSER_EXC;
    PARSER_EXT_t PARSER_EXT;
    PARSER_PTYPE_TCAM_t PARSER_PTYPE_TCAM;
    PARSER_PTYPE_RAM_t PARSER_PTYPE_RAM;
    PARSER_EXTRACT_CFG_t PARSER_EXTRACT_CFG;
    PARSER_COUNTERS_t PARSER_COUNTERS;
} mby_ppe_parser_map_hc_reg_read_t;

typedef struct packed {
    PARSER_PORT_CFG_t PARSER_PORT_CFG;
    PARSER_CSUM_CFG_t PARSER_CSUM_CFG;
    PARSER_IP_t PARSER_IP;
    PARSER_IM_t PARSER_IM;
    PARSER_KEY_W_t PARSER_KEY_W;
    PARSER_KEY_S_t PARSER_KEY_S;
    PARSER_ANA_W_t PARSER_ANA_W;
    PARSER_ANA_S_t PARSER_ANA_S;
    PARSER_EXC_t PARSER_EXC;
    PARSER_EXT_t PARSER_EXT;
    PARSER_PTYPE_TCAM_t PARSER_PTYPE_TCAM;
    PARSER_PTYPE_RAM_t PARSER_PTYPE_RAM;
    PARSER_EXTRACT_CFG_t PARSER_EXTRACT_CFG;
    PARSER_COUNTERS_t PARSER_COUNTERS;
} mby_ppe_parser_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_parser_map_pkg

`endif // MBY_PPE_PARSER_MAP_PKG_VH
