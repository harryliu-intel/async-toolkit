magic
tech scmos
timestamp 969938860
<< ndiffusion >>
rect -33 389 -31 393
rect -33 386 -29 389
rect -16 380 -8 381
rect -33 376 -29 379
rect -16 376 -8 377
<< pdiffusion >>
rect 31 389 33 393
rect 29 386 33 389
rect 8 380 16 381
rect 8 376 16 377
rect 29 376 33 382
<< ntransistor >>
rect -33 379 -29 386
rect -16 377 -8 380
<< ptransistor >>
rect 29 382 33 386
rect 8 377 16 380
<< polysilicon >>
rect -35 380 -33 386
rect -37 379 -33 380
rect -29 379 -25 386
rect -2 380 2 389
rect 25 382 29 386
rect 33 382 35 386
rect -20 377 -16 380
rect -8 377 8 380
rect 16 377 20 380
<< ndcontact >>
rect -31 389 -23 397
rect -16 381 -8 389
rect -33 368 -25 376
rect -16 368 -8 376
<< pdcontact >>
rect 23 389 31 397
rect 8 381 16 389
rect 8 368 16 376
rect 25 368 33 376
<< psubstratepcontact >>
rect -55 380 -47 388
<< nsubstratencontact >>
rect 47 380 55 388
<< polycontact >>
rect -4 389 4 397
rect -43 380 -35 388
rect 35 380 43 388
<< metal1 >>
rect -31 393 -4 397
rect -31 389 -23 393
rect 4 393 31 397
rect -4 389 4 392
rect 23 389 31 393
rect -55 376 -47 388
rect -43 385 -35 388
rect -16 385 -8 389
rect 8 385 16 389
rect 35 385 43 388
rect -43 381 43 385
rect -43 380 -35 381
rect 35 380 43 381
rect 47 376 55 388
rect -55 374 -3 376
rect -55 368 -21 374
rect 3 374 55 376
rect 21 368 55 374
<< m2contact >>
rect -4 392 4 398
rect -21 368 -3 374
rect 3 368 21 374
<< metal2 >>
rect -6 392 6 398
<< m3contact >>
rect -21 368 -3 374
rect 3 368 21 374
<< metal3 >>
rect -21 365 -3 401
rect 3 365 21 401
<< labels >>
rlabel ndcontact -12 372 -12 372 1 GND!
rlabel pdcontact 12 372 12 372 1 Vdd!
rlabel metal1 29 372 29 372 1 Vdd!
rlabel metal1 -29 372 -29 372 1 GND!
rlabel metal2 -6 392 -6 398 3 a
rlabel metal2 6 392 6 398 7 a
rlabel metal1 -51 384 -51 384 3 GND!
rlabel metal1 51 384 51 384 7 Vdd!
<< end >>
