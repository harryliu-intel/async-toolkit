// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

// -----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Subodh Nanal
// Created On   :  09/22/2018
// Description  :  Top Level Fuse Environment
// -----------------------------------------------------------------------------



`ifndef INC_FcFuseEnv
`define INC_FcFuseEnv

`define SLA_PATH_TO_STRING(SIG_PATH) `"SIG_PATH`"

`include "fusegen_param.vh"

class FcFuseEnv extends fuse_pkg::soc_fuses_extend_env;

    `ovm_component_utils_begin(FcFuseEnv)
    `ovm_component_utils_end

    `include "fusegen_api.vh"

    fc_tb_env   tb_env_ptr;
    fc_cfg_obj  fcCfgObj;  

    logic [31:0] idata;
    logic [31:0] soft_strap_base_addr;
    logic [31:0] soft_strap_addr;

    // ------------------------------------------------------------
    // constructor
    // ------------------------------------------------------------
    function new( string n="", ovm_component p = null);
        bit        rc;
        ovm_object temp;

        super.new( n, p);

        //Get a handle to the Flash Memory Space in the BFM.
        //nc = CGEnv::getAVMComponent("spis1");
        //if (!$cast(spis1, nc)) begin
        //    $display("could not get spis1 handle");
        //    $finish(0);
        //end      

        tb_env_ptr = fc_tb_env::get_tb_env();
        fcCfgObj = tb_env_ptr.get_cfg_obj_handle;

    endfunction : new

    // ------------------------------------------------------------
    // build
    // ------------------------------------------------------------
    function void build();
        super.build();
        `ovm_info(get_full_name(), $psprintf("FcFuseEnv: Start of build"), UVM_LOW)
        `ovm_info(get_full_name(), $psprintf("FcFuseEnv: End of build"), UVM_LOW)
    endfunction
    // 

    // ------------------------------------------------------------
    // connect
    // ------------------------------------------------------------
    function void connect();
        super.connect();
        `ovm_info(get_full_name(), $psprintf("FcFuseEnv: Start of connect"), UVM_LOW)
        `ovm_info(get_full_name(), $psprintf("FcFuseEnv: End of connect"), UVM_LOW)
    endfunction : connect

    //-----------------------------------------------------------
    // post_randomize
    //-----------------------------------------------------------
    function void post_randomize();
        //FC::EBGIp_t ip_e;

        super.post_randomize();
    endfunction

    //------------------------------------------------------------
    // Get the number of DW straps generated by fusegen
    //------------------------------------------------------------
    function int get_softstrap_row_count();
        return (1 + SOCFUSEGEN_SOFTSTRAPS_ROWEND - SOCFUSEGEN_SOFTSTRAPS_ROWBEGIN);
    endfunction : get_softstrap_row_count

endclass : FcFuseEnv
`endif //INC_FcFuseEnv

