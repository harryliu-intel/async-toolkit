///
///  INTEL CONFIDENTIAL
///
///  Copyright 2017 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
// ---------------------------------------------------------------------------------------------------------------------
// -- Author : Jim McCormick <jim.mccormick@intel.com>
// -- Project Name : ??? 
// -- Description  : Test execution loop 
// ---------------------------------------------------------------------------------------------------------------------

for (int loop=0; loop<loops; loop++) begin
    $display("---loop%0d start---",loop);

    env.reset();                    // reset the DUT and testbench
    env.load_stimulus(num_reqs);    // put stimulus in a testbench FIFO
    env.drive_stimulus();           // pull stimulus out of testbench FIFO and apply to DUT
    env.wait_done(10);              // wait for 10 clocks after done
    env.final_state_check();        // check for any irregularities in final state of DUT
    env.print_cfg();                // print configuration information
    env.print_stats();              // print statistics
    env.wait_delay(10);             // wait for 10 cycles
    $display("---loop%0d end---",loop);
end
