magic
tech scmos
timestamp 970030488
<< ndiffusion >>
rect -24 516 -8 517
rect -24 508 -8 513
rect -24 500 -8 505
rect -24 496 -8 497
rect -24 487 -8 488
<< pdiffusion >>
rect 8 516 34 517
rect 8 512 34 513
rect 8 503 34 504
rect 8 499 34 500
rect 22 491 34 499
rect 8 490 34 491
rect 8 486 34 487
<< ntransistor >>
rect -24 513 -8 516
rect -24 505 -8 508
rect -24 497 -8 500
<< ptransistor >>
rect 8 513 34 516
rect 8 500 34 503
rect 8 487 34 490
<< polysilicon >>
rect -28 513 -24 516
rect -8 513 8 516
rect 34 513 38 516
rect -28 505 -24 508
rect -8 505 6 508
rect 3 503 6 505
rect 3 500 8 503
rect 34 500 38 503
rect -28 497 -24 500
rect -8 497 -2 500
rect -5 490 -2 497
rect -5 487 8 490
rect 34 487 38 490
<< ndcontact >>
rect -24 517 -8 525
rect -24 488 -8 496
<< pdcontact >>
rect 8 517 34 525
rect 8 504 34 512
rect 8 491 22 499
rect 8 478 34 486
<< psubstratepcontact >>
rect -24 479 -8 487
<< nsubstratencontact >>
rect 43 486 51 494
<< polycontact >>
rect -36 513 -28 521
rect 38 500 46 508
rect -36 492 -28 500
<< metal1 >>
rect -36 519 -28 521
rect -24 517 34 525
rect -36 495 -28 500
rect -4 499 4 517
rect 8 504 34 512
rect -24 483 -8 496
rect -4 491 22 499
rect 26 494 34 504
rect 38 507 46 508
rect 38 500 46 501
rect 26 486 51 494
rect 8 483 34 486
rect -24 479 -21 483
rect 21 478 34 483
<< m2contact >>
rect -4 525 4 531
rect -36 513 -28 519
rect -36 489 -28 495
rect 38 501 46 507
rect -21 477 -3 483
rect 3 477 21 483
<< metal2 >>
rect -6 525 6 531
rect -36 513 0 519
rect 0 501 46 507
rect -36 489 0 495
<< m3contact >>
rect -21 477 -3 483
rect 3 477 21 483
<< metal3 >>
rect -21 474 -3 534
rect 3 474 21 534
<< labels >>
rlabel metal2 0 489 0 495 7 a
rlabel metal2 0 501 0 507 3 b
rlabel metal2 0 513 0 519 7 c
rlabel metal2 0 528 0 528 1 x
rlabel metal1 30 508 30 508 5 Vdd!
rlabel metal1 30 482 30 482 1 Vdd!
rlabel polysilicon 35 501 35 501 1 b
rlabel polysilicon 35 488 35 488 1 a
rlabel metal1 30 521 30 521 5 x
rlabel polysilicon 35 514 35 514 1 c
rlabel metal1 18 495 18 495 1 x
rlabel space 22 477 52 526 3 ^p
rlabel metal1 47 490 47 490 7 Vdd!
rlabel polysilicon -25 514 -25 514 3 c
rlabel polysilicon -25 506 -25 506 3 b
rlabel polysilicon -25 498 -25 498 3 a
rlabel metal1 -12 492 -12 492 1 GND!
rlabel metal1 -12 521 -12 521 1 x
rlabel space -37 478 -23 526 7 ^n
rlabel metal2 -32 516 -32 516 3 c
rlabel metal2 -32 492 -32 492 3 a
rlabel metal2 42 504 42 504 1 b
<< end >>
