// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Raghu P Gudla
// Created On   :  09/22/2018
// Description  :  CHI transaction sequence 
// ----------------------------------------------------------------------------------------------------

class fc_chi_txn_seq extends fc_chi_rn_basic_seq;

    `uvm_object_utils(fc_chi_txn_seq)

    rand svt_chi_rn_transaction::xact_type_enum        chi_xact_type;
   // rand svt_chi_rn_transaction::addr_enum        chi_addr;
rand bit [(`SVT_CHI_MAX_DATA_WIDTH-1):0] chi_data;
rand svt_chi_rn_transaction::data_size_enum        chi_size;
  rand bit [1023:0] data[];
  rand bit [63:0] chi_addr;


   
    // class constructor 
    function new(string name="fc_chi_txn_seq");
        super.new(name);
    endfunction

    virtual task body();
        svt_chi_rn_transaction  chi_tran ;
        svt_configuration get_cfg;
        bit status;
        int txn_id = 0;
        `uvm_info("body", "started running fc_chi_txn_seq..", UVM_LOW)

        super.body();

        // obtain a handle to the port configuration 
        p_sequencer.get_cfg(get_cfg);
        if (!$cast(cfg, get_cfg)) begin
            `uvm_fatal("body", "unable to $cast the configuration to a svt_axi_port_configuration class");
        end

      
      /** set up the write transaction */
      `uvm_create(chi_tran)
      chi_tran.cfg = this.cfg;
      chi_tran.txn_id = txn_id++;
      chi_tran.data_size = svt_chi_rn_transaction::SIZE_64BYTE;
     // chi_tran.addr         = 64'h0001_0000_0100_0010;
      chi_tran.addr      = chi_addr;

        chi_tran.xact_type    = chi_xact_type;

        chi_tran.data = chi_data;

      if(chi_tran.xact_type  == svt_chi_rn_transaction::WRITENOSNPFULL) begin 
        chi_tran.byte_enable = {`SVT_CHI_MAX_BE_WIDTH{1'b1}};
      chi_tran.snp_attr_snp_domain_type = svt_chi_transaction::INNER;
      chi_tran.exp_comp_ack = 1'b0;
      //chi_tran.is_likely_shared = 1'b0;
      //chi_tran.snp_attr_is_snoopable = 1'b0;
      chi_tran.mem_attr_is_early_wr_ack_allowed = 1'b1;
      chi_tran.mem_attr_mem_type = svt_chi_transaction::NORMAL;

      // construct dat_rsvdc to accomodate for the number of tx DAT
      // flits associated to this transaction and then setup the values.
      chi_tran.dat_rsvdc = new[chi_tran.compute_num_dat_flits()];
      foreach (chi_tran.dat_rsvdc[idx])
        chi_tran.dat_rsvdc[idx] = (idx+1);

      // adjust byte_enable field to make sure that the generated byte_enable
      // doesn't violate the protocol.
      chi_tran.post_randomize();
      
      `uvm_info("body", $sformatf("sending CHI WRITE transaction %0s", `SVT_CHI_PRINT_PREFIX(chi_tran)), UVM_LOW);
      end 
       
     else if( chi_xact_type ==  svt_chi_transaction::READNOSNP) begin

      chi_tran.xact_type    = svt_chi_transaction::READNOSNP;
      chi_tran.byte_enable = chi_tran.byte_enable;
      chi_tran.exp_comp_ack = 1'b1;
      chi_tran.is_likely_shared = 1'b0;
      chi_tran.snp_attr_is_snoopable = 1'b0;
      chi_tran.snp_attr_snp_domain_type = svt_chi_transaction::INNER;
      chi_tran.mem_attr_is_early_wr_ack_allowed = 1'b1;
      chi_tran.mem_attr_mem_type = svt_chi_transaction::NORMAL;

     `uvm_info("body", $sformatf("sending CHI READ transaction %0s", `SVT_CHI_PRINT_PREFIX(chi_tran)), UVM_LOW);
    end
   
        `uvm_send(chi_tran)
  
        // wait for the  transaction to complete 
        get_response(rsp);
       
        `uvm_info("body", "exiting...", UVM_LOW)
    endtask: body

endclass: fc_chi_txn_seq



