magic
tech scmos
timestamp 965071348
<< ndiffusion >>
rect -47 25 -39 26
rect -73 11 -61 12
rect -47 21 -39 22
rect -47 12 -39 13
rect -73 3 -61 8
rect -73 -10 -61 0
rect -47 8 -39 9
rect -47 -1 -39 0
rect -73 -18 -61 -13
rect -47 -5 -39 -4
rect -47 -14 -39 -13
rect -47 -18 -39 -17
<< pdiffusion >>
rect -123 25 -113 26
rect -23 25 -15 26
rect -123 21 -113 22
rect -123 12 -113 13
rect -123 8 -113 9
rect -23 21 -15 22
rect -23 12 -15 13
rect -115 0 -113 8
rect -100 5 -96 8
rect -123 -1 -113 0
rect -100 -1 -96 2
rect -123 -5 -113 -4
rect -100 -10 -89 -9
rect -23 8 -15 9
rect -23 -1 -15 0
rect -123 -14 -113 -13
rect -123 -18 -113 -17
rect -100 -18 -89 -13
rect -23 -5 -15 -4
rect -23 -14 -15 -13
rect -23 -18 -15 -17
<< ntransistor >>
rect -47 22 -39 25
rect -73 8 -61 11
rect -47 9 -39 12
rect -73 0 -61 3
rect -47 -4 -39 -1
rect -73 -13 -61 -10
rect -47 -17 -39 -14
<< ptransistor >>
rect -123 22 -113 25
rect -123 9 -113 12
rect -23 22 -15 25
rect -23 9 -15 12
rect -100 2 -96 5
rect -123 -4 -113 -1
rect -23 -4 -15 -1
rect -100 -13 -89 -10
rect -123 -17 -113 -14
rect -23 -17 -15 -14
<< polysilicon >>
rect -128 22 -123 25
rect -113 22 -75 25
rect -52 24 -47 25
rect -128 12 -125 22
rect -128 9 -123 12
rect -113 9 -109 12
rect -128 -1 -125 9
rect -78 11 -75 22
rect -51 22 -47 24
rect -39 22 -23 25
rect -15 22 -11 25
rect -51 16 -49 22
rect -52 12 -49 16
rect -78 8 -73 11
rect -61 8 -57 11
rect -52 9 -47 12
rect -39 9 -23 12
rect -15 9 -11 12
rect -104 2 -100 5
rect -96 3 -84 5
rect -96 2 -83 3
rect -87 0 -83 2
rect -128 -4 -123 -1
rect -113 -4 -109 -1
rect -128 -14 -125 -4
rect -75 0 -73 3
rect -61 0 -57 3
rect -52 -1 -49 9
rect -52 -4 -47 -1
rect -39 -4 -23 -1
rect -15 -4 -11 -1
rect -104 -13 -100 -10
rect -89 -13 -73 -10
rect -61 -13 -57 -10
rect -128 -17 -123 -14
rect -113 -17 -109 -14
rect -52 -14 -49 -4
rect -52 -17 -47 -14
rect -39 -17 -23 -14
rect -15 -17 -11 -14
<< ndcontact >>
rect -47 26 -39 34
rect -73 12 -61 20
rect -47 13 -39 21
rect -47 0 -39 8
rect -47 -13 -39 -5
rect -73 -26 -61 -18
rect -47 -26 -39 -18
<< pdcontact >>
rect -123 26 -113 34
rect -23 26 -15 34
rect -123 13 -113 21
rect -103 8 -95 16
rect -23 13 -15 21
rect -123 0 -115 8
rect -123 -13 -113 -5
rect -100 -9 -89 -1
rect -23 0 -15 8
rect -123 -26 -113 -18
rect -100 -26 -89 -18
rect -23 -13 -15 -5
rect -23 -26 -15 -18
<< polycontact >>
rect -59 16 -51 24
rect -83 -5 -75 3
<< metal1 >>
rect -123 26 -95 34
rect -47 26 -39 34
rect -23 26 -15 34
rect -123 17 -113 21
rect -123 13 -107 17
rect -123 0 -115 8
rect -111 -1 -107 13
rect -103 8 -95 26
rect -59 20 -51 24
rect -73 17 -51 20
rect -91 16 -51 17
rect -91 15 -52 16
rect -91 12 -61 15
rect -47 13 -15 21
rect -91 -1 -87 12
rect -111 -5 -87 -1
rect -83 -1 -75 3
rect -47 0 -39 8
rect -83 -5 -52 -1
rect -35 -5 -27 13
rect -23 0 -15 8
rect -123 -9 -87 -5
rect -56 -9 -15 -5
rect -123 -13 -113 -9
rect -47 -13 -15 -9
rect -123 -26 -89 -18
rect -73 -26 -39 -18
rect -23 -26 -15 -18
<< labels >>
rlabel metal1 -69 16 -69 16 1 _x
rlabel polysilicon -74 1 -74 1 1 x
rlabel polysilicon -74 9 -74 9 1 a
rlabel metal1 -69 -22 -69 -22 1 GND!
rlabel polysilicon -74 -12 -74 -12 1 _PReset!
rlabel polysilicon -124 -15 -124 -15 5 a
rlabel polysilicon -124 -2 -124 -2 5 a
rlabel metal1 -119 -22 -119 -22 1 Vdd!
rlabel polysilicon -124 23 -124 23 1 a
rlabel polysilicon -124 10 -124 10 1 a
rlabel metal1 -119 30 -119 30 5 Vdd!
rlabel metal1 -119 4 -119 4 1 Vdd!
rlabel metal1 -118 -9 -118 -9 5 _x
rlabel metal1 -118 17 -118 17 1 _x
rlabel metal1 -94 -22 -94 -22 1 Vdd!
rlabel polysilicon -88 -12 -88 -12 1 _PReset!
rlabel metal1 -95 -5 -95 -5 1 _x
rlabel polysilicon -101 3 -101 3 1 x
rlabel pdcontact -19 -9 -19 -9 5 x
rlabel pdcontact -19 -22 -19 -22 1 Vdd!
rlabel polysilicon -14 -15 -14 -15 5 _x
rlabel polysilicon -14 -2 -14 -2 5 _x
rlabel polysilicon -48 -15 -48 -15 3 _x
rlabel polysilicon -48 -2 -48 -2 3 _x
rlabel ndcontact -43 -22 -43 -22 1 GND!
rlabel ndcontact -43 -9 -43 -9 5 x
rlabel pdcontact -19 4 -19 4 1 Vdd!
rlabel pdcontact -19 17 -19 17 1 x
rlabel pdcontact -19 30 -19 30 5 Vdd!
rlabel polysilicon -14 23 -14 23 1 _x
rlabel polysilicon -14 10 -14 10 1 _x
rlabel polysilicon -48 23 -48 23 3 _x
rlabel polysilicon -48 10 -48 10 3 _x
rlabel ndcontact -43 30 -43 30 5 GND!
rlabel ndcontact -43 4 -43 4 1 GND!
rlabel ndcontact -43 17 -43 17 1 x
rlabel metal1 -99 12 -99 12 1 Vdd!
rlabel space -15 -26 -10 34 3 ^p2
rlabel space -39 -27 -9 35 3 ^n2
rlabel space -129 -26 -123 34 7 ^p1
<< end >>
