.SUBCKT nch_ulvt_mac s g d b 
.ENDS

.SUBCKT pch_ulvt_mac s g d b 
.ENDS

.SUBCKT ppode_ulvt_mac s g b 
.ENDS

.SUBCKT npode_ulvt_mac s g b 
.ENDS
