magic
tech scmos
timestamp 965070867
<< ndiffusion >>
rect 0 559 8 560
rect 0 551 8 556
rect 0 547 8 548
<< pdiffusion >>
rect 24 564 32 565
rect 24 560 32 561
rect 24 551 32 552
rect 24 547 32 548
<< ntransistor >>
rect 0 556 8 559
rect 0 548 8 551
<< ptransistor >>
rect 24 561 32 564
rect 24 548 32 551
<< polysilicon >>
rect 19 561 24 564
rect 32 561 36 564
rect 19 559 22 561
rect -4 556 0 559
rect 8 556 22 559
rect -4 548 0 551
rect 8 548 24 551
rect 32 548 36 551
<< ndcontact >>
rect 0 560 8 568
rect 0 539 8 547
<< pdcontact >>
rect 24 565 32 573
rect 24 552 32 560
rect 24 539 32 547
<< metal1 >>
rect 0 560 16 568
rect 24 565 32 573
rect 8 552 32 560
rect 0 539 8 547
rect 24 539 32 547
<< labels >>
rlabel metal1 28 556 28 556 1 x
rlabel metal1 28 569 28 569 5 Vdd!
rlabel metal1 28 543 28 543 1 Vdd!
rlabel metal1 4 564 4 564 1 x
rlabel metal1 4 543 4 543 1 GND!
rlabel polysilicon -1 549 -1 549 3 a
rlabel polysilicon -1 557 -1 557 3 b
rlabel polysilicon 33 562 33 562 1 b
rlabel polysilicon 33 549 33 549 1 a
rlabel space -5 539 0 568 7 ^n
rlabel space 32 539 37 573 3 ^p
<< end >>
