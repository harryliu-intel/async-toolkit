// -------------------------------------------------------------------------
// This file binds the formal assertions to the DUT 

   bind mby_top mby_checker mby_checker0 (.*);
