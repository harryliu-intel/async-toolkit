magic
tech scmos
timestamp 962519057
<< ndiffusion >>
rect 116 97 120 100
rect 166 98 170 99
rect 112 96 120 97
rect 112 93 120 94
rect 112 89 116 93
rect 112 88 120 89
rect 166 95 170 96
rect 166 90 170 91
rect 112 85 120 86
rect 116 81 120 85
rect 112 80 120 81
rect 166 87 170 88
rect 166 82 170 83
rect 112 74 120 78
rect 112 71 120 72
rect 166 79 170 80
rect 166 74 170 75
rect 166 71 170 72
<< pdiffusion >>
rect 150 98 154 99
rect 96 94 100 95
rect 96 88 100 92
rect 137 90 140 94
rect 133 88 140 90
rect 150 95 154 96
rect 150 90 154 91
rect 96 85 100 86
rect 96 80 100 81
rect 133 85 140 86
rect 137 82 140 85
rect 150 87 154 88
rect 150 82 154 83
rect 133 80 137 81
rect 96 74 100 78
rect 96 71 100 72
rect 133 71 137 78
rect 150 79 154 80
rect 150 74 154 75
rect 150 71 154 72
<< ntransistor >>
rect 166 96 170 98
rect 112 94 120 96
rect 166 88 170 90
rect 112 86 120 88
rect 166 80 170 82
rect 112 78 120 80
rect 112 72 120 74
rect 166 72 170 74
<< ptransistor >>
rect 150 96 154 98
rect 96 92 100 94
rect 150 88 154 90
rect 96 86 100 88
rect 133 86 140 88
rect 150 80 154 82
rect 96 78 100 80
rect 133 78 137 80
rect 96 72 100 74
rect 150 72 154 74
<< polysilicon >>
rect 146 96 150 98
rect 154 96 166 98
rect 170 96 174 98
rect 108 94 112 96
rect 120 94 123 96
rect 93 92 96 94
rect 100 92 110 94
rect 146 90 148 96
rect 172 90 174 96
rect 146 88 150 90
rect 154 88 166 90
rect 170 88 174 90
rect 93 86 96 88
rect 100 86 112 88
rect 120 86 123 88
rect 130 86 133 88
rect 140 86 143 88
rect 146 82 148 88
rect 172 82 174 88
rect 146 80 150 82
rect 154 80 166 82
rect 170 80 174 82
rect 93 78 96 80
rect 100 78 103 80
rect 109 78 112 80
rect 120 78 133 80
rect 137 78 140 80
rect 93 72 96 74
rect 100 72 103 74
rect 109 72 112 74
rect 120 72 123 74
rect 146 74 148 80
rect 172 74 174 80
rect 146 72 150 74
rect 154 72 166 74
rect 170 72 174 74
<< ndcontact >>
rect 112 97 116 101
rect 166 99 170 103
rect 116 89 120 93
rect 166 91 170 95
rect 112 81 116 85
rect 166 83 170 87
rect 112 67 120 71
rect 166 75 170 79
rect 166 67 170 71
<< pdcontact >>
rect 96 95 100 99
rect 150 99 154 103
rect 133 90 137 94
rect 150 91 154 95
rect 96 81 100 85
rect 133 81 137 85
rect 150 83 154 87
rect 96 67 100 71
rect 150 75 154 79
rect 133 67 137 71
rect 150 67 154 71
<< polycontact >>
rect 142 92 146 96
rect 127 74 131 78
<< metal1 >>
rect 112 100 116 101
rect 96 95 100 99
rect 109 97 116 100
rect 133 99 154 103
rect 166 99 170 103
rect 96 81 100 85
rect 109 85 112 97
rect 116 92 120 93
rect 116 89 123 92
rect 133 90 137 99
rect 142 92 146 96
rect 120 86 123 89
rect 143 86 146 92
rect 150 91 170 95
rect 109 82 116 85
rect 112 81 116 82
rect 133 81 137 85
rect 142 83 146 86
rect 150 83 154 87
rect 158 79 162 91
rect 166 83 170 87
rect 150 78 170 79
rect 127 75 170 78
rect 127 74 131 75
rect 96 67 100 71
rect 112 67 120 71
rect 133 67 154 71
rect 166 67 170 71
<< m2contact >>
rect 100 81 105 86
rect 120 81 125 86
rect 137 81 142 86
<< metal2 >>
rect 100 82 142 86
rect 100 81 105 82
rect 120 81 125 82
rect 137 81 142 82
<< labels >>
rlabel space 169 66 174 104 3 ^n2
rlabel space 153 65 175 105 3 ^p2
rlabel polysilicon 132 87 132 87 1 _PReset!
rlabel polysilicon 95 93 95 93 3 b
rlabel polysilicon 95 87 95 87 3 a
rlabel polysilicon 95 79 95 79 3 b
rlabel polysilicon 95 73 95 73 3 a
rlabel polysilicon 111 73 111 73 1 _PReset!
rlabel space 92 67 96 99 7 ^p1
rlabel pdcontact 152 101 152 101 5 Vdd!
rlabel pdcontact 152 93 152 93 1 x
rlabel pdcontact 152 85 152 85 5 Vdd!
rlabel pdcontact 152 77 152 77 1 x
rlabel pdcontact 152 69 152 69 1 Vdd!
rlabel ndcontact 168 93 168 93 1 x
rlabel ndcontact 168 101 168 101 5 GND!
rlabel ndcontact 168 77 168 77 1 x
rlabel ndcontact 168 85 168 85 5 GND!
rlabel ndcontact 168 69 168 69 1 GND!
rlabel pdcontact 135 92 135 92 1 Vdd!
rlabel pdcontact 98 69 98 69 1 Vdd!
rlabel pdcontact 98 83 98 83 1 _x
rlabel pdcontact 98 97 98 97 5 Vdd!
rlabel ndcontact 116 69 116 69 1 GND!
rlabel pdcontact 135 83 135 83 6 _x
rlabel ndcontact 118 91 118 91 5 _x
rlabel polycontact 129 76 129 76 1 x
rlabel polycontact 144 94 144 94 5 _x
<< end >>
