magic
tech scmos
timestamp 950177980
<< ntransistor >>
rect 63 8 69 10
rect 4 6 8 8
rect 4 0 8 2
rect 48 0 51 8
rect 63 0 69 2
<< ptransistor >>
rect 81 8 85 10
rect 20 6 24 8
rect 33 5 36 8
rect 20 0 24 2
rect 81 0 85 2
<< ndiffusion >>
rect 4 8 8 9
rect 63 11 65 15
rect 63 10 69 11
rect 48 8 51 9
rect 4 2 8 6
rect 4 -1 8 0
rect 63 7 69 8
rect 63 3 65 7
rect 63 2 69 3
rect 48 -1 51 0
rect 63 -1 69 0
<< pdiffusion >>
rect 20 8 24 9
rect 33 8 36 9
rect 81 10 85 11
rect 20 2 24 6
rect 20 -1 24 0
rect 33 -1 36 5
rect 81 7 85 8
rect 81 2 85 3
rect 81 -1 85 0
<< ndcontact >>
rect 4 9 8 13
rect 48 9 52 13
rect 65 11 69 15
rect 4 -5 8 -1
rect 65 3 69 7
rect 48 -5 52 -1
rect 63 -5 69 -1
<< pdcontact >>
rect 20 9 24 13
rect 32 9 36 13
rect 81 11 85 15
rect 81 3 85 7
rect 20 -5 24 -1
rect 81 -5 85 -1
<< nsubstratencontact >>
rect 29 -5 36 -1
<< polysilicon >>
rect 60 8 63 10
rect 69 8 81 10
rect 85 8 88 10
rect 1 6 4 8
rect 8 6 20 8
rect 24 6 27 8
rect 30 5 33 8
rect 36 6 48 8
rect 36 5 39 6
rect 1 0 4 2
rect 8 0 20 2
rect 24 0 27 2
rect 45 0 48 6
rect 51 6 54 8
rect 51 2 52 6
rect 60 2 62 8
rect 86 2 88 8
rect 51 0 54 2
rect 60 0 63 2
rect 69 0 81 2
rect 85 0 88 2
<< polycontact >>
rect 58 10 62 14
rect 52 2 56 6
<< metal1 >>
rect 8 10 20 13
rect 24 10 32 13
rect 36 10 48 13
rect 52 10 58 13
rect 56 3 65 6
rect 69 3 81 7
rect 24 -5 29 -1
<< labels >>
rlabel ndcontact 67 -3 67 -3 1 GND!
rlabel ndcontact 67 13 67 13 5 GND!
rlabel pdcontact 83 5 83 5 1 x
rlabel ndcontact 67 5 67 5 1 x
rlabel pdcontact 83 13 83 13 5 Vdd!
rlabel ndcontact 50 -3 50 -3 1 GND!
rlabel pdcontact 34 11 34 11 4 _x
rlabel nsubstratencontact 34 -3 34 -3 1 Vdd!
rlabel ndcontact 50 11 50 11 5 _x
rlabel pdcontact 22 -3 22 -3 1 Vdd!
rlabel pdcontact 22 11 22 11 1 _x
rlabel pdcontact 83 -3 83 -3 1 Vdd!
rlabel space 84 -6 89 16 3 ^p2
rlabel space 68 -7 90 17 3 ^n2
rlabel ndcontact 6 -3 6 -3 1 GND!
rlabel polysilicon 3 1 3 1 3 a
rlabel polysilicon 3 7 3 7 3 b
rlabel ndcontact 6 11 6 11 1 _x
rlabel space 0 -5 4 13 7 ^n1
rlabel space -1 -6 20 14 7 ^p1
<< end >>
