///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_rx_stats_map_pkg.vh                                
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_RX_STATS_MAP_PKG_VH
`define MBY_PPE_RX_STATS_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_rx_stats_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_rx_stats_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_rx_stats_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_rx_stats_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] FRAME_COUNTER;  // RW/V
} RX_STATS_BANK_FRAME_t;

localparam RX_STATS_BANK_FRAME_REG_STRIDE = 48'h8;
localparam RX_STATS_BANK_FRAME_REG_ENTRIES = 144;
localparam RX_STATS_BANK_FRAME_REGFILE_STRIDE = 48'h1000;
localparam RX_STATS_BANK_FRAME_REGFILE_ENTRIES = 4;
localparam RX_STATS_BANK_FRAME_CR_ADDR = 48'h0;
localparam RX_STATS_BANK_FRAME_SIZE = 64;
localparam RX_STATS_BANK_FRAME_FRAME_COUNTER_LO = 0;
localparam RX_STATS_BANK_FRAME_FRAME_COUNTER_HI = 47;
localparam RX_STATS_BANK_FRAME_FRAME_COUNTER_RESET = 48'h0;
localparam RX_STATS_BANK_FRAME_USEMASK = 64'hFFFFFFFFFFFF;
localparam RX_STATS_BANK_FRAME_RO_MASK = 64'h0;
localparam RX_STATS_BANK_FRAME_WO_MASK = 64'h0;
localparam RX_STATS_BANK_FRAME_RESET = 64'h0;

typedef struct packed {
    logic  [7:0] reserved0;  // RSVD
    logic [55:0] BYTE_COUNTER;  // RW/V
} RX_STATS_BANK_BYTE_t;

localparam RX_STATS_BANK_BYTE_REG_STRIDE = 48'h8;
localparam RX_STATS_BANK_BYTE_REG_ENTRIES = 144;
localparam RX_STATS_BANK_BYTE_REGFILE_STRIDE = 48'h1000;
localparam RX_STATS_BANK_BYTE_REGFILE_ENTRIES = 4;
localparam RX_STATS_BANK_BYTE_CR_ADDR = 48'h4000;
localparam RX_STATS_BANK_BYTE_SIZE = 64;
localparam RX_STATS_BANK_BYTE_BYTE_COUNTER_LO = 0;
localparam RX_STATS_BANK_BYTE_BYTE_COUNTER_HI = 55;
localparam RX_STATS_BANK_BYTE_BYTE_COUNTER_RESET = 56'h0;
localparam RX_STATS_BANK_BYTE_USEMASK = 64'hFFFFFFFFFFFFFF;
localparam RX_STATS_BANK_BYTE_RO_MASK = 64'h0;
localparam RX_STATS_BANK_BYTE_WO_MASK = 64'h0;
localparam RX_STATS_BANK_BYTE_RESET = 64'h0;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic [35:0] FRAME_COUNTER;  // RW/V
} RX_STATS_VLAN_FRAME_t;

localparam RX_STATS_VLAN_FRAME_REG_STRIDE = 48'h8;
localparam RX_STATS_VLAN_FRAME_REG_ENTRIES = 16128;
localparam RX_STATS_VLAN_FRAME_CR_ADDR = 48'h8000;
localparam RX_STATS_VLAN_FRAME_SIZE = 64;
localparam RX_STATS_VLAN_FRAME_FRAME_COUNTER_LO = 0;
localparam RX_STATS_VLAN_FRAME_FRAME_COUNTER_HI = 35;
localparam RX_STATS_VLAN_FRAME_FRAME_COUNTER_RESET = 36'h0;
localparam RX_STATS_VLAN_FRAME_USEMASK = 64'hFFFFFFFFF;
localparam RX_STATS_VLAN_FRAME_RO_MASK = 64'h0;
localparam RX_STATS_VLAN_FRAME_WO_MASK = 64'h0;
localparam RX_STATS_VLAN_FRAME_RESET = 64'h0;

typedef struct packed {
    logic [19:0] reserved0;  // RSVD
    logic [43:0] BYTE_COUNTER;  // RW/V
} RX_STATS_VLAN_BYTE_t;

localparam RX_STATS_VLAN_BYTE_REG_STRIDE = 48'h8;
localparam RX_STATS_VLAN_BYTE_REG_ENTRIES = 16128;
localparam RX_STATS_VLAN_BYTE_CR_ADDR = 48'h28000;
localparam RX_STATS_VLAN_BYTE_SIZE = 64;
localparam RX_STATS_VLAN_BYTE_BYTE_COUNTER_LO = 0;
localparam RX_STATS_VLAN_BYTE_BYTE_COUNTER_HI = 43;
localparam RX_STATS_VLAN_BYTE_BYTE_COUNTER_RESET = 44'h0;
localparam RX_STATS_VLAN_BYTE_USEMASK = 64'hFFFFFFFFFFF;
localparam RX_STATS_VLAN_BYTE_RO_MASK = 64'h0;
localparam RX_STATS_VLAN_BYTE_WO_MASK = 64'h0;
localparam RX_STATS_VLAN_BYTE_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_RX_STATS_BANK_FRAME_t;

typedef logic [7:0] we_RX_STATS_BANK_BYTE_t;

typedef logic [7:0] we_RX_STATS_VLAN_FRAME_t;

typedef logic [7:0] we_RX_STATS_VLAN_BYTE_t;

typedef struct packed {
    we_RX_STATS_BANK_FRAME_t RX_STATS_BANK_FRAME;
    we_RX_STATS_BANK_BYTE_t RX_STATS_BANK_BYTE;
    we_RX_STATS_VLAN_FRAME_t RX_STATS_VLAN_FRAME;
    we_RX_STATS_VLAN_BYTE_t RX_STATS_VLAN_BYTE;
} mby_ppe_rx_stats_map_handcoded_t;

typedef logic [7:0] re_RX_STATS_BANK_FRAME_t;

typedef logic [7:0] re_RX_STATS_BANK_BYTE_t;

typedef logic [7:0] re_RX_STATS_VLAN_FRAME_t;

typedef logic [7:0] re_RX_STATS_VLAN_BYTE_t;

typedef struct packed {
    re_RX_STATS_BANK_FRAME_t RX_STATS_BANK_FRAME;
    re_RX_STATS_BANK_BYTE_t RX_STATS_BANK_BYTE;
    re_RX_STATS_VLAN_FRAME_t RX_STATS_VLAN_FRAME;
    re_RX_STATS_VLAN_BYTE_t RX_STATS_VLAN_BYTE;
} mby_ppe_rx_stats_map_hc_re_t;

typedef logic handcode_rvalid_RX_STATS_BANK_FRAME_t;

typedef logic handcode_rvalid_RX_STATS_BANK_BYTE_t;

typedef logic handcode_rvalid_RX_STATS_VLAN_FRAME_t;

typedef logic handcode_rvalid_RX_STATS_VLAN_BYTE_t;

typedef struct packed {
    handcode_rvalid_RX_STATS_BANK_FRAME_t RX_STATS_BANK_FRAME;
    handcode_rvalid_RX_STATS_BANK_BYTE_t RX_STATS_BANK_BYTE;
    handcode_rvalid_RX_STATS_VLAN_FRAME_t RX_STATS_VLAN_FRAME;
    handcode_rvalid_RX_STATS_VLAN_BYTE_t RX_STATS_VLAN_BYTE;
} mby_ppe_rx_stats_map_hc_rvalid_t;

typedef logic handcode_wvalid_RX_STATS_BANK_FRAME_t;

typedef logic handcode_wvalid_RX_STATS_BANK_BYTE_t;

typedef logic handcode_wvalid_RX_STATS_VLAN_FRAME_t;

typedef logic handcode_wvalid_RX_STATS_VLAN_BYTE_t;

typedef struct packed {
    handcode_wvalid_RX_STATS_BANK_FRAME_t RX_STATS_BANK_FRAME;
    handcode_wvalid_RX_STATS_BANK_BYTE_t RX_STATS_BANK_BYTE;
    handcode_wvalid_RX_STATS_VLAN_FRAME_t RX_STATS_VLAN_FRAME;
    handcode_wvalid_RX_STATS_VLAN_BYTE_t RX_STATS_VLAN_BYTE;
} mby_ppe_rx_stats_map_hc_wvalid_t;

typedef logic handcode_error_RX_STATS_BANK_FRAME_t;

typedef logic handcode_error_RX_STATS_BANK_BYTE_t;

typedef logic handcode_error_RX_STATS_VLAN_FRAME_t;

typedef logic handcode_error_RX_STATS_VLAN_BYTE_t;

typedef struct packed {
    handcode_error_RX_STATS_BANK_FRAME_t RX_STATS_BANK_FRAME;
    handcode_error_RX_STATS_BANK_BYTE_t RX_STATS_BANK_BYTE;
    handcode_error_RX_STATS_VLAN_FRAME_t RX_STATS_VLAN_FRAME;
    handcode_error_RX_STATS_VLAN_BYTE_t RX_STATS_VLAN_BYTE;
} mby_ppe_rx_stats_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    RX_STATS_BANK_FRAME_t RX_STATS_BANK_FRAME;
    RX_STATS_BANK_BYTE_t RX_STATS_BANK_BYTE;
    RX_STATS_VLAN_FRAME_t RX_STATS_VLAN_FRAME;
    RX_STATS_VLAN_BYTE_t RX_STATS_VLAN_BYTE;
} mby_ppe_rx_stats_map_hc_reg_read_t;

typedef struct packed {
    RX_STATS_BANK_FRAME_t RX_STATS_BANK_FRAME;
    RX_STATS_BANK_BYTE_t RX_STATS_BANK_BYTE;
    RX_STATS_VLAN_FRAME_t RX_STATS_VLAN_FRAME;
    RX_STATS_VLAN_BYTE_t RX_STATS_VLAN_BYTE;
} mby_ppe_rx_stats_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_rx_stats_map_pkg

`endif // MBY_PPE_RX_STATS_MAP_PKG_VH
