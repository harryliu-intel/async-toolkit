magic
tech scmos
timestamp 962798678
<< ndiffusion >>
rect -118 49 -110 50
rect -95 57 -87 58
rect -95 49 -87 54
rect -118 45 -110 46
rect -95 45 -87 46
<< pdiffusion >>
rect -18 62 -10 63
rect -18 58 -10 59
rect -65 54 -61 57
rect -65 45 -61 50
rect -48 49 -40 50
rect -18 49 -10 50
rect -48 45 -40 46
rect -18 45 -10 46
<< ntransistor >>
rect -95 54 -87 57
rect -118 46 -110 49
rect -95 46 -87 49
<< ptransistor >>
rect -18 59 -10 62
rect -65 50 -61 54
rect -48 46 -40 49
rect -18 46 -10 49
<< polysilicon >>
rect -108 49 -105 65
rect -85 67 -51 70
rect -85 57 -82 67
rect -54 65 -51 67
rect -99 54 -95 57
rect -87 54 -82 57
rect -54 62 -20 65
rect -23 59 -18 62
rect -10 59 -5 62
rect -122 46 -118 49
rect -110 46 -105 49
rect -99 46 -95 49
rect -87 46 -77 49
rect -69 50 -65 54
rect -61 50 -57 54
rect -8 49 -5 59
rect -52 46 -48 49
rect -40 46 -33 49
rect -22 46 -18 49
rect -10 46 -5 49
<< ndcontact >>
rect -118 50 -110 58
rect -95 58 -87 66
rect -118 37 -110 45
rect -95 37 -87 45
<< pdcontact >>
rect -65 57 -57 65
rect -18 63 -10 71
rect -48 50 -40 58
rect -18 50 -10 58
rect -65 37 -57 45
rect -48 37 -40 45
rect -18 37 -10 45
<< polycontact >>
rect -105 62 -97 70
rect -77 46 -69 54
rect -36 49 -28 57
<< metal1 >>
rect -105 67 -97 70
rect -105 62 -30 67
rect -18 63 -10 71
rect -95 58 -87 62
rect -118 54 -110 58
rect -65 57 -57 62
rect -118 53 -69 54
rect -48 53 -40 58
rect -118 50 -40 53
rect -36 57 -30 62
rect -18 57 -10 58
rect -36 51 -10 57
rect -77 49 -44 50
rect -36 49 -28 51
rect -18 50 -10 51
rect -77 46 -69 49
rect -118 37 -87 45
rect -65 37 -10 45
<< labels >>
rlabel pdcontact -44 41 -44 41 1 Vdd!
rlabel polysilicon -86 55 -86 55 1 a
rlabel metal1 -91 41 -91 41 1 GND!
rlabel metal1 -61 41 -61 41 1 Vdd!
rlabel ndcontact -114 41 -114 41 1 GND!
rlabel polysilicon -9 60 -9 60 1 a
rlabel polysilicon -9 47 -9 47 1 a
rlabel metal1 -14 67 -14 67 5 Vdd!
rlabel metal1 -14 41 -14 41 1 Vdd!
rlabel space -10 37 -4 71 3 ^p
rlabel metal1 -14 54 -14 54 1 x
rlabel metal1 -61 61 -61 61 1 x
rlabel metal1 -91 62 -91 62 1 x
<< end >>
