* CB clock wire test
.temp 25
.param vhi=0.75

.param tcyc=1.0/1.6e9
.param ttran=50p
.param when=tcyc*10

.option resmin=1e-9 accurate delmax=10e-9
.option CSDF probe=0

.include "dut_model.inc"

X1 in out dut_model

* control voltage for load
V1 in 0 PWL (
+     0                                                       0
+    ttran                                                    vhi
+ '  tcyc/2'                                                  vhi
+ 'tcyc/2+ttran'                                              0
+ tcyc                                                        0
+ R
+)

.TRAN step=1e-12 stop='4*when'

.probe tran v(in)
.probe tran v(out)

.end

