///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_trig_apply_misc_map_pkg.vh                         
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_TRIG_APPLY_MISC_MAP_PKG_VH
`define MBY_PPE_TRIG_APPLY_MISC_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_trig_apply_misc_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_trig_apply_misc_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_trig_apply_misc_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_trig_apply_misc_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic [23:0] DROP_MASK;  // RW
} TRIGGER_RATE_LIM_CFG_2_t;

localparam TRIGGER_RATE_LIM_CFG_2_REG_STRIDE = 48'h8;
localparam TRIGGER_RATE_LIM_CFG_2_REG_ENTRIES = 16;
localparam TRIGGER_RATE_LIM_CFG_2_CR_ADDR = 48'h0;
localparam TRIGGER_RATE_LIM_CFG_2_SIZE = 64;
localparam TRIGGER_RATE_LIM_CFG_2_DROP_MASK_LO = 0;
localparam TRIGGER_RATE_LIM_CFG_2_DROP_MASK_HI = 23;
localparam TRIGGER_RATE_LIM_CFG_2_DROP_MASK_RESET = 24'h0;
localparam TRIGGER_RATE_LIM_CFG_2_USEMASK = 64'hFFFFFF;
localparam TRIGGER_RATE_LIM_CFG_2_RO_MASK = 64'h0;
localparam TRIGGER_RATE_LIM_CFG_2_WO_MASK = 64'h0;
localparam TRIGGER_RATE_LIM_CFG_2_RESET = 64'h0;

typedef struct packed {
    logic [63:0] METADATA_MASK;  // RW
} TRIGGER_ACTION_METADATA_MASK_t;

localparam TRIGGER_ACTION_METADATA_MASK_REG_STRIDE = 48'h8;
localparam TRIGGER_ACTION_METADATA_MASK_REG_ENTRIES = 4;
localparam TRIGGER_ACTION_METADATA_MASK_REGFILE_STRIDE = 48'h20;
localparam TRIGGER_ACTION_METADATA_MASK_REGFILE_ENTRIES = 2;
localparam TRIGGER_ACTION_METADATA_MASK_CR_ADDR = 48'h80;
localparam TRIGGER_ACTION_METADATA_MASK_SIZE = 64;
localparam TRIGGER_ACTION_METADATA_MASK_METADATA_MASK_LO = 0;
localparam TRIGGER_ACTION_METADATA_MASK_METADATA_MASK_HI = 63;
localparam TRIGGER_ACTION_METADATA_MASK_METADATA_MASK_RESET = 64'h0;
localparam TRIGGER_ACTION_METADATA_MASK_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_ACTION_METADATA_MASK_RO_MASK = 64'h0;
localparam TRIGGER_ACTION_METADATA_MASK_WO_MASK = 64'h0;
localparam TRIGGER_ACTION_METADATA_MASK_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] PENDING;  // RW/1C/V
} TRIGGER_IP_t;

localparam TRIGGER_IP_REG_STRIDE = 48'h8;
localparam TRIGGER_IP_REG_ENTRIES = 2;
localparam [1:0][47:0] TRIGGER_IP_CR_ADDR = {48'hC8, 48'hC0};
localparam TRIGGER_IP_SIZE = 64;
localparam TRIGGER_IP_PENDING_LO = 0;
localparam TRIGGER_IP_PENDING_HI = 47;
localparam TRIGGER_IP_PENDING_RESET = 48'h0;
localparam TRIGGER_IP_USEMASK = 64'hFFFFFFFFFFFF;
localparam TRIGGER_IP_RO_MASK = 64'h0;
localparam TRIGGER_IP_WO_MASK = 64'h0;
localparam TRIGGER_IP_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] MASK;  // RW
} TRIGGER_IM_t;

localparam TRIGGER_IM_REG_STRIDE = 48'h8;
localparam TRIGGER_IM_REG_ENTRIES = 2;
localparam [1:0][47:0] TRIGGER_IM_CR_ADDR = {48'hD8, 48'hD0};
localparam TRIGGER_IM_SIZE = 64;
localparam TRIGGER_IM_MASK_LO = 0;
localparam TRIGGER_IM_MASK_HI = 47;
localparam TRIGGER_IM_MASK_RESET = 48'hffffffffffff;
localparam TRIGGER_IM_USEMASK = 64'hFFFFFFFFFFFF;
localparam TRIGGER_IM_RO_MASK = 64'h0;
localparam TRIGGER_IM_WO_MASK = 64'h0;
localparam TRIGGER_IM_RESET = 64'hFFFFFFFFFFFF;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] EMPTY;  // RO/V
} TRIGGER_RATE_LIM_EMPTY_t;

localparam TRIGGER_RATE_LIM_EMPTY_REG_STRIDE = 48'h8;
localparam TRIGGER_RATE_LIM_EMPTY_REG_ENTRIES = 1;
localparam [47:0] TRIGGER_RATE_LIM_EMPTY_CR_ADDR = 48'hE0;
localparam TRIGGER_RATE_LIM_EMPTY_SIZE = 64;
localparam TRIGGER_RATE_LIM_EMPTY_EMPTY_LO = 0;
localparam TRIGGER_RATE_LIM_EMPTY_EMPTY_HI = 15;
localparam TRIGGER_RATE_LIM_EMPTY_EMPTY_RESET = 16'hffff;
localparam TRIGGER_RATE_LIM_EMPTY_USEMASK = 64'hFFFF;
localparam TRIGGER_RATE_LIM_EMPTY_RO_MASK = 64'hFFFF;
localparam TRIGGER_RATE_LIM_EMPTY_WO_MASK = 64'h0;
localparam TRIGGER_RATE_LIM_EMPTY_RESET = 64'hFFFF;

typedef struct packed {
    logic [10:0] reserved0;  // RSVD
    logic  [4:0] PORT;  // RO/V
    logic [47:0] MAC_ADDRESS;  // RO/V
} MA_TCN_FIFO_0_t;

localparam MA_TCN_FIFO_0_REG_STRIDE = 48'h8;
localparam MA_TCN_FIFO_0_REG_ENTRIES = 512;
localparam MA_TCN_FIFO_0_CR_ADDR = 48'h100;
localparam MA_TCN_FIFO_0_SIZE = 64;
localparam MA_TCN_FIFO_0_PORT_LO = 48;
localparam MA_TCN_FIFO_0_PORT_HI = 52;
localparam MA_TCN_FIFO_0_PORT_RESET = 5'h0;
localparam MA_TCN_FIFO_0_MAC_ADDRESS_LO = 0;
localparam MA_TCN_FIFO_0_MAC_ADDRESS_HI = 47;
localparam MA_TCN_FIFO_0_MAC_ADDRESS_RESET = 48'h0;
localparam MA_TCN_FIFO_0_USEMASK = 64'h1FFFFFFFFFFFFF;
localparam MA_TCN_FIFO_0_RO_MASK = 64'h1FFFFFFFFFFFFF;
localparam MA_TCN_FIFO_0_WO_MASK = 64'h0;
localparam MA_TCN_FIFO_0_RESET = 64'h0;

typedef struct packed {
    logic [43:0] reserved0;  // RSVD
    logic  [7:0] L2_DOMAIN;  // RO/V
    logic [11:0] VID;  // RO/V
} MA_TCN_FIFO_1_t;

localparam MA_TCN_FIFO_1_REG_STRIDE = 48'h8;
localparam MA_TCN_FIFO_1_REG_ENTRIES = 512;
localparam MA_TCN_FIFO_1_CR_ADDR = 48'h1100;
localparam MA_TCN_FIFO_1_SIZE = 64;
localparam MA_TCN_FIFO_1_L2_DOMAIN_LO = 12;
localparam MA_TCN_FIFO_1_L2_DOMAIN_HI = 19;
localparam MA_TCN_FIFO_1_L2_DOMAIN_RESET = 8'h0;
localparam MA_TCN_FIFO_1_VID_LO = 0;
localparam MA_TCN_FIFO_1_VID_HI = 11;
localparam MA_TCN_FIFO_1_VID_RESET = 12'h0;
localparam MA_TCN_FIFO_1_USEMASK = 64'hFFFFF;
localparam MA_TCN_FIFO_1_RO_MASK = 64'hFFFFF;
localparam MA_TCN_FIFO_1_WO_MASK = 64'h0;
localparam MA_TCN_FIFO_1_RESET = 64'h0;

typedef struct packed {
    logic [62:0] reserved0;  // RSVD
    logic  [0:0] READY;  // RW/V
} MA_TCN_DEQUEUE_t;

localparam MA_TCN_DEQUEUE_REG_STRIDE = 48'h8;
localparam MA_TCN_DEQUEUE_REG_ENTRIES = 1;
localparam MA_TCN_DEQUEUE_CR_ADDR = 48'h2100;
localparam MA_TCN_DEQUEUE_SIZE = 64;
localparam MA_TCN_DEQUEUE_READY_LO = 0;
localparam MA_TCN_DEQUEUE_READY_HI = 0;
localparam MA_TCN_DEQUEUE_READY_RESET = 1'h0;
localparam MA_TCN_DEQUEUE_USEMASK = 64'h1;
localparam MA_TCN_DEQUEUE_RO_MASK = 64'h0;
localparam MA_TCN_DEQUEUE_WO_MASK = 64'h0;
localparam MA_TCN_DEQUEUE_RESET = 64'h0;

typedef struct packed {
    logic  [9:0] reserved0;  // RSVD
    logic  [0:0] VALID;  // RO/V
    logic  [4:0] PORT;  // RO/V
    logic [47:0] MAC_ADDRESS;  // RO/V
} MA_TCN_DATA_0_t;

localparam MA_TCN_DATA_0_REG_STRIDE = 48'h8;
localparam MA_TCN_DATA_0_REG_ENTRIES = 1;
localparam MA_TCN_DATA_0_CR_ADDR = 48'h2108;
localparam MA_TCN_DATA_0_SIZE = 64;
localparam MA_TCN_DATA_0_VALID_LO = 53;
localparam MA_TCN_DATA_0_VALID_HI = 53;
localparam MA_TCN_DATA_0_VALID_RESET = 1'h0;
localparam MA_TCN_DATA_0_PORT_LO = 48;
localparam MA_TCN_DATA_0_PORT_HI = 52;
localparam MA_TCN_DATA_0_PORT_RESET = 5'h0;
localparam MA_TCN_DATA_0_MAC_ADDRESS_LO = 0;
localparam MA_TCN_DATA_0_MAC_ADDRESS_HI = 47;
localparam MA_TCN_DATA_0_MAC_ADDRESS_RESET = 48'h0;
localparam MA_TCN_DATA_0_USEMASK = 64'h3FFFFFFFFFFFFF;
localparam MA_TCN_DATA_0_RO_MASK = 64'h3FFFFFFFFFFFFF;
localparam MA_TCN_DATA_0_WO_MASK = 64'h0;
localparam MA_TCN_DATA_0_RESET = 64'h0;

typedef struct packed {
    logic [43:0] reserved0;  // RSVD
    logic  [7:0] L2_DOMAIN;  // RO/V
    logic [11:0] VID;  // RO/V
} MA_TCN_DATA_1_t;

localparam MA_TCN_DATA_1_REG_STRIDE = 48'h8;
localparam MA_TCN_DATA_1_REG_ENTRIES = 1;
localparam MA_TCN_DATA_1_CR_ADDR = 48'h2110;
localparam MA_TCN_DATA_1_SIZE = 64;
localparam MA_TCN_DATA_1_L2_DOMAIN_LO = 12;
localparam MA_TCN_DATA_1_L2_DOMAIN_HI = 19;
localparam MA_TCN_DATA_1_L2_DOMAIN_RESET = 8'h0;
localparam MA_TCN_DATA_1_VID_LO = 0;
localparam MA_TCN_DATA_1_VID_HI = 11;
localparam MA_TCN_DATA_1_VID_RESET = 12'h0;
localparam MA_TCN_DATA_1_USEMASK = 64'hFFFFF;
localparam MA_TCN_DATA_1_RO_MASK = 64'hFFFFF;
localparam MA_TCN_DATA_1_WO_MASK = 64'h0;
localparam MA_TCN_DATA_1_RESET = 64'h0;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [8:0] HEAD;  // RW/V
} MA_TCN_PTR_HEAD_t;

localparam MA_TCN_PTR_HEAD_REG_STRIDE = 48'h8;
localparam MA_TCN_PTR_HEAD_REG_ENTRIES = 1;
localparam MA_TCN_PTR_HEAD_CR_ADDR = 48'h2118;
localparam MA_TCN_PTR_HEAD_SIZE = 64;
localparam MA_TCN_PTR_HEAD_HEAD_LO = 0;
localparam MA_TCN_PTR_HEAD_HEAD_HI = 8;
localparam MA_TCN_PTR_HEAD_HEAD_RESET = 9'h0;
localparam MA_TCN_PTR_HEAD_USEMASK = 64'h1FF;
localparam MA_TCN_PTR_HEAD_RO_MASK = 64'h0;
localparam MA_TCN_PTR_HEAD_WO_MASK = 64'h0;
localparam MA_TCN_PTR_HEAD_RESET = 64'h0;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [8:0] TAIL;  // RW/V
} MA_TCN_PTR_TAIL_t;

localparam MA_TCN_PTR_TAIL_REG_STRIDE = 48'h8;
localparam MA_TCN_PTR_TAIL_REG_ENTRIES = 1;
localparam MA_TCN_PTR_TAIL_CR_ADDR = 48'h2120;
localparam MA_TCN_PTR_TAIL_SIZE = 64;
localparam MA_TCN_PTR_TAIL_TAIL_LO = 0;
localparam MA_TCN_PTR_TAIL_TAIL_HI = 8;
localparam MA_TCN_PTR_TAIL_TAIL_RESET = 9'h0;
localparam MA_TCN_PTR_TAIL_USEMASK = 64'h1FF;
localparam MA_TCN_PTR_TAIL_RO_MASK = 64'h0;
localparam MA_TCN_PTR_TAIL_WO_MASK = 64'h0;
localparam MA_TCN_PTR_TAIL_RESET = 64'h0;

typedef struct packed {
    logic [61:0] reserved0;  // RSVD
    logic  [0:0] PENDING_EVENTS;  // RW/1C/V
    logic  [0:0] TCN_OVERFLOW;  // RW/1C/V
} MA_TCN_IP_t;

localparam MA_TCN_IP_REG_STRIDE = 48'h8;
localparam MA_TCN_IP_REG_ENTRIES = 1;
localparam [47:0] MA_TCN_IP_CR_ADDR = 48'h2128;
localparam MA_TCN_IP_SIZE = 64;
localparam MA_TCN_IP_PENDING_EVENTS_LO = 1;
localparam MA_TCN_IP_PENDING_EVENTS_HI = 1;
localparam MA_TCN_IP_PENDING_EVENTS_RESET = 1'h0;
localparam MA_TCN_IP_TCN_OVERFLOW_LO = 0;
localparam MA_TCN_IP_TCN_OVERFLOW_HI = 0;
localparam MA_TCN_IP_TCN_OVERFLOW_RESET = 1'h0;
localparam MA_TCN_IP_USEMASK = 64'h3;
localparam MA_TCN_IP_RO_MASK = 64'h0;
localparam MA_TCN_IP_WO_MASK = 64'h0;
localparam MA_TCN_IP_RESET = 64'h0;

typedef struct packed {
    logic [61:0] reserved0;  // RSVD
    logic  [0:0] PENDING_EVENTS;  // RW
    logic  [0:0] TCN_OVERFLOW;  // RW
} MA_TCN_IM_t;

localparam MA_TCN_IM_REG_STRIDE = 48'h8;
localparam MA_TCN_IM_REG_ENTRIES = 1;
localparam [47:0] MA_TCN_IM_CR_ADDR = 48'h2130;
localparam MA_TCN_IM_SIZE = 64;
localparam MA_TCN_IM_PENDING_EVENTS_LO = 1;
localparam MA_TCN_IM_PENDING_EVENTS_HI = 1;
localparam MA_TCN_IM_PENDING_EVENTS_RESET = 1'h1;
localparam MA_TCN_IM_TCN_OVERFLOW_LO = 0;
localparam MA_TCN_IM_TCN_OVERFLOW_HI = 0;
localparam MA_TCN_IM_TCN_OVERFLOW_RESET = 1'h1;
localparam MA_TCN_IM_USEMASK = 64'h3;
localparam MA_TCN_IM_RO_MASK = 64'h0;
localparam MA_TCN_IM_WO_MASK = 64'h0;
localparam MA_TCN_IM_RESET = 64'h3;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [8:0] WM;  // RW
} MA_TCN_WM_t;

localparam MA_TCN_WM_REG_STRIDE = 48'h8;
localparam MA_TCN_WM_REG_ENTRIES = 17;
localparam [16:0][47:0] MA_TCN_WM_CR_ADDR = {48'h21C0, 48'h21B8, 48'h21B0, 48'h21A8, 48'h21A0, 48'h2198, 48'h2190, 48'h2188, 48'h2180, 48'h2178, 48'h2170, 48'h2168, 48'h2160, 48'h2158, 48'h2150, 48'h2148, 48'h2140};
localparam MA_TCN_WM_SIZE = 64;
localparam MA_TCN_WM_WM_LO = 0;
localparam MA_TCN_WM_WM_HI = 8;
localparam MA_TCN_WM_WM_RESET = 9'h1e;
localparam MA_TCN_WM_USEMASK = 64'h1FF;
localparam MA_TCN_WM_RO_MASK = 64'h0;
localparam MA_TCN_WM_WO_MASK = 64'h0;
localparam MA_TCN_WM_RESET = 64'h1E;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [8:0] USAGE;  // RW
} MA_TCN_USAGE_t;

localparam MA_TCN_USAGE_REG_STRIDE = 48'h8;
localparam MA_TCN_USAGE_REG_ENTRIES = 17;
localparam [16:0][47:0] MA_TCN_USAGE_CR_ADDR = {48'h2250, 48'h2248, 48'h2240, 48'h2238, 48'h2230, 48'h2228, 48'h2220, 48'h2218, 48'h2210, 48'h2208, 48'h2200, 48'h21F8, 48'h21F0, 48'h21E8, 48'h21E0, 48'h21D8, 48'h21D0};
localparam MA_TCN_USAGE_SIZE = 64;
localparam MA_TCN_USAGE_USAGE_LO = 0;
localparam MA_TCN_USAGE_USAGE_HI = 8;
localparam MA_TCN_USAGE_USAGE_RESET = 9'h0;
localparam MA_TCN_USAGE_USEMASK = 64'h1FF;
localparam MA_TCN_USAGE_RO_MASK = 64'h0;
localparam MA_TCN_USAGE_WO_MASK = 64'h0;
localparam MA_TCN_USAGE_RESET = 64'h0;

typedef struct packed {
    TRIGGER_IP_t [1:0] TRIGGER_IP;
    TRIGGER_IM_t [1:0] TRIGGER_IM;
    TRIGGER_RATE_LIM_EMPTY_t  TRIGGER_RATE_LIM_EMPTY;
    MA_TCN_IP_t  MA_TCN_IP;
    MA_TCN_IM_t  MA_TCN_IM;
    MA_TCN_WM_t [16:0] MA_TCN_WM;
    MA_TCN_USAGE_t [16:0] MA_TCN_USAGE;
} mby_ppe_trig_apply_misc_map_registers_t;

// ===================================================
// load

typedef struct packed {
    logic  [0:0] PENDING;  // RW/1C/V
} load_TRIGGER_IP_t;

typedef struct packed {
    logic  [0:0] PENDING_EVENTS;  // RW/1C/V
    logic  [0:0] TCN_OVERFLOW;  // RW/1C/V
} load_MA_TCN_IP_t;

typedef struct packed {
    load_TRIGGER_IP_t [1:0] TRIGGER_IP;
    load_MA_TCN_IP_t  MA_TCN_IP;
} mby_ppe_trig_apply_misc_map_load_t;

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

typedef struct packed {
    logic [47:0] PENDING;  // RW/1C/V
} new_TRIGGER_IP_t;

typedef struct packed {
    logic [15:0] EMPTY;  // RO/V
} new_TRIGGER_RATE_LIM_EMPTY_t;

typedef struct packed {
    logic  [0:0] PENDING_EVENTS;  // RW/1C/V
    logic  [0:0] TCN_OVERFLOW;  // RW/1C/V
} new_MA_TCN_IP_t;

typedef struct packed {
    new_TRIGGER_IP_t [1:0] TRIGGER_IP;
    new_TRIGGER_RATE_LIM_EMPTY_t  TRIGGER_RATE_LIM_EMPTY;
    new_MA_TCN_IP_t  MA_TCN_IP;
} mby_ppe_trig_apply_misc_map_new_t;

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_TRIGGER_RATE_LIM_CFG_2_t;

typedef logic [7:0] we_TRIGGER_ACTION_METADATA_MASK_t;

typedef logic [7:0] we_MA_TCN_FIFO_0_t;

typedef logic [7:0] we_MA_TCN_FIFO_1_t;

typedef logic [7:0] we_MA_TCN_DEQUEUE_t;

typedef logic [7:0] we_MA_TCN_DATA_0_t;

typedef logic [7:0] we_MA_TCN_DATA_1_t;

typedef logic [7:0] we_MA_TCN_PTR_HEAD_t;

typedef logic [7:0] we_MA_TCN_PTR_TAIL_t;

typedef struct packed {
    we_TRIGGER_RATE_LIM_CFG_2_t TRIGGER_RATE_LIM_CFG_2;
    we_TRIGGER_ACTION_METADATA_MASK_t TRIGGER_ACTION_METADATA_MASK;
    we_MA_TCN_FIFO_0_t MA_TCN_FIFO_0;
    we_MA_TCN_FIFO_1_t MA_TCN_FIFO_1;
    we_MA_TCN_DEQUEUE_t MA_TCN_DEQUEUE;
    we_MA_TCN_DATA_0_t MA_TCN_DATA_0;
    we_MA_TCN_DATA_1_t MA_TCN_DATA_1;
    we_MA_TCN_PTR_HEAD_t MA_TCN_PTR_HEAD;
    we_MA_TCN_PTR_TAIL_t MA_TCN_PTR_TAIL;
} mby_ppe_trig_apply_misc_map_handcoded_t;

typedef logic [7:0] re_TRIGGER_RATE_LIM_CFG_2_t;

typedef logic [7:0] re_TRIGGER_ACTION_METADATA_MASK_t;

typedef logic [7:0] re_MA_TCN_FIFO_0_t;

typedef logic [7:0] re_MA_TCN_FIFO_1_t;

typedef logic [7:0] re_MA_TCN_DEQUEUE_t;

typedef logic [7:0] re_MA_TCN_DATA_0_t;

typedef logic [7:0] re_MA_TCN_DATA_1_t;

typedef logic [7:0] re_MA_TCN_PTR_HEAD_t;

typedef logic [7:0] re_MA_TCN_PTR_TAIL_t;

typedef struct packed {
    re_TRIGGER_RATE_LIM_CFG_2_t TRIGGER_RATE_LIM_CFG_2;
    re_TRIGGER_ACTION_METADATA_MASK_t TRIGGER_ACTION_METADATA_MASK;
    re_MA_TCN_FIFO_0_t MA_TCN_FIFO_0;
    re_MA_TCN_FIFO_1_t MA_TCN_FIFO_1;
    re_MA_TCN_DEQUEUE_t MA_TCN_DEQUEUE;
    re_MA_TCN_DATA_0_t MA_TCN_DATA_0;
    re_MA_TCN_DATA_1_t MA_TCN_DATA_1;
    re_MA_TCN_PTR_HEAD_t MA_TCN_PTR_HEAD;
    re_MA_TCN_PTR_TAIL_t MA_TCN_PTR_TAIL;
} mby_ppe_trig_apply_misc_map_hc_re_t;

typedef logic handcode_rvalid_TRIGGER_RATE_LIM_CFG_2_t;

typedef logic handcode_rvalid_TRIGGER_ACTION_METADATA_MASK_t;

typedef logic handcode_rvalid_MA_TCN_FIFO_0_t;

typedef logic handcode_rvalid_MA_TCN_FIFO_1_t;

typedef logic handcode_rvalid_MA_TCN_DEQUEUE_t;

typedef logic handcode_rvalid_MA_TCN_DATA_0_t;

typedef logic handcode_rvalid_MA_TCN_DATA_1_t;

typedef logic handcode_rvalid_MA_TCN_PTR_HEAD_t;

typedef logic handcode_rvalid_MA_TCN_PTR_TAIL_t;

typedef struct packed {
    handcode_rvalid_TRIGGER_RATE_LIM_CFG_2_t TRIGGER_RATE_LIM_CFG_2;
    handcode_rvalid_TRIGGER_ACTION_METADATA_MASK_t TRIGGER_ACTION_METADATA_MASK;
    handcode_rvalid_MA_TCN_FIFO_0_t MA_TCN_FIFO_0;
    handcode_rvalid_MA_TCN_FIFO_1_t MA_TCN_FIFO_1;
    handcode_rvalid_MA_TCN_DEQUEUE_t MA_TCN_DEQUEUE;
    handcode_rvalid_MA_TCN_DATA_0_t MA_TCN_DATA_0;
    handcode_rvalid_MA_TCN_DATA_1_t MA_TCN_DATA_1;
    handcode_rvalid_MA_TCN_PTR_HEAD_t MA_TCN_PTR_HEAD;
    handcode_rvalid_MA_TCN_PTR_TAIL_t MA_TCN_PTR_TAIL;
} mby_ppe_trig_apply_misc_map_hc_rvalid_t;

typedef logic handcode_wvalid_TRIGGER_RATE_LIM_CFG_2_t;

typedef logic handcode_wvalid_TRIGGER_ACTION_METADATA_MASK_t;

typedef logic handcode_wvalid_MA_TCN_FIFO_0_t;

typedef logic handcode_wvalid_MA_TCN_FIFO_1_t;

typedef logic handcode_wvalid_MA_TCN_DEQUEUE_t;

typedef logic handcode_wvalid_MA_TCN_DATA_0_t;

typedef logic handcode_wvalid_MA_TCN_DATA_1_t;

typedef logic handcode_wvalid_MA_TCN_PTR_HEAD_t;

typedef logic handcode_wvalid_MA_TCN_PTR_TAIL_t;

typedef struct packed {
    handcode_wvalid_TRIGGER_RATE_LIM_CFG_2_t TRIGGER_RATE_LIM_CFG_2;
    handcode_wvalid_TRIGGER_ACTION_METADATA_MASK_t TRIGGER_ACTION_METADATA_MASK;
    handcode_wvalid_MA_TCN_FIFO_0_t MA_TCN_FIFO_0;
    handcode_wvalid_MA_TCN_FIFO_1_t MA_TCN_FIFO_1;
    handcode_wvalid_MA_TCN_DEQUEUE_t MA_TCN_DEQUEUE;
    handcode_wvalid_MA_TCN_DATA_0_t MA_TCN_DATA_0;
    handcode_wvalid_MA_TCN_DATA_1_t MA_TCN_DATA_1;
    handcode_wvalid_MA_TCN_PTR_HEAD_t MA_TCN_PTR_HEAD;
    handcode_wvalid_MA_TCN_PTR_TAIL_t MA_TCN_PTR_TAIL;
} mby_ppe_trig_apply_misc_map_hc_wvalid_t;

typedef logic handcode_error_TRIGGER_RATE_LIM_CFG_2_t;

typedef logic handcode_error_TRIGGER_ACTION_METADATA_MASK_t;

typedef logic handcode_error_MA_TCN_FIFO_0_t;

typedef logic handcode_error_MA_TCN_FIFO_1_t;

typedef logic handcode_error_MA_TCN_DEQUEUE_t;

typedef logic handcode_error_MA_TCN_DATA_0_t;

typedef logic handcode_error_MA_TCN_DATA_1_t;

typedef logic handcode_error_MA_TCN_PTR_HEAD_t;

typedef logic handcode_error_MA_TCN_PTR_TAIL_t;

typedef struct packed {
    handcode_error_TRIGGER_RATE_LIM_CFG_2_t TRIGGER_RATE_LIM_CFG_2;
    handcode_error_TRIGGER_ACTION_METADATA_MASK_t TRIGGER_ACTION_METADATA_MASK;
    handcode_error_MA_TCN_FIFO_0_t MA_TCN_FIFO_0;
    handcode_error_MA_TCN_FIFO_1_t MA_TCN_FIFO_1;
    handcode_error_MA_TCN_DEQUEUE_t MA_TCN_DEQUEUE;
    handcode_error_MA_TCN_DATA_0_t MA_TCN_DATA_0;
    handcode_error_MA_TCN_DATA_1_t MA_TCN_DATA_1;
    handcode_error_MA_TCN_PTR_HEAD_t MA_TCN_PTR_HEAD;
    handcode_error_MA_TCN_PTR_TAIL_t MA_TCN_PTR_TAIL;
} mby_ppe_trig_apply_misc_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    TRIGGER_RATE_LIM_CFG_2_t TRIGGER_RATE_LIM_CFG_2;
    TRIGGER_ACTION_METADATA_MASK_t TRIGGER_ACTION_METADATA_MASK;
    MA_TCN_FIFO_0_t MA_TCN_FIFO_0;
    MA_TCN_FIFO_1_t MA_TCN_FIFO_1;
    MA_TCN_DEQUEUE_t MA_TCN_DEQUEUE;
    MA_TCN_DATA_0_t MA_TCN_DATA_0;
    MA_TCN_DATA_1_t MA_TCN_DATA_1;
    MA_TCN_PTR_HEAD_t MA_TCN_PTR_HEAD;
    MA_TCN_PTR_TAIL_t MA_TCN_PTR_TAIL;
} mby_ppe_trig_apply_misc_map_hc_reg_read_t;

typedef struct packed {
    TRIGGER_RATE_LIM_CFG_2_t TRIGGER_RATE_LIM_CFG_2;
    TRIGGER_ACTION_METADATA_MASK_t TRIGGER_ACTION_METADATA_MASK;
    MA_TCN_FIFO_0_t MA_TCN_FIFO_0;
    MA_TCN_FIFO_1_t MA_TCN_FIFO_1;
    MA_TCN_DEQUEUE_t MA_TCN_DEQUEUE;
    MA_TCN_DATA_0_t MA_TCN_DATA_0;
    MA_TCN_DATA_1_t MA_TCN_DATA_1;
    MA_TCN_PTR_HEAD_t MA_TCN_PTR_HEAD;
    MA_TCN_PTR_TAIL_t MA_TCN_PTR_TAIL;
} mby_ppe_trig_apply_misc_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_trig_apply_misc_map_pkg

`endif // MBY_PPE_TRIG_APPLY_MISC_MAP_PKG_VH
