///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cgrp_em_map_pkg.vh                                 
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_CGRP_EM_MAP_PKG_VH
`define MBY_PPE_CGRP_EM_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_cgrp_em_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_cgrp_em_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_cgrp_em_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_cgrp_em_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [63:0] DATA;  // RW
} HASH_CAM_t;

localparam HASH_CAM_REG_STRIDE = 48'h8;
localparam HASH_CAM_REG_ENTRIES = 8;
localparam HASH_CAM_REGFILE_STRIDE = 48'h40;
localparam HASH_CAM_REGFILE_ENTRIES = 32;
localparam HASH_CAM_CR_ADDR = 48'h0;
localparam HASH_CAM_SIZE = 64;
localparam HASH_CAM_DATA_LO = 0;
localparam HASH_CAM_DATA_HI = 63;
localparam HASH_CAM_DATA_RESET = 64'h0;
localparam HASH_CAM_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam HASH_CAM_RO_MASK = 64'h0;
localparam HASH_CAM_WO_MASK = 64'h0;
localparam HASH_CAM_RESET = 64'h0;

typedef struct packed {
    logic [63:0] MASK;  // RW
} HASH_CAM_EN_t;

localparam HASH_CAM_EN_REG_STRIDE = 48'h8;
localparam HASH_CAM_EN_REG_ENTRIES = 32;
localparam HASH_CAM_EN_REGFILE_STRIDE = 48'h100;
localparam HASH_CAM_EN_REGFILE_ENTRIES = 2;
localparam HASH_CAM_EN_CR_ADDR = 48'h800;
localparam HASH_CAM_EN_SIZE = 64;
localparam HASH_CAM_EN_MASK_LO = 0;
localparam HASH_CAM_EN_MASK_HI = 63;
localparam HASH_CAM_EN_MASK_RESET = 64'h0;
localparam HASH_CAM_EN_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam HASH_CAM_EN_RO_MASK = 64'h0;
localparam HASH_CAM_EN_WO_MASK = 64'h0;
localparam HASH_CAM_EN_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [31:0] KEY8_MASK;  // RW
} KEY_SEL0_t;

localparam KEY_SEL0_REG_STRIDE = 48'h8;
localparam KEY_SEL0_REG_ENTRIES = 64;
localparam KEY_SEL0_REGFILE_STRIDE = 48'h200;
localparam KEY_SEL0_REGFILE_ENTRIES = 2;
localparam KEY_SEL0_CR_ADDR = 48'hC00;
localparam KEY_SEL0_SIZE = 64;
localparam KEY_SEL0_KEY8_MASK_LO = 0;
localparam KEY_SEL0_KEY8_MASK_HI = 31;
localparam KEY_SEL0_KEY8_MASK_RESET = 32'h0;
localparam KEY_SEL0_USEMASK = 64'hFFFFFFFF;
localparam KEY_SEL0_RO_MASK = 64'h0;
localparam KEY_SEL0_WO_MASK = 64'h0;
localparam KEY_SEL0_RESET = 64'h0;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic  [3:0] KEY_MASK_SEL;  // RW
    logic [15:0] KEY32_MASK;  // RW
    logic [31:0] KEY16_MASK;  // RW
} KEY_SEL1_t;

localparam KEY_SEL1_REG_STRIDE = 48'h8;
localparam KEY_SEL1_REG_ENTRIES = 64;
localparam KEY_SEL1_REGFILE_STRIDE = 48'h200;
localparam KEY_SEL1_REGFILE_ENTRIES = 2;
localparam KEY_SEL1_CR_ADDR = 48'h1000;
localparam KEY_SEL1_SIZE = 64;
localparam KEY_SEL1_KEY_MASK_SEL_LO = 48;
localparam KEY_SEL1_KEY_MASK_SEL_HI = 51;
localparam KEY_SEL1_KEY_MASK_SEL_RESET = 4'h0;
localparam KEY_SEL1_KEY32_MASK_LO = 32;
localparam KEY_SEL1_KEY32_MASK_HI = 47;
localparam KEY_SEL1_KEY32_MASK_RESET = 16'h0;
localparam KEY_SEL1_KEY16_MASK_LO = 0;
localparam KEY_SEL1_KEY16_MASK_HI = 31;
localparam KEY_SEL1_KEY16_MASK_RESET = 32'h0;
localparam KEY_SEL1_USEMASK = 64'hFFFFFFFFFFFFF;
localparam KEY_SEL1_RO_MASK = 64'h0;
localparam KEY_SEL1_WO_MASK = 64'h0;
localparam KEY_SEL1_RESET = 64'h0;

typedef struct packed {
    logic [63:0] MASK;  // RW
} KEY_MASK_t;

localparam KEY_MASK_REG_STRIDE = 48'h8;
localparam KEY_MASK_REG_ENTRIES = 32;
localparam KEY_MASK_REGFILE_STRIDE = 48'h100;
localparam KEY_MASK_REGFILE_ENTRIES = 2;
localparam KEY_MASK_CR_ADDR = 48'h1400;
localparam KEY_MASK_SIZE = 64;
localparam KEY_MASK_MASK_LO = 0;
localparam KEY_MASK_MASK_HI = 63;
localparam KEY_MASK_MASK_RESET = 64'h0;
localparam KEY_MASK_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam KEY_MASK_RO_MASK = 64'h0;
localparam KEY_MASK_WO_MASK = 64'h0;
localparam KEY_MASK_RESET = 64'h0;

typedef struct packed {
    logic [31:0] ACTION1;  // RW
    logic [31:0] ACTION0;  // RW
} HASH_MISS_t;

localparam HASH_MISS_REG_STRIDE = 48'h8;
localparam HASH_MISS_REG_ENTRIES = 64;
localparam HASH_MISS_REGFILE_STRIDE = 48'h200;
localparam HASH_MISS_REGFILE_ENTRIES = 2;
localparam HASH_MISS_CR_ADDR = 48'h1800;
localparam HASH_MISS_SIZE = 64;
localparam HASH_MISS_ACTION1_LO = 32;
localparam HASH_MISS_ACTION1_HI = 63;
localparam HASH_MISS_ACTION1_RESET = 32'h0;
localparam HASH_MISS_ACTION0_LO = 0;
localparam HASH_MISS_ACTION0_HI = 31;
localparam HASH_MISS_ACTION0_RESET = 32'h0;
localparam HASH_MISS_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam HASH_MISS_RO_MASK = 64'h0;
localparam HASH_MISS_WO_MASK = 64'h0;
localparam HASH_MISS_RESET = 64'h0;

typedef struct packed {
    logic [14:0] reserved0;  // RSVD
    logic  [0:0] HASH_HI;  // RW
    logic  [0:0] HASH_LO;  // RW
    logic  [0:0] MODE;  // RW
    logic [12:0] BASE_PTR_0;  // RW
    logic [12:0] BASE_PTR_1;  // RW
    logic  [4:0] HASH_SIZE_0;  // RW
    logic  [4:0] HASH_SIZE_1;  // RW
    logic  [4:0] ENTRY_SIZE_0;  // RW
    logic  [4:0] ENTRY_SIZE_1;  // RW
} HASH_CFG_t;

localparam HASH_CFG_REG_STRIDE = 48'h8;
localparam HASH_CFG_REG_ENTRIES = 64;
localparam HASH_CFG_CR_ADDR = 48'h1C00;
localparam HASH_CFG_SIZE = 64;
localparam HASH_CFG_HASH_HI_LO = 48;
localparam HASH_CFG_HASH_HI_HI = 48;
localparam HASH_CFG_HASH_HI_RESET = 1'h0;
localparam HASH_CFG_HASH_LO_LO = 47;
localparam HASH_CFG_HASH_LO_HI = 47;
localparam HASH_CFG_HASH_LO_RESET = 1'h0;
localparam HASH_CFG_MODE_LO = 46;
localparam HASH_CFG_MODE_HI = 46;
localparam HASH_CFG_MODE_RESET = 1'h0;
localparam HASH_CFG_BASE_PTR_0_LO = 33;
localparam HASH_CFG_BASE_PTR_0_HI = 45;
localparam HASH_CFG_BASE_PTR_0_RESET = 13'h0;
localparam HASH_CFG_BASE_PTR_1_LO = 20;
localparam HASH_CFG_BASE_PTR_1_HI = 32;
localparam HASH_CFG_BASE_PTR_1_RESET = 13'h0;
localparam HASH_CFG_HASH_SIZE_0_LO = 15;
localparam HASH_CFG_HASH_SIZE_0_HI = 19;
localparam HASH_CFG_HASH_SIZE_0_RESET = 5'h0;
localparam HASH_CFG_HASH_SIZE_1_LO = 10;
localparam HASH_CFG_HASH_SIZE_1_HI = 14;
localparam HASH_CFG_HASH_SIZE_1_RESET = 5'h0;
localparam HASH_CFG_ENTRY_SIZE_0_LO = 5;
localparam HASH_CFG_ENTRY_SIZE_0_HI = 9;
localparam HASH_CFG_ENTRY_SIZE_0_RESET = 5'h0;
localparam HASH_CFG_ENTRY_SIZE_1_LO = 0;
localparam HASH_CFG_ENTRY_SIZE_1_HI = 4;
localparam HASH_CFG_ENTRY_SIZE_1_RESET = 5'h0;
localparam HASH_CFG_USEMASK = 64'h1FFFFFFFFFFFF;
localparam HASH_CFG_RO_MASK = 64'h0;
localparam HASH_CFG_WO_MASK = 64'h0;
localparam HASH_CFG_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_HASH_CAM_t;

typedef logic [7:0] we_HASH_CAM_EN_t;

typedef logic [7:0] we_KEY_SEL0_t;

typedef logic [7:0] we_KEY_SEL1_t;

typedef logic [7:0] we_KEY_MASK_t;

typedef logic [7:0] we_HASH_MISS_t;

typedef logic [7:0] we_HASH_CFG_t;

typedef struct packed {
    we_HASH_CAM_t HASH_CAM;
    we_HASH_CAM_EN_t HASH_CAM_EN;
    we_KEY_SEL0_t KEY_SEL0;
    we_KEY_SEL1_t KEY_SEL1;
    we_KEY_MASK_t KEY_MASK;
    we_HASH_MISS_t HASH_MISS;
    we_HASH_CFG_t HASH_CFG;
} mby_ppe_cgrp_em_map_handcoded_t;

typedef logic [7:0] re_HASH_CAM_t;

typedef logic [7:0] re_HASH_CAM_EN_t;

typedef logic [7:0] re_KEY_SEL0_t;

typedef logic [7:0] re_KEY_SEL1_t;

typedef logic [7:0] re_KEY_MASK_t;

typedef logic [7:0] re_HASH_MISS_t;

typedef logic [7:0] re_HASH_CFG_t;

typedef struct packed {
    re_HASH_CAM_t HASH_CAM;
    re_HASH_CAM_EN_t HASH_CAM_EN;
    re_KEY_SEL0_t KEY_SEL0;
    re_KEY_SEL1_t KEY_SEL1;
    re_KEY_MASK_t KEY_MASK;
    re_HASH_MISS_t HASH_MISS;
    re_HASH_CFG_t HASH_CFG;
} mby_ppe_cgrp_em_map_hc_re_t;

typedef logic handcode_rvalid_HASH_CAM_t;

typedef logic handcode_rvalid_HASH_CAM_EN_t;

typedef logic handcode_rvalid_KEY_SEL0_t;

typedef logic handcode_rvalid_KEY_SEL1_t;

typedef logic handcode_rvalid_KEY_MASK_t;

typedef logic handcode_rvalid_HASH_MISS_t;

typedef logic handcode_rvalid_HASH_CFG_t;

typedef struct packed {
    handcode_rvalid_HASH_CAM_t HASH_CAM;
    handcode_rvalid_HASH_CAM_EN_t HASH_CAM_EN;
    handcode_rvalid_KEY_SEL0_t KEY_SEL0;
    handcode_rvalid_KEY_SEL1_t KEY_SEL1;
    handcode_rvalid_KEY_MASK_t KEY_MASK;
    handcode_rvalid_HASH_MISS_t HASH_MISS;
    handcode_rvalid_HASH_CFG_t HASH_CFG;
} mby_ppe_cgrp_em_map_hc_rvalid_t;

typedef logic handcode_wvalid_HASH_CAM_t;

typedef logic handcode_wvalid_HASH_CAM_EN_t;

typedef logic handcode_wvalid_KEY_SEL0_t;

typedef logic handcode_wvalid_KEY_SEL1_t;

typedef logic handcode_wvalid_KEY_MASK_t;

typedef logic handcode_wvalid_HASH_MISS_t;

typedef logic handcode_wvalid_HASH_CFG_t;

typedef struct packed {
    handcode_wvalid_HASH_CAM_t HASH_CAM;
    handcode_wvalid_HASH_CAM_EN_t HASH_CAM_EN;
    handcode_wvalid_KEY_SEL0_t KEY_SEL0;
    handcode_wvalid_KEY_SEL1_t KEY_SEL1;
    handcode_wvalid_KEY_MASK_t KEY_MASK;
    handcode_wvalid_HASH_MISS_t HASH_MISS;
    handcode_wvalid_HASH_CFG_t HASH_CFG;
} mby_ppe_cgrp_em_map_hc_wvalid_t;

typedef logic handcode_error_HASH_CAM_t;

typedef logic handcode_error_HASH_CAM_EN_t;

typedef logic handcode_error_KEY_SEL0_t;

typedef logic handcode_error_KEY_SEL1_t;

typedef logic handcode_error_KEY_MASK_t;

typedef logic handcode_error_HASH_MISS_t;

typedef logic handcode_error_HASH_CFG_t;

typedef struct packed {
    handcode_error_HASH_CAM_t HASH_CAM;
    handcode_error_HASH_CAM_EN_t HASH_CAM_EN;
    handcode_error_KEY_SEL0_t KEY_SEL0;
    handcode_error_KEY_SEL1_t KEY_SEL1;
    handcode_error_KEY_MASK_t KEY_MASK;
    handcode_error_HASH_MISS_t HASH_MISS;
    handcode_error_HASH_CFG_t HASH_CFG;
} mby_ppe_cgrp_em_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    HASH_CAM_t HASH_CAM;
    HASH_CAM_EN_t HASH_CAM_EN;
    KEY_SEL0_t KEY_SEL0;
    KEY_SEL1_t KEY_SEL1;
    KEY_MASK_t KEY_MASK;
    HASH_MISS_t HASH_MISS;
    HASH_CFG_t HASH_CFG;
} mby_ppe_cgrp_em_map_hc_reg_read_t;

typedef struct packed {
    HASH_CAM_t HASH_CAM;
    HASH_CAM_EN_t HASH_CAM_EN;
    KEY_SEL0_t KEY_SEL0;
    KEY_SEL1_t KEY_SEL1;
    KEY_MASK_t KEY_MASK;
    HASH_MISS_t HASH_MISS;
    HASH_CFG_t HASH_CFG;
} mby_ppe_cgrp_em_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_cgrp_em_map_pkg

`endif // MBY_PPE_CGRP_EM_MAP_PKG_VH
