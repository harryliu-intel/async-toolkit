///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_nexthop_map.sv                                     
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_nexthop_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_FF
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_FF

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_RSTD


module rtlgen_mby_ppe_nexthop_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_nexthop_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_PH2_FF
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_NEXTHOP_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_NEXTHOP_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_nexthop_map ( //lintra s-2096
    // Clocks


    // Resets



    // Register Inputs
    handcode_reg_rdata_FLOOD_GLORT_TABLE,
    handcode_reg_rdata_INGRESS_VID_TABLE,
    handcode_reg_rdata_MTU_TABLE,
    handcode_reg_rdata_NH_CONFIG,
    handcode_reg_rdata_NH_GROUPS_0,
    handcode_reg_rdata_NH_GROUPS_1,
    handcode_reg_rdata_NH_GROUP_MIN,
    handcode_reg_rdata_NH_NEIGHBORS_0,
    handcode_reg_rdata_NH_NEIGHBORS_1,
    handcode_reg_rdata_NH_PATH_CTRS,
    handcode_reg_rdata_NH_ROUTES,
    handcode_reg_rdata_NH_STATUS,
    handcode_reg_rdata_NH_USED,
    handcode_reg_rdata_NH_WEIGHTS,

    handcode_rvalid_FLOOD_GLORT_TABLE,
    handcode_rvalid_INGRESS_VID_TABLE,
    handcode_rvalid_MTU_TABLE,
    handcode_rvalid_NH_CONFIG,
    handcode_rvalid_NH_GROUPS_0,
    handcode_rvalid_NH_GROUPS_1,
    handcode_rvalid_NH_GROUP_MIN,
    handcode_rvalid_NH_NEIGHBORS_0,
    handcode_rvalid_NH_NEIGHBORS_1,
    handcode_rvalid_NH_PATH_CTRS,
    handcode_rvalid_NH_ROUTES,
    handcode_rvalid_NH_STATUS,
    handcode_rvalid_NH_USED,
    handcode_rvalid_NH_WEIGHTS,

    handcode_wvalid_FLOOD_GLORT_TABLE,
    handcode_wvalid_INGRESS_VID_TABLE,
    handcode_wvalid_MTU_TABLE,
    handcode_wvalid_NH_CONFIG,
    handcode_wvalid_NH_GROUPS_0,
    handcode_wvalid_NH_GROUPS_1,
    handcode_wvalid_NH_GROUP_MIN,
    handcode_wvalid_NH_NEIGHBORS_0,
    handcode_wvalid_NH_NEIGHBORS_1,
    handcode_wvalid_NH_PATH_CTRS,
    handcode_wvalid_NH_ROUTES,
    handcode_wvalid_NH_STATUS,
    handcode_wvalid_NH_USED,
    handcode_wvalid_NH_WEIGHTS,

    handcode_error_FLOOD_GLORT_TABLE,
    handcode_error_INGRESS_VID_TABLE,
    handcode_error_MTU_TABLE,
    handcode_error_NH_CONFIG,
    handcode_error_NH_GROUPS_0,
    handcode_error_NH_GROUPS_1,
    handcode_error_NH_GROUP_MIN,
    handcode_error_NH_NEIGHBORS_0,
    handcode_error_NH_NEIGHBORS_1,
    handcode_error_NH_PATH_CTRS,
    handcode_error_NH_ROUTES,
    handcode_error_NH_STATUS,
    handcode_error_NH_USED,
    handcode_error_NH_WEIGHTS,


    // Register Outputs

    // Register signals for HandCoded registers
    handcode_reg_wdata_FLOOD_GLORT_TABLE,
    handcode_reg_wdata_INGRESS_VID_TABLE,
    handcode_reg_wdata_MTU_TABLE,
    handcode_reg_wdata_NH_CONFIG,
    handcode_reg_wdata_NH_GROUPS_0,
    handcode_reg_wdata_NH_GROUPS_1,
    handcode_reg_wdata_NH_GROUP_MIN,
    handcode_reg_wdata_NH_NEIGHBORS_0,
    handcode_reg_wdata_NH_NEIGHBORS_1,
    handcode_reg_wdata_NH_PATH_CTRS,
    handcode_reg_wdata_NH_ROUTES,
    handcode_reg_wdata_NH_STATUS,
    handcode_reg_wdata_NH_USED,
    handcode_reg_wdata_NH_WEIGHTS,

    we_FLOOD_GLORT_TABLE,
    we_INGRESS_VID_TABLE,
    we_MTU_TABLE,
    we_NH_CONFIG,
    we_NH_GROUPS_0,
    we_NH_GROUPS_1,
    we_NH_GROUP_MIN,
    we_NH_NEIGHBORS_0,
    we_NH_NEIGHBORS_1,
    we_NH_PATH_CTRS,
    we_NH_ROUTES,
    we_NH_STATUS,
    we_NH_USED,
    we_NH_WEIGHTS,

    re_FLOOD_GLORT_TABLE,
    re_INGRESS_VID_TABLE,
    re_MTU_TABLE,
    re_NH_CONFIG,
    re_NH_GROUPS_0,
    re_NH_GROUPS_1,
    re_NH_GROUP_MIN,
    re_NH_NEIGHBORS_0,
    re_NH_NEIGHBORS_1,
    re_NH_PATH_CTRS,
    re_NH_ROUTES,
    re_NH_STATUS,
    re_NH_USED,
    re_NH_WEIGHTS,




    // Config Access
    req,
    ack
    

);

import mby_ppe_nexthop_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:0] MBY_PPE_NEXTHOP_MAP_OFFSET = {MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] NEXTHOP_SB_BAR = 3'b0;
parameter [7:0] NEXTHOP_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;

    // Clocks


    // Resets



    // Register Inputs
input FLOOD_GLORT_TABLE_t  handcode_reg_rdata_FLOOD_GLORT_TABLE;
input INGRESS_VID_TABLE_t  handcode_reg_rdata_INGRESS_VID_TABLE;
input MTU_TABLE_t  handcode_reg_rdata_MTU_TABLE;
input NH_CONFIG_t  handcode_reg_rdata_NH_CONFIG;
input NH_GROUPS_0_t  handcode_reg_rdata_NH_GROUPS_0;
input NH_GROUPS_1_t  handcode_reg_rdata_NH_GROUPS_1;
input NH_GROUP_MIN_t  handcode_reg_rdata_NH_GROUP_MIN;
input NH_NEIGHBORS_0_t  handcode_reg_rdata_NH_NEIGHBORS_0;
input NH_NEIGHBORS_1_t  handcode_reg_rdata_NH_NEIGHBORS_1;
input NH_PATH_CTRS_t  handcode_reg_rdata_NH_PATH_CTRS;
input NH_ROUTES_t  handcode_reg_rdata_NH_ROUTES;
input NH_STATUS_t  handcode_reg_rdata_NH_STATUS;
input NH_USED_t  handcode_reg_rdata_NH_USED;
input NH_WEIGHTS_t  handcode_reg_rdata_NH_WEIGHTS;

input handcode_rvalid_FLOOD_GLORT_TABLE_t  handcode_rvalid_FLOOD_GLORT_TABLE;
input handcode_rvalid_INGRESS_VID_TABLE_t  handcode_rvalid_INGRESS_VID_TABLE;
input handcode_rvalid_MTU_TABLE_t  handcode_rvalid_MTU_TABLE;
input handcode_rvalid_NH_CONFIG_t  handcode_rvalid_NH_CONFIG;
input handcode_rvalid_NH_GROUPS_0_t  handcode_rvalid_NH_GROUPS_0;
input handcode_rvalid_NH_GROUPS_1_t  handcode_rvalid_NH_GROUPS_1;
input handcode_rvalid_NH_GROUP_MIN_t  handcode_rvalid_NH_GROUP_MIN;
input handcode_rvalid_NH_NEIGHBORS_0_t  handcode_rvalid_NH_NEIGHBORS_0;
input handcode_rvalid_NH_NEIGHBORS_1_t  handcode_rvalid_NH_NEIGHBORS_1;
input handcode_rvalid_NH_PATH_CTRS_t  handcode_rvalid_NH_PATH_CTRS;
input handcode_rvalid_NH_ROUTES_t  handcode_rvalid_NH_ROUTES;
input handcode_rvalid_NH_STATUS_t  handcode_rvalid_NH_STATUS;
input handcode_rvalid_NH_USED_t  handcode_rvalid_NH_USED;
input handcode_rvalid_NH_WEIGHTS_t  handcode_rvalid_NH_WEIGHTS;

input handcode_wvalid_FLOOD_GLORT_TABLE_t  handcode_wvalid_FLOOD_GLORT_TABLE;
input handcode_wvalid_INGRESS_VID_TABLE_t  handcode_wvalid_INGRESS_VID_TABLE;
input handcode_wvalid_MTU_TABLE_t  handcode_wvalid_MTU_TABLE;
input handcode_wvalid_NH_CONFIG_t  handcode_wvalid_NH_CONFIG;
input handcode_wvalid_NH_GROUPS_0_t  handcode_wvalid_NH_GROUPS_0;
input handcode_wvalid_NH_GROUPS_1_t  handcode_wvalid_NH_GROUPS_1;
input handcode_wvalid_NH_GROUP_MIN_t  handcode_wvalid_NH_GROUP_MIN;
input handcode_wvalid_NH_NEIGHBORS_0_t  handcode_wvalid_NH_NEIGHBORS_0;
input handcode_wvalid_NH_NEIGHBORS_1_t  handcode_wvalid_NH_NEIGHBORS_1;
input handcode_wvalid_NH_PATH_CTRS_t  handcode_wvalid_NH_PATH_CTRS;
input handcode_wvalid_NH_ROUTES_t  handcode_wvalid_NH_ROUTES;
input handcode_wvalid_NH_STATUS_t  handcode_wvalid_NH_STATUS;
input handcode_wvalid_NH_USED_t  handcode_wvalid_NH_USED;
input handcode_wvalid_NH_WEIGHTS_t  handcode_wvalid_NH_WEIGHTS;

input handcode_error_FLOOD_GLORT_TABLE_t  handcode_error_FLOOD_GLORT_TABLE;
input handcode_error_INGRESS_VID_TABLE_t  handcode_error_INGRESS_VID_TABLE;
input handcode_error_MTU_TABLE_t  handcode_error_MTU_TABLE;
input handcode_error_NH_CONFIG_t  handcode_error_NH_CONFIG;
input handcode_error_NH_GROUPS_0_t  handcode_error_NH_GROUPS_0;
input handcode_error_NH_GROUPS_1_t  handcode_error_NH_GROUPS_1;
input handcode_error_NH_GROUP_MIN_t  handcode_error_NH_GROUP_MIN;
input handcode_error_NH_NEIGHBORS_0_t  handcode_error_NH_NEIGHBORS_0;
input handcode_error_NH_NEIGHBORS_1_t  handcode_error_NH_NEIGHBORS_1;
input handcode_error_NH_PATH_CTRS_t  handcode_error_NH_PATH_CTRS;
input handcode_error_NH_ROUTES_t  handcode_error_NH_ROUTES;
input handcode_error_NH_STATUS_t  handcode_error_NH_STATUS;
input handcode_error_NH_USED_t  handcode_error_NH_USED;
input handcode_error_NH_WEIGHTS_t  handcode_error_NH_WEIGHTS;


    // Register Outputs

    // Register signals for HandCoded registers
output FLOOD_GLORT_TABLE_t  handcode_reg_wdata_FLOOD_GLORT_TABLE;
output INGRESS_VID_TABLE_t  handcode_reg_wdata_INGRESS_VID_TABLE;
output MTU_TABLE_t  handcode_reg_wdata_MTU_TABLE;
output NH_CONFIG_t  handcode_reg_wdata_NH_CONFIG;
output NH_GROUPS_0_t  handcode_reg_wdata_NH_GROUPS_0;
output NH_GROUPS_1_t  handcode_reg_wdata_NH_GROUPS_1;
output NH_GROUP_MIN_t  handcode_reg_wdata_NH_GROUP_MIN;
output NH_NEIGHBORS_0_t  handcode_reg_wdata_NH_NEIGHBORS_0;
output NH_NEIGHBORS_1_t  handcode_reg_wdata_NH_NEIGHBORS_1;
output NH_PATH_CTRS_t  handcode_reg_wdata_NH_PATH_CTRS;
output NH_ROUTES_t  handcode_reg_wdata_NH_ROUTES;
output NH_STATUS_t  handcode_reg_wdata_NH_STATUS;
output NH_USED_t  handcode_reg_wdata_NH_USED;
output NH_WEIGHTS_t  handcode_reg_wdata_NH_WEIGHTS;

output we_FLOOD_GLORT_TABLE_t  we_FLOOD_GLORT_TABLE;
output we_INGRESS_VID_TABLE_t  we_INGRESS_VID_TABLE;
output we_MTU_TABLE_t  we_MTU_TABLE;
output we_NH_CONFIG_t  we_NH_CONFIG;
output we_NH_GROUPS_0_t  we_NH_GROUPS_0;
output we_NH_GROUPS_1_t  we_NH_GROUPS_1;
output we_NH_GROUP_MIN_t  we_NH_GROUP_MIN;
output we_NH_NEIGHBORS_0_t  we_NH_NEIGHBORS_0;
output we_NH_NEIGHBORS_1_t  we_NH_NEIGHBORS_1;
output we_NH_PATH_CTRS_t  we_NH_PATH_CTRS;
output we_NH_ROUTES_t  we_NH_ROUTES;
output we_NH_STATUS_t  we_NH_STATUS;
output we_NH_USED_t  we_NH_USED;
output we_NH_WEIGHTS_t  we_NH_WEIGHTS;

output re_FLOOD_GLORT_TABLE_t  re_FLOOD_GLORT_TABLE;
output re_INGRESS_VID_TABLE_t  re_INGRESS_VID_TABLE;
output re_MTU_TABLE_t  re_MTU_TABLE;
output re_NH_CONFIG_t  re_NH_CONFIG;
output re_NH_GROUPS_0_t  re_NH_GROUPS_0;
output re_NH_GROUPS_1_t  re_NH_GROUPS_1;
output re_NH_GROUP_MIN_t  re_NH_GROUP_MIN;
output re_NH_NEIGHBORS_0_t  re_NH_NEIGHBORS_0;
output re_NH_NEIGHBORS_1_t  re_NH_NEIGHBORS_1;
output re_NH_PATH_CTRS_t  re_NH_PATH_CTRS;
output re_NH_ROUTES_t  re_NH_ROUTES;
output re_NH_STATUS_t  re_NH_STATUS;
output re_NH_USED_t  re_NH_USED;
output re_NH_WEIGHTS_t  re_NH_WEIGHTS;




    // Config Access
input mby_ppe_nexthop_map_cr_req_t  req;
output mby_ppe_nexthop_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_nexthop_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_NEXTHOP_MAP_MEM;
assign case_req_addr_MBY_PPE_NEXTHOP_MAP_MEM = req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_nexthop;
always_comb begin : sb_fid_cond_nexthop_BLOCK
    unique casez (req_fid) 
		NEXTHOP_SB_FID: sb_fid_cond_nexthop = 1;
		default: sb_fid_cond_nexthop = 0;
    endcase 
end


logic sb_bar_cond_nexthop;
always_comb begin : sb_bar_cond_nexthop_BLOCK
    unique casez (req_bar) 
		NEXTHOP_SB_BAR: sb_bar_cond_nexthop = 1;
		default: sb_bar_cond_nexthop = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// NH_CONFIG using HANDCODED_REG template.
logic addr_decode_NH_CONFIG;
logic write_req_NH_CONFIG;
logic read_req_NH_CONFIG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h0,1'b0}: 
         addr_decode_NH_CONFIG = req.valid;
      default: 
         addr_decode_NH_CONFIG = 1'b0; 
   endcase
end

always_comb write_req_NH_CONFIG = f_IsMEMWr(req_opcode) && addr_decode_NH_CONFIG ;
always_comb read_req_NH_CONFIG  = f_IsMEMRd(req_opcode) && addr_decode_NH_CONFIG ;

always_comb we_NH_CONFIG = {8{write_req_NH_CONFIG}} & be;
always_comb re_NH_CONFIG = {8{read_req_NH_CONFIG}} & be;
always_comb handcode_reg_wdata_NH_CONFIG = write_data;


// ----------------------------------------------------------------------
// NH_STATUS using HANDCODED_REG template.
logic addr_decode_NH_STATUS;
logic write_req_NH_STATUS;
logic read_req_NH_STATUS;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h0,1'b1}: 
         addr_decode_NH_STATUS = req.valid;
      default: 
         addr_decode_NH_STATUS = 1'b0; 
   endcase
end

always_comb write_req_NH_STATUS = f_IsMEMWr(req_opcode) && addr_decode_NH_STATUS ;
always_comb read_req_NH_STATUS  = f_IsMEMRd(req_opcode) && addr_decode_NH_STATUS ;

always_comb we_NH_STATUS = {8{write_req_NH_STATUS}} & be;
always_comb re_NH_STATUS = {8{read_req_NH_STATUS}} & be;
always_comb handcode_reg_wdata_NH_STATUS = write_data;


// ----------------------------------------------------------------------
// NH_NEIGHBORS_0 using HANDCODED_REG template.
logic addr_decode_NH_NEIGHBORS_0;
logic write_req_NH_NEIGHBORS_0;
logic read_req_NH_NEIGHBORS_0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b1?,12'h???,1'b?}: 
         addr_decode_NH_NEIGHBORS_0 = req.valid;
      default: 
         addr_decode_NH_NEIGHBORS_0 = 1'b0; 
   endcase
end

always_comb write_req_NH_NEIGHBORS_0 = f_IsMEMWr(req_opcode) && addr_decode_NH_NEIGHBORS_0 ;
always_comb read_req_NH_NEIGHBORS_0  = f_IsMEMRd(req_opcode) && addr_decode_NH_NEIGHBORS_0 ;

always_comb we_NH_NEIGHBORS_0 = {8{write_req_NH_NEIGHBORS_0}} & be;
always_comb re_NH_NEIGHBORS_0 = {8{read_req_NH_NEIGHBORS_0}} & be;
always_comb handcode_reg_wdata_NH_NEIGHBORS_0 = write_data;


// ----------------------------------------------------------------------
// NH_NEIGHBORS_1 using HANDCODED_REG template.
logic addr_decode_NH_NEIGHBORS_1;
logic write_req_NH_NEIGHBORS_1;
logic read_req_NH_NEIGHBORS_1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b10?,12'h???,1'b?}: 
         addr_decode_NH_NEIGHBORS_1 = req.valid;
      default: 
         addr_decode_NH_NEIGHBORS_1 = 1'b0; 
   endcase
end

always_comb write_req_NH_NEIGHBORS_1 = f_IsMEMWr(req_opcode) && addr_decode_NH_NEIGHBORS_1 ;
always_comb read_req_NH_NEIGHBORS_1  = f_IsMEMRd(req_opcode) && addr_decode_NH_NEIGHBORS_1 ;

always_comb we_NH_NEIGHBORS_1 = {8{write_req_NH_NEIGHBORS_1}} & be;
always_comb re_NH_NEIGHBORS_1 = {8{read_req_NH_NEIGHBORS_1}} & be;
always_comb handcode_reg_wdata_NH_NEIGHBORS_1 = write_data;


// ----------------------------------------------------------------------
// NH_GROUPS_0 using HANDCODED_REG template.
logic addr_decode_NH_GROUPS_0;
logic write_req_NH_GROUPS_0;
logic read_req_NH_GROUPS_0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h6,4'b0???,8'h??,1'b?}: 
         addr_decode_NH_GROUPS_0 = req.valid;
      default: 
         addr_decode_NH_GROUPS_0 = 1'b0; 
   endcase
end

always_comb write_req_NH_GROUPS_0 = f_IsMEMWr(req_opcode) && addr_decode_NH_GROUPS_0 ;
always_comb read_req_NH_GROUPS_0  = f_IsMEMRd(req_opcode) && addr_decode_NH_GROUPS_0 ;

always_comb we_NH_GROUPS_0 = {8{write_req_NH_GROUPS_0}} & be;
always_comb re_NH_GROUPS_0 = {8{read_req_NH_GROUPS_0}} & be;
always_comb handcode_reg_wdata_NH_GROUPS_0 = write_data;


// ----------------------------------------------------------------------
// NH_GROUPS_1 using HANDCODED_REG template.
logic addr_decode_NH_GROUPS_1;
logic write_req_NH_GROUPS_1;
logic read_req_NH_GROUPS_1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h6,4'b1???,8'h??,1'b?}: 
         addr_decode_NH_GROUPS_1 = req.valid;
      default: 
         addr_decode_NH_GROUPS_1 = 1'b0; 
   endcase
end

always_comb write_req_NH_GROUPS_1 = f_IsMEMWr(req_opcode) && addr_decode_NH_GROUPS_1 ;
always_comb read_req_NH_GROUPS_1  = f_IsMEMRd(req_opcode) && addr_decode_NH_GROUPS_1 ;

always_comb we_NH_GROUPS_1 = {8{write_req_NH_GROUPS_1}} & be;
always_comb re_NH_GROUPS_1 = {8{read_req_NH_GROUPS_1}} & be;
always_comb handcode_reg_wdata_NH_GROUPS_1 = write_data;


// ----------------------------------------------------------------------
// NH_ROUTES using HANDCODED_REG template.
logic addr_decode_NH_ROUTES;
logic write_req_NH_ROUTES;
logic read_req_NH_ROUTES;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b100?,12'h???,1'b?}: 
         addr_decode_NH_ROUTES = req.valid;
      default: 
         addr_decode_NH_ROUTES = 1'b0; 
   endcase
end

always_comb write_req_NH_ROUTES = f_IsMEMWr(req_opcode) && addr_decode_NH_ROUTES ;
always_comb read_req_NH_ROUTES  = f_IsMEMRd(req_opcode) && addr_decode_NH_ROUTES ;

always_comb we_NH_ROUTES = {8{write_req_NH_ROUTES}} & be;
always_comb re_NH_ROUTES = {8{read_req_NH_ROUTES}} & be;
always_comb handcode_reg_wdata_NH_ROUTES = write_data;


// ----------------------------------------------------------------------
// NH_WEIGHTS using HANDCODED_REG template.
logic addr_decode_NH_WEIGHTS;
logic write_req_NH_WEIGHTS;
logic read_req_NH_WEIGHTS;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b101?,12'h???,1'b?}: 
         addr_decode_NH_WEIGHTS = req.valid;
      default: 
         addr_decode_NH_WEIGHTS = 1'b0; 
   endcase
end

always_comb write_req_NH_WEIGHTS = f_IsMEMWr(req_opcode) && addr_decode_NH_WEIGHTS ;
always_comb read_req_NH_WEIGHTS  = f_IsMEMRd(req_opcode) && addr_decode_NH_WEIGHTS ;

always_comb we_NH_WEIGHTS = {8{write_req_NH_WEIGHTS}} & be;
always_comb re_NH_WEIGHTS = {8{read_req_NH_WEIGHTS}} & be;
always_comb handcode_reg_wdata_NH_WEIGHTS = write_data;


// ----------------------------------------------------------------------
// INGRESS_VID_TABLE using HANDCODED_REG template.
logic addr_decode_INGRESS_VID_TABLE;
logic write_req_INGRESS_VID_TABLE;
logic read_req_INGRESS_VID_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'hC,4'b0???,8'h??,1'b?}: 
         addr_decode_INGRESS_VID_TABLE = req.valid;
      default: 
         addr_decode_INGRESS_VID_TABLE = 1'b0; 
   endcase
end

always_comb write_req_INGRESS_VID_TABLE = f_IsMEMWr(req_opcode) && addr_decode_INGRESS_VID_TABLE ;
always_comb read_req_INGRESS_VID_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_INGRESS_VID_TABLE ;

always_comb we_INGRESS_VID_TABLE = {8{write_req_INGRESS_VID_TABLE}} & be;
always_comb re_INGRESS_VID_TABLE = {8{read_req_INGRESS_VID_TABLE}} & be;
always_comb handcode_reg_wdata_INGRESS_VID_TABLE = write_data;


// ----------------------------------------------------------------------
// FLOOD_GLORT_TABLE using HANDCODED_REG template.
logic addr_decode_FLOOD_GLORT_TABLE;
logic write_req_FLOOD_GLORT_TABLE;
logic read_req_FLOOD_GLORT_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'hC8,4'b0???,4'h?,1'b?}: 
         addr_decode_FLOOD_GLORT_TABLE = req.valid;
      default: 
         addr_decode_FLOOD_GLORT_TABLE = 1'b0; 
   endcase
end

always_comb write_req_FLOOD_GLORT_TABLE = f_IsMEMWr(req_opcode) && addr_decode_FLOOD_GLORT_TABLE ;
always_comb read_req_FLOOD_GLORT_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_FLOOD_GLORT_TABLE ;

always_comb we_FLOOD_GLORT_TABLE = {8{write_req_FLOOD_GLORT_TABLE}} & be;
always_comb re_FLOOD_GLORT_TABLE = {8{read_req_FLOOD_GLORT_TABLE}} & be;
always_comb handcode_reg_wdata_FLOOD_GLORT_TABLE = write_data;


// ----------------------------------------------------------------------
// NH_USED using HANDCODED_REG template.
logic addr_decode_NH_USED;
logic write_req_NH_USED;
logic read_req_NH_USED;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'hC8,4'b1???,4'h?,1'b?}: 
         addr_decode_NH_USED = req.valid;
      default: 
         addr_decode_NH_USED = 1'b0; 
   endcase
end

always_comb write_req_NH_USED = f_IsMEMWr(req_opcode) && addr_decode_NH_USED ;
always_comb read_req_NH_USED  = f_IsMEMRd(req_opcode) && addr_decode_NH_USED ;

always_comb we_NH_USED = {8{write_req_NH_USED}} & be;
always_comb re_NH_USED = {8{read_req_NH_USED}} & be;
always_comb handcode_reg_wdata_NH_USED = write_data;


// ----------------------------------------------------------------------
// NH_PATH_CTRS using HANDCODED_REG template.
logic addr_decode_NH_PATH_CTRS;
logic write_req_NH_PATH_CTRS;
logic read_req_NH_PATH_CTRS;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b111?,12'h???,1'b?}: 
         addr_decode_NH_PATH_CTRS = req.valid;
      default: 
         addr_decode_NH_PATH_CTRS = 1'b0; 
   endcase
end

always_comb write_req_NH_PATH_CTRS = f_IsMEMWr(req_opcode) && addr_decode_NH_PATH_CTRS ;
always_comb read_req_NH_PATH_CTRS  = f_IsMEMRd(req_opcode) && addr_decode_NH_PATH_CTRS ;

always_comb we_NH_PATH_CTRS = {8{write_req_NH_PATH_CTRS}} & be;
always_comb re_NH_PATH_CTRS = {8{read_req_NH_PATH_CTRS}} & be;
always_comb handcode_reg_wdata_NH_PATH_CTRS = write_data;


// ----------------------------------------------------------------------
// NH_GROUP_MIN using HANDCODED_REG template.
logic addr_decode_NH_GROUP_MIN;
logic write_req_NH_GROUP_MIN;
logic read_req_NH_GROUP_MIN;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h100??,1'b?}: 
         addr_decode_NH_GROUP_MIN = req.valid;
      default: 
         addr_decode_NH_GROUP_MIN = 1'b0; 
   endcase
end

always_comb write_req_NH_GROUP_MIN = f_IsMEMWr(req_opcode) && addr_decode_NH_GROUP_MIN ;
always_comb read_req_NH_GROUP_MIN  = f_IsMEMRd(req_opcode) && addr_decode_NH_GROUP_MIN ;

always_comb we_NH_GROUP_MIN = {8{write_req_NH_GROUP_MIN}} & be;
always_comb re_NH_GROUP_MIN = {8{read_req_NH_GROUP_MIN}} & be;
always_comb handcode_reg_wdata_NH_GROUP_MIN = write_data;


// ----------------------------------------------------------------------
// MTU_TABLE using HANDCODED_REG template.
logic addr_decode_MTU_TABLE;
logic write_req_MTU_TABLE;
logic read_req_MTU_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_NEXTHOP_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h1010,4'b00??,1'b?}: 
         addr_decode_MTU_TABLE = req.valid;
      default: 
         addr_decode_MTU_TABLE = 1'b0; 
   endcase
end

always_comb write_req_MTU_TABLE = f_IsMEMWr(req_opcode) && addr_decode_MTU_TABLE ;
always_comb read_req_MTU_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_MTU_TABLE ;

always_comb we_MTU_TABLE = {8{write_req_MTU_TABLE}} & be;
always_comb re_MTU_TABLE = {8{read_req_MTU_TABLE}} & be;
always_comb handcode_reg_wdata_MTU_TABLE = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_NEXTHOP_MAP_MEM) 
           {44'h0,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_CONFIG;
                    ack.read_miss = handcode_error_NH_CONFIG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h0,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_STATUS;
                    ack.read_miss = handcode_error_NH_STATUS;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b1?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_NEIGHBORS_0;
                    ack.read_miss = handcode_error_NH_NEIGHBORS_0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b10?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_NEIGHBORS_1;
                    ack.read_miss = handcode_error_NH_NEIGHBORS_1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h6,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_GROUPS_0;
                    ack.read_miss = handcode_error_NH_GROUPS_0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h6,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_GROUPS_1;
                    ack.read_miss = handcode_error_NH_GROUPS_1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b100?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_ROUTES;
                    ack.read_miss = handcode_error_NH_ROUTES;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b101?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_WEIGHTS;
                    ack.read_miss = handcode_error_NH_WEIGHTS;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'hC,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_INGRESS_VID_TABLE;
                    ack.read_miss = handcode_error_INGRESS_VID_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'hC8,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_FLOOD_GLORT_TABLE;
                    ack.read_miss = handcode_error_FLOOD_GLORT_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'hC8,4'b1???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_USED;
                    ack.read_miss = handcode_error_NH_USED;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b111?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_PATH_CTRS;
                    ack.read_miss = handcode_error_NH_PATH_CTRS;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h100??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_NH_GROUP_MIN;
                    ack.read_miss = handcode_error_NH_GROUP_MIN;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h1010,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MTU_TABLE;
                    ack.read_miss = handcode_error_MTU_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_NEXTHOP_MAP_MEM) 
           {44'h0,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_CONFIG;
                    ack.write_miss = handcode_error_NH_CONFIG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h0,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_STATUS;
                    ack.write_miss = handcode_error_NH_STATUS;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b1?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_NEIGHBORS_0;
                    ack.write_miss = handcode_error_NH_NEIGHBORS_0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b10?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_NEIGHBORS_1;
                    ack.write_miss = handcode_error_NH_NEIGHBORS_1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h6,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_GROUPS_0;
                    ack.write_miss = handcode_error_NH_GROUPS_0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h6,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_GROUPS_1;
                    ack.write_miss = handcode_error_NH_GROUPS_1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b100?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_ROUTES;
                    ack.write_miss = handcode_error_NH_ROUTES;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b101?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_WEIGHTS;
                    ack.write_miss = handcode_error_NH_WEIGHTS;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'hC,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_INGRESS_VID_TABLE;
                    ack.write_miss = handcode_error_INGRESS_VID_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'hC8,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_FLOOD_GLORT_TABLE;
                    ack.write_miss = handcode_error_FLOOD_GLORT_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'hC8,4'b1???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_USED;
                    ack.write_miss = handcode_error_NH_USED;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b111?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_PATH_CTRS;
                    ack.write_miss = handcode_error_NH_PATH_CTRS;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h100??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_NH_GROUP_MIN;
                    ack.write_miss = handcode_error_NH_GROUP_MIN;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h1010,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MTU_TABLE;
                    ack.write_miss = handcode_error_MTU_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_NEXTHOP_MAP_MEM) 
           {44'h0,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_CONFIG;
                 default: read_data = '0;
              endcase
           end
           {44'h0,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_STATUS;
                 default: read_data = '0;
              endcase
           end
           {32'b1?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_NEIGHBORS_0;
                 default: read_data = '0;
              endcase
           end
           {32'b10?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_NEIGHBORS_1;
                 default: read_data = '0;
              endcase
           end
           {32'h6,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_GROUPS_0;
                 default: read_data = '0;
              endcase
           end
           {32'h6,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_GROUPS_1;
                 default: read_data = '0;
              endcase
           end
           {32'b100?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_ROUTES;
                 default: read_data = '0;
              endcase
           end
           {32'b101?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_WEIGHTS;
                 default: read_data = '0;
              endcase
           end
           {32'hC,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_INGRESS_VID_TABLE;
                 default: read_data = '0;
              endcase
           end
           {36'hC8,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_FLOOD_GLORT_TABLE;
                 default: read_data = '0;
              endcase
           end
           {36'hC8,4'b1???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_USED;
                 default: read_data = '0;
              endcase
           end
           {32'b111?,12'h???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_PATH_CTRS;
                 default: read_data = '0;
              endcase
           end
           {44'h100??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_NH_GROUP_MIN;
                 default: read_data = '0;
              endcase
           end
           {40'h1010,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {NEXTHOP_SB_FID,NEXTHOP_SB_BAR}: read_data = handcode_reg_rdata_MTU_TABLE;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {


// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
