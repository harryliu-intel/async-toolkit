//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors. The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//   Author        : Akshay Kotian
//   Project       : MBY
//   Description   : Placeholder for any systemverilog interface which might 
//                  be required to pass information within the TB. 
//------------------------------------------------------------------------------


module mby_wm_tb_top();

//   import uvm_pkg::*;
//  `include "uvm_macros.svh"
//   import sla_pkg::*;
//  `include "sla_macros.svh"

//    mby_wm_intf wm_intf();
//
//    // Add handler of testbench interface
//    initial begin
//        `uvm_info("tb_top", "Setting virtual interfaces", UVM_LOW)
//        slu_resource_db #(virtual mby_wm_intf)::add({"wm_env", ".wm_intf"}, wm_intf, `__FILE__, `__LINE__);
//    end


endmodule

// vim: noai : tw=80 : ts=3 : sw=3 : expandtab : ft=systemverilog

