magic
tech scmos
timestamp 964081429
<< ndiffusion >>
rect 98 144 106 149
rect 140 151 148 152
rect 90 143 106 144
rect 140 143 148 148
rect 90 135 106 140
rect 140 135 148 140
rect 90 130 106 132
rect 90 122 98 130
rect 140 127 148 132
rect 90 121 106 122
rect 90 117 106 118
rect 98 109 106 117
rect 140 123 148 124
rect 140 114 148 115
rect 90 108 106 109
rect 90 100 106 105
rect 140 106 148 111
rect 140 98 148 103
rect 90 96 106 97
rect 90 88 92 96
rect 140 90 148 95
rect 90 87 106 88
rect 90 83 106 84
rect 98 78 106 83
rect 140 86 148 87
rect 140 75 148 76
rect 140 67 148 72
rect 140 59 148 64
rect 140 51 148 56
rect 140 47 148 48
rect 140 38 148 39
rect 140 30 148 35
rect 140 22 148 27
rect 140 14 148 19
rect 140 10 148 11
<< pdiffusion >>
rect 171 155 187 156
rect 209 155 233 156
rect 171 151 187 152
rect 171 142 187 143
rect 209 151 233 152
rect 217 143 233 151
rect 209 142 233 143
rect 171 138 187 139
rect 171 130 179 138
rect 209 138 233 139
rect 171 129 187 130
rect 209 130 217 138
rect 225 130 233 138
rect 209 129 233 130
rect 171 125 187 126
rect 171 116 187 117
rect 209 125 233 126
rect 217 117 233 125
rect 209 116 233 117
rect 171 112 187 113
rect 171 104 179 112
rect 171 103 187 104
rect 209 112 233 113
rect 209 104 217 112
rect 225 104 233 112
rect 209 103 233 104
rect 171 99 187 100
rect 209 99 233 100
rect 171 90 187 91
rect 209 91 217 99
rect 231 91 233 99
rect 209 90 233 91
rect 171 86 187 87
rect 171 77 187 78
rect 209 86 233 87
rect 209 81 225 86
rect 171 73 187 74
rect 171 64 187 65
rect 171 60 187 61
rect 171 52 179 60
rect 171 51 187 52
rect 171 47 187 48
rect 171 38 187 39
rect 171 34 187 35
rect 171 26 179 34
rect 171 25 187 26
rect 171 21 187 22
rect 171 12 187 13
rect 171 8 187 9
<< ntransistor >>
rect 140 148 148 151
rect 90 140 106 143
rect 140 140 148 143
rect 90 132 106 135
rect 140 132 148 135
rect 140 124 148 127
rect 90 118 106 121
rect 90 105 106 108
rect 140 111 148 114
rect 140 103 148 106
rect 90 97 106 100
rect 140 95 148 98
rect 140 87 148 90
rect 90 84 106 87
rect 140 72 148 75
rect 140 64 148 67
rect 140 56 148 59
rect 140 48 148 51
rect 140 35 148 38
rect 140 27 148 30
rect 140 19 148 22
rect 140 11 148 14
<< ptransistor >>
rect 171 152 187 155
rect 209 152 233 155
rect 171 139 187 142
rect 209 139 233 142
rect 171 126 187 129
rect 209 126 233 129
rect 171 113 187 116
rect 209 113 233 116
rect 171 100 187 103
rect 209 100 233 103
rect 171 87 187 90
rect 209 87 233 90
rect 171 74 187 77
rect 171 61 187 64
rect 171 48 187 51
rect 171 35 187 38
rect 171 22 187 25
rect 171 9 187 12
<< polysilicon >>
rect 117 153 138 156
rect 135 151 138 153
rect 166 152 171 155
rect 187 152 192 155
rect 205 152 209 155
rect 233 152 237 155
rect 135 148 140 151
rect 148 148 152 151
rect 86 140 90 143
rect 106 140 122 143
rect 166 143 169 152
rect 130 140 140 143
rect 148 142 169 143
rect 189 142 192 152
rect 148 140 171 142
rect 166 139 171 140
rect 187 139 209 142
rect 233 139 237 142
rect 86 132 90 135
rect 106 132 140 135
rect 148 132 161 135
rect 158 129 161 132
rect 135 124 140 127
rect 148 124 153 127
rect 158 126 171 129
rect 187 126 191 129
rect 199 126 209 129
rect 233 126 237 129
rect 135 121 138 124
rect 86 118 90 121
rect 106 118 138 121
rect 135 114 138 118
rect 150 119 153 124
rect 150 114 157 119
rect 86 105 90 108
rect 106 105 109 108
rect 135 111 140 114
rect 148 111 157 114
rect 165 113 171 116
rect 187 113 209 116
rect 233 113 237 116
rect 165 111 169 113
rect 130 103 140 106
rect 148 103 152 106
rect 166 103 169 111
rect 88 97 90 100
rect 106 97 110 100
rect 166 100 171 103
rect 187 100 191 103
rect 205 100 209 103
rect 233 100 235 103
rect 136 95 140 98
rect 148 95 161 98
rect 158 90 161 95
rect 135 87 140 90
rect 148 87 152 90
rect 158 87 171 90
rect 187 87 191 90
rect 204 87 209 90
rect 233 87 237 90
rect 86 84 90 87
rect 106 84 110 87
rect 135 75 138 87
rect 204 79 207 87
rect 117 72 140 75
rect 148 72 152 75
rect 165 74 171 77
rect 187 74 191 77
rect 204 76 209 79
rect 157 67 160 69
rect 136 64 140 67
rect 148 64 160 67
rect 166 61 171 64
rect 187 61 191 64
rect 166 59 169 61
rect 136 56 140 59
rect 148 56 169 59
rect 130 48 140 51
rect 148 48 171 51
rect 187 48 191 51
rect 130 43 138 48
rect 135 38 138 43
rect 135 35 140 38
rect 148 35 171 38
rect 187 35 191 38
rect 136 27 140 30
rect 148 27 169 30
rect 166 25 169 27
rect 166 22 171 25
rect 187 22 191 25
rect 136 19 140 22
rect 148 19 160 22
rect 157 17 160 19
rect 117 11 140 14
rect 148 11 152 14
rect 165 9 171 12
rect 187 9 191 12
<< ndcontact >>
rect 90 144 98 152
rect 140 152 148 160
rect 98 122 106 130
rect 90 109 98 117
rect 140 115 148 123
rect 92 88 106 96
rect 90 75 98 83
rect 140 76 148 86
rect 140 39 148 47
rect 140 2 148 10
<< pdcontact >>
rect 171 156 187 164
rect 209 156 233 164
rect 171 143 187 151
rect 209 143 217 151
rect 179 130 187 138
rect 217 130 225 138
rect 171 117 187 125
rect 209 117 217 125
rect 179 104 187 112
rect 217 104 225 112
rect 171 91 187 99
rect 217 91 231 99
rect 171 78 187 86
rect 171 65 187 73
rect 225 78 233 86
rect 179 52 187 60
rect 171 39 187 47
rect 179 26 187 34
rect 171 13 187 21
rect 171 0 187 8
<< polycontact >>
rect 109 148 117 156
rect 122 140 130 148
rect 191 126 199 134
rect 109 105 117 113
rect 157 111 165 119
rect 122 103 130 111
rect 80 92 88 100
rect 191 87 199 95
rect 235 95 243 103
rect 109 70 117 78
rect 157 69 165 77
rect 209 71 217 79
rect 191 61 199 69
rect 122 43 130 51
rect 191 22 199 30
rect 109 11 117 19
rect 157 9 165 17
<< metal1 >>
rect 90 144 98 152
rect 109 148 117 156
rect 140 152 148 160
rect 171 156 187 164
rect 209 156 233 164
rect 90 117 94 144
rect 98 122 106 130
rect 90 109 98 117
rect 110 113 116 148
rect 122 140 130 148
rect 171 143 187 151
rect 209 143 217 151
rect 109 105 117 113
rect 123 111 129 140
rect 171 125 175 143
rect 179 130 187 138
rect 191 126 199 134
rect 140 115 148 123
rect 157 111 165 119
rect 171 117 187 125
rect 80 92 88 95
rect 84 83 88 92
rect 92 88 106 96
rect 84 79 98 83
rect 90 75 98 79
rect 110 78 116 105
rect 122 103 130 111
rect 109 70 117 78
rect 110 19 116 70
rect 123 51 129 103
rect 140 76 148 86
rect 157 77 163 111
rect 171 99 175 117
rect 179 104 187 112
rect 171 91 187 99
rect 192 95 198 126
rect 209 125 213 143
rect 217 130 225 138
rect 209 117 217 125
rect 191 87 199 95
rect 171 78 187 86
rect 157 69 165 77
rect 122 43 130 51
rect 140 39 148 47
rect 109 11 117 19
rect 157 17 163 69
rect 171 65 187 73
rect 192 69 198 87
rect 209 79 213 117
rect 221 112 225 130
rect 217 104 225 112
rect 217 91 231 99
rect 235 86 239 95
rect 225 82 239 86
rect 209 71 217 79
rect 225 78 233 82
rect 171 47 175 65
rect 191 61 199 69
rect 179 52 187 60
rect 171 39 187 47
rect 171 21 175 39
rect 179 26 187 34
rect 192 30 198 61
rect 191 22 199 30
rect 140 2 148 10
rect 157 9 165 17
rect 171 13 187 21
rect 171 0 187 8
<< m2contact >>
rect 80 95 88 103
rect 235 95 243 103
<< metal2 >>
rect 80 102 88 103
rect 235 102 243 103
rect 80 96 243 102
rect 80 95 88 96
rect 235 95 243 96
<< labels >>
rlabel polysilicon 170 10 170 10 1 a
rlabel polysilicon 170 75 170 75 1 a
rlabel metal1 175 82 175 82 1 Vdd!
rlabel metal1 175 4 175 4 1 Vdd!
rlabel polysilicon 170 36 170 36 5 _b1
rlabel polysilicon 170 62 170 62 1 _b0
rlabel polysilicon 170 49 170 49 5 _b1
rlabel metal1 175 160 175 160 5 Vdd!
rlabel polysilicon 170 115 170 115 5 a
rlabel polysilicon 170 102 170 102 5 a
rlabel polysilicon 170 153 170 153 1 _b1
rlabel polysilicon 170 140 170 140 1 _b1
rlabel polysilicon 170 127 170 127 1 _b0
rlabel polysilicon 170 88 170 88 1 _b0
rlabel metal1 144 119 144 119 1 x
rlabel polysilicon 139 149 139 149 1 _SReset!
rlabel polysilicon 139 133 139 133 1 _b0
rlabel polysilicon 139 141 139 141 1 _b1
rlabel polysilicon 139 125 139 125 1 a
rlabel polysilicon 139 88 139 88 1 _SReset!
rlabel polysilicon 139 112 139 112 5 a
rlabel metal1 144 156 144 156 1 GND!
rlabel polysilicon 170 23 170 23 1 _b0
rlabel polysilicon 139 96 139 96 1 _b0
rlabel polysilicon 139 104 139 104 1 _b1
rlabel polysilicon 139 20 139 20 1 a
rlabel polysilicon 139 12 139 12 1 _SReset!
rlabel polysilicon 139 65 139 65 5 a
rlabel polysilicon 139 49 139 49 5 _b1
rlabel polysilicon 139 57 139 57 5 _b0
rlabel polysilicon 139 36 139 36 1 _b1
rlabel polysilicon 139 28 139 28 1 _b0
rlabel polysilicon 139 73 139 73 1 _SReset!
rlabel metal1 144 6 144 6 1 GND!
rlabel metal1 144 43 144 43 1 x
rlabel metal1 144 81 144 81 1 GND!
rlabel ndcontact 102 126 102 126 1 x
rlabel polysilicon 107 106 107 106 1 _SReset!
rlabel polysilicon 107 141 107 141 1 _b1
rlabel polysilicon 107 133 107 133 1 _b0
rlabel polysilicon 107 119 107 119 1 a
rlabel polysilicon 107 86 107 86 5 x
rlabel metal1 96 92 96 92 1 GND!
rlabel metal1 221 95 221 95 5 Vdd!
rlabel polysilicon 234 89 234 89 7 x
rlabel metal1 220 160 220 160 5 Vdd!
rlabel polysilicon 234 154 234 154 5 _PReset!
rlabel metal1 213 147 213 147 1 x
rlabel metal1 213 121 213 121 1 x
rlabel polysilicon 234 114 234 114 1 a
rlabel polysilicon 234 127 234 127 1 _b0
rlabel polysilicon 234 140 234 140 1 _b1
rlabel metal1 183 30 183 30 1 x
rlabel metal1 183 56 183 56 1 x
rlabel metal1 183 108 183 108 5 x
rlabel metal1 183 134 183 134 5 Vdd!
rlabel metal1 213 75 213 75 1 x
rlabel space 180 -1 244 165 3 ^p
rlabel space 79 -2 141 161 7 ^n
<< end >>
