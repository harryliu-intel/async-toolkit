///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Mike Jarvis <michael.a.jarvis.com> 
// -- Project Name : MBY 
// -- Description  : mpp (MegaPort Pair) netlist. 
// ------------------------------------------------------------------- 

module mpp (
//Input List
input                   arst_n,                                   //Asynchronous negedge reset     
input                   cclk,                                     
input                   clk,                                      
input            [7:0]  epl0_igr0_rx_data_valid,                  
input         [0:7][71:0]  epl0_igr0_rx_data_w_ecc,                  
input            [7:0]  epl0_igr0_rx_ecc,                         
input            [2:0]  epl0_igr0_rx_flow_control_tc,             
input           [23:0]  epl0_igr0_rx_metadata,                    
input                   epl0_igr0_rx_pfc_xoff,                    
input            [1:0]  epl0_igr0_rx_port_num,                    
input           [35:0]  epl0_igr0_rx_time_stamp,                  
input            [7:0]  epl0_igr1_rx_data_valid,                  
input         [0:7][71:0]  epl0_igr1_rx_data_w_ecc,                  
input            [7:0]  epl0_igr1_rx_ecc,                         
input            [2:0]  epl0_igr1_rx_flow_control_tc,             
input           [23:0]  epl0_igr1_rx_metadata,                    
input                   epl0_igr1_rx_pfc_xoff,                    
input            [1:0]  epl0_igr1_rx_port_num,                    
input           [35:0]  epl0_igr1_rx_time_stamp,                  
input            [7:0]  epl1_igr0_rx_data_valid,                  
input         [0:7][71:0]  epl1_igr0_rx_data_w_ecc,                  
input            [7:0]  epl1_igr0_rx_ecc,                         
input            [2:0]  epl1_igr0_rx_flow_control_tc,             
input           [23:0]  epl1_igr0_rx_metadata,                    
input                   epl1_igr0_rx_pfc_xoff,                    
input            [1:0]  epl1_igr0_rx_port_num,                    
input           [35:0]  epl1_igr0_rx_time_stamp,                  
input            [7:0]  epl1_igr1_rx_data_valid,                  
input         [0:7][71:0]  epl1_igr1_rx_data_w_ecc,                  
input            [7:0]  epl1_igr1_rx_ecc,                         
input            [2:0]  epl1_igr1_rx_flow_control_tc,             
input           [23:0]  epl1_igr1_rx_metadata,                    
input                   epl1_igr1_rx_pfc_xoff,                    
input            [1:0]  epl1_igr1_rx_port_num,                    
input           [35:0]  epl1_igr1_rx_time_stamp,                  
input            [7:0]  epl2_igr0_rx_data_valid,                  
input         [0:7][71:0]  epl2_igr0_rx_data_w_ecc,                  
input            [7:0]  epl2_igr0_rx_ecc,                         
input            [2:0]  epl2_igr0_rx_flow_control_tc,             
input           [23:0]  epl2_igr0_rx_metadata,                    
input                   epl2_igr0_rx_pfc_xoff,                    
input            [1:0]  epl2_igr0_rx_port_num,                    
input           [35:0]  epl2_igr0_rx_time_stamp,                  
input            [7:0]  epl2_igr1_rx_data_valid,                  
input         [0:7][71:0]  epl2_igr1_rx_data_w_ecc,                  
input            [7:0]  epl2_igr1_rx_ecc,                         
input            [2:0]  epl2_igr1_rx_flow_control_tc,             
input           [23:0]  epl2_igr1_rx_metadata,                    
input                   epl2_igr1_rx_pfc_xoff,                    
input            [1:0]  epl2_igr1_rx_port_num,                    
input           [35:0]  epl2_igr1_rx_time_stamp,                  
input            [7:0]  epl3_igr0_rx_data_valid,                  
input         [0:7][71:0]  epl3_igr0_rx_data_w_ecc,                  
input            [7:0]  epl3_igr0_rx_ecc,                         
input            [2:0]  epl3_igr0_rx_flow_control_tc,             
input           [23:0]  epl3_igr0_rx_metadata,                    
input                   epl3_igr0_rx_pfc_xoff,                    
input            [1:0]  epl3_igr0_rx_port_num,                    
input           [35:0]  epl3_igr0_rx_time_stamp,                  
input            [7:0]  epl3_igr1_rx_data_valid,                  
input         [0:7][71:0]  epl3_igr1_rx_data_w_ecc,                  
input            [7:0]  epl3_igr1_rx_ecc,                         
input            [2:0]  epl3_igr1_rx_flow_control_tc,             
input           [23:0]  epl3_igr1_rx_metadata,                    
input                   epl3_igr1_rx_pfc_xoff,                    
input            [1:0]  epl3_igr1_rx_port_num,                    
input           [35:0]  epl3_igr1_rx_time_stamp,                  
input           [19:0]  igr0_vp_cpp_rx_metadata,                  
input            [7:0]  igr0_vp_rx_data_valid,                    
input         [0:7][71:0]  igr0_vp_rx_data_w_ecc,                    
input            [7:0]  igr0_vp_rx_ecc,                           
input            [2:0]  igr0_vp_rx_flow_control_tc,               
input           [23:0]  igr0_vp_rx_metadata,                      
input            [1:0]  igr0_vp_rx_port_num,                      
input           [35:0]  igr0_vp_rx_time_stamp,                    
input           [19:0]  igr1_vp_cpp_rx_metadata,                  
input            [7:0]  igr1_vp_rx_data_valid,                    
input         [0:7][71:0]  igr1_vp_rx_data_w_ecc,                    
input            [7:0]  igr1_vp_rx_ecc,                           
input            [2:0]  igr1_vp_rx_flow_control_tc,               
input           [23:0]  igr1_vp_rx_metadata,                      
input            [1:0]  igr1_vp_rx_port_num,                      
input           [35:0]  igr1_vp_rx_time_stamp,                    
input                   reset,                                    
input                   rst_n,                                    //taken from HLP active low for MBY?  

//Interface List
ahb_rx_ppe_if.ppe                 ahb0_rx_ppe_if,  
ahb_rx_ppe_if.ppe                 ahb0_txppe0_if,  
ahb_rx_ppe_if.ppe                 ahb0_txppe1_if,  
ahb_rx_ppe_if.ppe                 ahb1_rx_ppe_if,  
ahb_rx_ppe_if.ppe                 ahb1_txppe0_if,  
ahb_rx_ppe_if.ppe                 ahb1_txppe1_if,  
egr_ahb_if.egr                    egr0_ahb_if,  //EGR-AHB and DFx Interface  
egr_mc_table_if.egr               egr0_mc_table_if0,  //EGR-MultiCast Shared Table 0 Interface  
egr_mc_table_if.egr               egr0_mc_table_if1,  //EGR-MultiCast Shared Table 1 Interface  
egr_pod_if.egr                    egr0_pod_if,  //EGR-Pod Ring Interface  
egr_ppe_stm_if.egr                egr0_ppestm_if0,  //EGR-PPE Shared Table Memory 0 Interface   
egr_ppe_stm_if.egr                egr0_ppestm_if1,  //EGR-PPE Shared Table Memory 1 Interface  
egr_smm_readarb_if.egr            egr0_smm_readarb_if,  //EGR-SMM_Read_Arb Interface  
egr_smm_writearb_if.egr           egr0_smm_writearb_if,  //EGR-SMM_Write_Arb Interface  
egr_statsmgmt_if.egr              egr0_statsmgmt_if,  //EGR-Stats Management Interface  
egr_tagring_if.egr                egr0_tagring_if,  //EGR-Tag Ring Interface  
egr_vp_if.egr                     egr0_vp_if0,  //EGR-VP0 Interface  
egr_vp_if.egr                     egr0_vp_if1,  //EGR-VP1 Interface  
egr_ahb_if.egr                    egr1_ahb_if,  //EGR-AHB and DFx Interface  
egr_mc_table_if.egr               egr1_mc_table_if0,  //EGR-MultiCast Shared Table 0 Interface  
egr_mc_table_if.egr               egr1_mc_table_if1,  //EGR-MultiCast Shared Table 1 Interface  
egr_pod_if.egr                    egr1_pod_if,  //EGR-Pod Ring Interface  
egr_ppe_stm_if.egr                egr1_ppestm_if0,  //EGR-PPE Shared Table Memory 0 Interface   
egr_ppe_stm_if.egr                egr1_ppestm_if1,  //EGR-PPE Shared Table Memory 1 Interface  
egr_smm_readarb_if.egr            egr1_smm_readarb_if,  //EGR-SMM_Read_Arb Interface  
egr_smm_writearb_if.egr           egr1_smm_writearb_if,  //EGR-SMM_Write_Arb Interface  
egr_statsmgmt_if.egr              egr1_statsmgmt_if,  //EGR-Stats Management Interface  
egr_tagring_if.egr                egr1_tagring_if,  //EGR-Tag Ring Interface  
egr_vp_if.egr                     egr1_vp_if0,  //EGR-VP0 Interface  
egr_vp_if.egr                     egr1_vp_if1,  //EGR-VP1 Interface  
egr_ppe_stm_if.stm                egr_ppe_stm_if,  
glb_rx_ppe_if.ppe                 glb0_rx_ppe_if,  
glb_rx_ppe_if.ppe                 glb0_txppe0_if,  
glb_rx_ppe_if.ppe                 glb0_txppe1_if,  
glb_rx_ppe_if.ppe                 glb1_rx_ppe_if,  
glb_rx_ppe_if.ppe                 glb1_txppe0_if,  
glb_rx_ppe_if.ppe                 glb1_txppe1_if,  

//Output List
output                  igr0_vp_tx_pfc_xoff,                      //FIXME should this be [1:0] for 2 VP   
output                  igr1_vp_tx_pfc_xoff                       //FIXME should this be [1:0] for 2 VP   
);

egr_epl_if                       egr_();
egr_igr_if                       egr_igr_if();
rx_ppe_ppe_stm_if                rx_ppe_ppe_stm_if();


// module mgp0    from mgp using mgp.map 0
mgp    mgp0(
/* input  logic                      */ .arst_n                       (arst_n),                                 //Asynchronous negedge reset     
/* input  logic                      */ .cclk                         (cclk),                                   
/* input  logic                      */ .clk                          (clk),                                    
/* input  logic                [7:0] */ .epl0_igr_rx_data_valid       (epl0_igr0_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl0_igr_rx_data_w_ecc       (epl0_igr0_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl0_igr_rx_ecc              (epl0_igr0_rx_ecc),                       
/* input  logic                [2:0] */ .epl0_igr_rx_flow_control_tc  (epl0_igr0_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl0_igr_rx_metadata         (epl0_igr0_rx_metadata),                  
/* input  logic                      */ .epl0_igr_rx_pfc_xoff         (epl0_igr0_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl0_igr_rx_port_num         (epl0_igr0_rx_port_num),                  
/* input  logic               [35:0] */ .epl0_igr_rx_time_stamp       (epl0_igr0_rx_time_stamp),                
/* input  logic                [7:0] */ .epl1_igr_rx_data_valid       (epl1_igr0_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl1_igr_rx_data_w_ecc       (epl1_igr0_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl1_igr_rx_ecc              (epl1_igr0_rx_ecc),                       
/* input  logic                [2:0] */ .epl1_igr_rx_flow_control_tc  (epl1_igr0_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl1_igr_rx_metadata         (epl1_igr0_rx_metadata),                  
/* input  logic                      */ .epl1_igr_rx_pfc_xoff         (epl1_igr0_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl1_igr_rx_port_num         (epl1_igr0_rx_port_num),                  
/* input  logic               [35:0] */ .epl1_igr_rx_time_stamp       (epl1_igr0_rx_time_stamp),                
/* input  logic                [7:0] */ .epl2_igr_rx_data_valid       (epl2_igr0_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl2_igr_rx_data_w_ecc       (epl2_igr0_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl2_igr_rx_ecc              (epl2_igr0_rx_ecc),                       
/* input  logic                [2:0] */ .epl2_igr_rx_flow_control_tc  (epl2_igr0_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl2_igr_rx_metadata         (epl2_igr0_rx_metadata),                  
/* input  logic                      */ .epl2_igr_rx_pfc_xoff         (epl2_igr0_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl2_igr_rx_port_num         (epl2_igr0_rx_port_num),                  
/* input  logic               [35:0] */ .epl2_igr_rx_time_stamp       (epl2_igr0_rx_time_stamp),                
/* input  logic                [7:0] */ .epl3_igr_rx_data_valid       (epl3_igr0_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl3_igr_rx_data_w_ecc       (epl3_igr0_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl3_igr_rx_ecc              (epl3_igr0_rx_ecc),                       
/* input  logic                [2:0] */ .epl3_igr_rx_flow_control_tc  (epl3_igr0_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl3_igr_rx_metadata         (epl3_igr0_rx_metadata),                  
/* input  logic                      */ .epl3_igr_rx_pfc_xoff         (epl3_igr0_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl3_igr_rx_port_num         (epl3_igr0_rx_port_num),                  
/* input  logic               [35:0] */ .epl3_igr_rx_time_stamp       (epl3_igr0_rx_time_stamp),                
/* input  logic               [19:0] */ .igr_vp_cpp_rx_metadata       (igr0_vp_cpp_rx_metadata),                
/* input  logic                [7:0] */ .igr_vp_rx_data_valid         (igr0_vp_rx_data_valid),                  
/* input  logic          [0:7][71:0] */ .igr_vp_rx_data_w_ecc         (igr0_vp_rx_data_w_ecc),                  
/* input  logic                [7:0] */ .igr_vp_rx_ecc                (igr0_vp_rx_ecc),                         
/* input  logic                [2:0] */ .igr_vp_rx_flow_control_tc    (igr0_vp_rx_flow_control_tc),             
/* input  logic               [23:0] */ .igr_vp_rx_metadata           (igr0_vp_rx_metadata),                    
/* input  logic                [1:0] */ .igr_vp_rx_port_num           (igr0_vp_rx_port_num),                    
/* input  logic               [35:0] */ .igr_vp_rx_time_stamp         (igr0_vp_rx_time_stamp),                  
/* input  logic                      */ .reset                        (reset),                                  
/* input  logic                      */ .rst_n                        (rst_n),                                  //taken from HLP active low for MBY?  
/* Interface ahb_rx_ppe_if.ppe       */ .ahb_rx_ppe_if                (ahb0_rx_ppe_if),                         
/* Interface ahb_rx_ppe_if.ppe       */ .ahb_txppe0_if                (ahb0_txppe0_if),                         
/* Interface ahb_rx_ppe_if.ppe       */ .ahb_txppe1_if                (ahb0_txppe1_if),                         
/* Interface egr_ahb_if.egr          */ .egr_ahb_if                   (egr0_ahb_if),                            
/* Interface egr_epl_if.egr          */ .egr_epl0_if                  (egr_),                                   
/* Interface egr_epl_if.egr          */ .egr_epl1_if                  (egr_),                                   
/* Interface egr_epl_if.egr          */ .egr_epl2_if                  (egr_),                                   
/* Interface egr_epl_if.egr          */ .egr_epl3_if                  (egr_),                                   
/* Interface egr_igr_if.egr          */ .egr_igr_if                   (egr_igr_if),                             
/* Interface egr_mc_table_if.egr     */ .egr_mc_table_if0             (egr0_mc_table_if0),                      
/* Interface egr_mc_table_if.egr     */ .egr_mc_table_if1             (egr0_mc_table_if1),                      
/* Interface egr_pod_if.egr          */ .egr_pod_if                   (egr0_pod_if),                            
/* Interface egr_ppe_stm_if.egr      */ .egr_ppestm_if0               (egr0_ppestm_if0),                        
/* Interface egr_ppe_stm_if.egr      */ .egr_ppestm_if1               (egr0_ppestm_if1),                        
/* Interface egr_smm_readarb_if.egr  */ .egr_smm_readarb_if           (egr0_smm_readarb_if),                    
/* Interface egr_smm_writearb_if.egr */ .egr_smm_writearb_if          (egr0_smm_writearb_if),                   
/* Interface egr_statsmgmt_if.egr    */ .egr_statsmgmt_if             (egr0_statsmgmt_if),                      
/* Interface egr_tagring_if.egr      */ .egr_tagring_if               (egr0_tagring_if),                        
/* Interface egr_vp_if.egr           */ .egr_vp_if0                   (egr0_vp_if0),                            
/* Interface egr_vp_if.egr           */ .egr_vp_if1                   (egr0_vp_if1),                            
/* Interface glb_rx_ppe_if.ppe       */ .glb_rx_ppe_if                (glb0_rx_ppe_if),                         
/* Interface glb_rx_ppe_if.ppe       */ .glb_txppe0_if                (glb0_txppe0_if),                         
/* Interface glb_rx_ppe_if.ppe       */ .glb_txppe1_if                (glb0_txppe1_if),                         
/* Interface rx_ppe_ppe_stm_if.ppe   */ .rx_ppe_ppe_stm_if            (rx_ppe_ppe_stm_if),                      
/* output logic                      */ .igr_vp_tx_pfc_xoff           (igr0_vp_tx_pfc_xoff));                    //FIXME should this be [1:0] for 2 VP   
// End of module mgp0 from mgp


// module mgp1    from mgp using mgp.map 1
mgp    mgp1(
/* input  logic                      */ .arst_n                       (arst_n),                                 //Asynchronous negedge reset     
/* input  logic                      */ .cclk                         (cclk),                                   
/* input  logic                      */ .clk                          (clk),                                    
/* input  logic                [7:0] */ .epl0_igr_rx_data_valid       (epl0_igr1_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl0_igr_rx_data_w_ecc       (epl0_igr1_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl0_igr_rx_ecc              (epl0_igr1_rx_ecc),                       
/* input  logic                [2:0] */ .epl0_igr_rx_flow_control_tc  (epl0_igr1_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl0_igr_rx_metadata         (epl0_igr1_rx_metadata),                  
/* input  logic                      */ .epl0_igr_rx_pfc_xoff         (epl0_igr1_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl0_igr_rx_port_num         (epl0_igr1_rx_port_num),                  
/* input  logic               [35:0] */ .epl0_igr_rx_time_stamp       (epl0_igr1_rx_time_stamp),                
/* input  logic                [7:0] */ .epl1_igr_rx_data_valid       (epl1_igr1_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl1_igr_rx_data_w_ecc       (epl1_igr1_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl1_igr_rx_ecc              (epl1_igr1_rx_ecc),                       
/* input  logic                [2:0] */ .epl1_igr_rx_flow_control_tc  (epl1_igr1_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl1_igr_rx_metadata         (epl1_igr1_rx_metadata),                  
/* input  logic                      */ .epl1_igr_rx_pfc_xoff         (epl1_igr1_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl1_igr_rx_port_num         (epl1_igr1_rx_port_num),                  
/* input  logic               [35:0] */ .epl1_igr_rx_time_stamp       (epl1_igr1_rx_time_stamp),                
/* input  logic                [7:0] */ .epl2_igr_rx_data_valid       (epl2_igr1_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl2_igr_rx_data_w_ecc       (epl2_igr1_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl2_igr_rx_ecc              (epl2_igr1_rx_ecc),                       
/* input  logic                [2:0] */ .epl2_igr_rx_flow_control_tc  (epl2_igr1_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl2_igr_rx_metadata         (epl2_igr1_rx_metadata),                  
/* input  logic                      */ .epl2_igr_rx_pfc_xoff         (epl2_igr1_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl2_igr_rx_port_num         (epl2_igr1_rx_port_num),                  
/* input  logic               [35:0] */ .epl2_igr_rx_time_stamp       (epl2_igr1_rx_time_stamp),                
/* input  logic                [7:0] */ .epl3_igr_rx_data_valid       (epl3_igr1_rx_data_valid),                
/* input  logic          [0:7][71:0] */ .epl3_igr_rx_data_w_ecc       (epl3_igr1_rx_data_w_ecc),                
/* input  logic                [7:0] */ .epl3_igr_rx_ecc              (epl3_igr1_rx_ecc),                       
/* input  logic                [2:0] */ .epl3_igr_rx_flow_control_tc  (epl3_igr1_rx_flow_control_tc),           
/* input  logic               [23:0] */ .epl3_igr_rx_metadata         (epl3_igr1_rx_metadata),                  
/* input  logic                      */ .epl3_igr_rx_pfc_xoff         (epl3_igr1_rx_pfc_xoff),                  
/* input  logic                [1:0] */ .epl3_igr_rx_port_num         (epl3_igr1_rx_port_num),                  
/* input  logic               [35:0] */ .epl3_igr_rx_time_stamp       (epl3_igr1_rx_time_stamp),                
/* input  logic               [19:0] */ .igr_vp_cpp_rx_metadata       (igr1_vp_cpp_rx_metadata),                
/* input  logic                [7:0] */ .igr_vp_rx_data_valid         (igr1_vp_rx_data_valid),                  
/* input  logic          [0:7][71:0] */ .igr_vp_rx_data_w_ecc         (igr1_vp_rx_data_w_ecc),                  
/* input  logic                [7:0] */ .igr_vp_rx_ecc                (igr1_vp_rx_ecc),                         
/* input  logic                [2:0] */ .igr_vp_rx_flow_control_tc    (igr1_vp_rx_flow_control_tc),             
/* input  logic               [23:0] */ .igr_vp_rx_metadata           (igr1_vp_rx_metadata),                    
/* input  logic                [1:0] */ .igr_vp_rx_port_num           (igr1_vp_rx_port_num),                    
/* input  logic               [35:0] */ .igr_vp_rx_time_stamp         (igr1_vp_rx_time_stamp),                  
/* input  logic                      */ .reset                        (reset),                                  
/* input  logic                      */ .rst_n                        (rst_n),                                  //taken from HLP active low for MBY?  
/* Interface ahb_rx_ppe_if.ppe       */ .ahb_rx_ppe_if                (ahb1_rx_ppe_if),                         
/* Interface ahb_rx_ppe_if.ppe       */ .ahb_txppe0_if                (ahb1_txppe0_if),                         
/* Interface ahb_rx_ppe_if.ppe       */ .ahb_txppe1_if                (ahb1_txppe1_if),                         
/* Interface egr_ahb_if.egr          */ .egr_ahb_if                   (egr1_ahb_if),                            
/* Interface egr_epl_if.egr          */ .egr_epl0_if                  (egr_),                                   
/* Interface egr_epl_if.egr          */ .egr_epl1_if                  (egr_),                                   
/* Interface egr_epl_if.egr          */ .egr_epl2_if                  (egr_),                                   
/* Interface egr_epl_if.egr          */ .egr_epl3_if                  (egr_),                                   
/* Interface egr_igr_if.egr          */ .egr_igr_if                   (egr_igr_if),                             
/* Interface egr_mc_table_if.egr     */ .egr_mc_table_if0             (egr1_mc_table_if0),                      
/* Interface egr_mc_table_if.egr     */ .egr_mc_table_if1             (egr1_mc_table_if1),                      
/* Interface egr_pod_if.egr          */ .egr_pod_if                   (egr1_pod_if),                            
/* Interface egr_ppe_stm_if.egr      */ .egr_ppestm_if0               (egr1_ppestm_if0),                        
/* Interface egr_ppe_stm_if.egr      */ .egr_ppestm_if1               (egr1_ppestm_if1),                        
/* Interface egr_smm_readarb_if.egr  */ .egr_smm_readarb_if           (egr1_smm_readarb_if),                    
/* Interface egr_smm_writearb_if.egr */ .egr_smm_writearb_if          (egr1_smm_writearb_if),                   
/* Interface egr_statsmgmt_if.egr    */ .egr_statsmgmt_if             (egr1_statsmgmt_if),                      
/* Interface egr_tagring_if.egr      */ .egr_tagring_if               (egr1_tagring_if),                        
/* Interface egr_vp_if.egr           */ .egr_vp_if0                   (egr1_vp_if0),                            
/* Interface egr_vp_if.egr           */ .egr_vp_if1                   (egr1_vp_if1),                            
/* Interface glb_rx_ppe_if.ppe       */ .glb_rx_ppe_if                (glb1_rx_ppe_if),                         
/* Interface glb_rx_ppe_if.ppe       */ .glb_txppe0_if                (glb1_txppe0_if),                         
/* Interface glb_rx_ppe_if.ppe       */ .glb_txppe1_if                (glb1_txppe1_if),                         
/* Interface rx_ppe_ppe_stm_if.ppe   */ .rx_ppe_ppe_stm_if            (rx_ppe_ppe_stm_if),                      
/* output logic                      */ .igr_vp_tx_pfc_xoff           (igr1_vp_tx_pfc_xoff));                    //FIXME should this be [1:0] for 2 VP   
// End of module mgp1 from mgp


// module ppestm    from ppe_stm_top using ppestm.map 
ppe_stm_top    ppestm(
/* input  logic                    */ .reset                        (reset),                                  
/* Interface rx_ppe_ppe_stm_if.stm */ .rx_ppe_ppe_stm_if            (rx_ppe_ppe_stm_if),                      
/* Interface egr_ppe_stm_if.stm    */ .egr_ppe_stm_if               (egr_ppe_stm_if),                         
/* input  logic                    */ .cclk                         (cclk));                                   
// End of module ppestm from ppe_stm_top

endmodule // mpp
