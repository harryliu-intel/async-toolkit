///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cm_apply_map_pkg.vh                                
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_CM_APPLY_MAP_PKG_VH
`define MBY_PPE_CM_APPLY_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_cm_apply_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_cm_apply_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_cm_apply_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_cm_apply_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [61:0] reserved0;  // RSVD
    logic  [0:0] SOFT_DROP_ON_PRIVATE;  // RW
    logic  [0:0] SOFT_DROP_ON_SMP_FREE;  // RW
} CM_APPLY_TX_SOFTDROP_CFG_t;

localparam CM_APPLY_TX_SOFTDROP_CFG_REG_STRIDE = 48'h8;
localparam CM_APPLY_TX_SOFTDROP_CFG_REG_ENTRIES = 8;
localparam CM_APPLY_TX_SOFTDROP_CFG_REGFILE_STRIDE = 48'h40;
localparam CM_APPLY_TX_SOFTDROP_CFG_REGFILE_ENTRIES = 64;
localparam CM_APPLY_TX_SOFTDROP_CFG_CR_ADDR = 48'h0;
localparam CM_APPLY_TX_SOFTDROP_CFG_SIZE = 64;
localparam CM_APPLY_TX_SOFTDROP_CFG_SOFT_DROP_ON_PRIVATE_LO = 1;
localparam CM_APPLY_TX_SOFTDROP_CFG_SOFT_DROP_ON_PRIVATE_HI = 1;
localparam CM_APPLY_TX_SOFTDROP_CFG_SOFT_DROP_ON_PRIVATE_RESET = 1'h0;
localparam CM_APPLY_TX_SOFTDROP_CFG_SOFT_DROP_ON_SMP_FREE_LO = 0;
localparam CM_APPLY_TX_SOFTDROP_CFG_SOFT_DROP_ON_SMP_FREE_HI = 0;
localparam CM_APPLY_TX_SOFTDROP_CFG_SOFT_DROP_ON_SMP_FREE_RESET = 1'h0;
localparam CM_APPLY_TX_SOFTDROP_CFG_USEMASK = 64'h3;
localparam CM_APPLY_TX_SOFTDROP_CFG_RO_MASK = 64'h0;
localparam CM_APPLY_TX_SOFTDROP_CFG_WO_MASK = 64'h0;
localparam CM_APPLY_TX_SOFTDROP_CFG_RESET = 64'h0;

typedef struct packed {
    logic [44:0] reserved0;  // RSVD
    logic [14:0] QUEUE_DEPTH;  // RO/V
    logic  [0:0] OVER_SMP_FREE2;  // RO/V
    logic  [0:0] OVER_SMP_FREE;  // RO/V
    logic  [0:0] TX_HOG;  // RO/V
    logic  [0:0] TX_PRIVATE;  // RO/V
} CM_APPLY_TX_TC_STATE_t;

localparam CM_APPLY_TX_TC_STATE_REG_STRIDE = 48'h8;
localparam CM_APPLY_TX_TC_STATE_REG_ENTRIES = 8;
localparam CM_APPLY_TX_TC_STATE_REGFILE_STRIDE = 48'h40;
localparam CM_APPLY_TX_TC_STATE_REGFILE_ENTRIES = 64;
localparam CM_APPLY_TX_TC_STATE_CR_ADDR = 48'h1000;
localparam CM_APPLY_TX_TC_STATE_SIZE = 64;
localparam CM_APPLY_TX_TC_STATE_QUEUE_DEPTH_LO = 4;
localparam CM_APPLY_TX_TC_STATE_QUEUE_DEPTH_HI = 18;
localparam CM_APPLY_TX_TC_STATE_QUEUE_DEPTH_RESET = 15'h0;
localparam CM_APPLY_TX_TC_STATE_OVER_SMP_FREE2_LO = 3;
localparam CM_APPLY_TX_TC_STATE_OVER_SMP_FREE2_HI = 3;
localparam CM_APPLY_TX_TC_STATE_OVER_SMP_FREE2_RESET = 1'h0;
localparam CM_APPLY_TX_TC_STATE_OVER_SMP_FREE_LO = 2;
localparam CM_APPLY_TX_TC_STATE_OVER_SMP_FREE_HI = 2;
localparam CM_APPLY_TX_TC_STATE_OVER_SMP_FREE_RESET = 1'h0;
localparam CM_APPLY_TX_TC_STATE_TX_HOG_LO = 1;
localparam CM_APPLY_TX_TC_STATE_TX_HOG_HI = 1;
localparam CM_APPLY_TX_TC_STATE_TX_HOG_RESET = 1'h0;
localparam CM_APPLY_TX_TC_STATE_TX_PRIVATE_LO = 0;
localparam CM_APPLY_TX_TC_STATE_TX_PRIVATE_HI = 0;
localparam CM_APPLY_TX_TC_STATE_TX_PRIVATE_RESET = 1'h0;
localparam CM_APPLY_TX_TC_STATE_USEMASK = 64'h7FFFF;
localparam CM_APPLY_TX_TC_STATE_RO_MASK = 64'h7FFFF;
localparam CM_APPLY_TX_TC_STATE_WO_MASK = 64'h0;
localparam CM_APPLY_TX_TC_STATE_RESET = 64'h0;

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic [14:0] WM_THRESHOLD;  // RW
} CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t;

localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_REG_STRIDE = 48'h8;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_REG_ENTRIES = 8;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_REGFILE_STRIDE = 48'h40;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_REGFILE_ENTRIES = 64;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_CR_ADDR = 48'h2000;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_SIZE = 64;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_WM_THRESHOLD_LO = 0;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_WM_THRESHOLD_HI = 14;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_WM_THRESHOLD_RESET = 15'h0;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_USEMASK = 64'h7FFF;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_RO_MASK = 64'h0;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_WO_MASK = 64'h0;
localparam CM_APPLY_TX_TC_QCN_WM_THRESHOLD_RESET = 64'h0;

typedef struct packed {
    logic [61:0] reserved0;  // RSVD
    logic  [0:0] RX_HOG;  // RO/V
    logic  [0:0] RX_PRIVATE;  // RO/V
} CM_APPLY_RX_SMP_STATE_t;

localparam CM_APPLY_RX_SMP_STATE_REG_STRIDE = 48'h8;
localparam CM_APPLY_RX_SMP_STATE_REG_ENTRIES = 2;
localparam CM_APPLY_RX_SMP_STATE_REGFILE_STRIDE = 48'h10;
localparam CM_APPLY_RX_SMP_STATE_REGFILE_ENTRIES = 32;
localparam CM_APPLY_RX_SMP_STATE_CR_ADDR = 48'h3000;
localparam CM_APPLY_RX_SMP_STATE_SIZE = 64;
localparam CM_APPLY_RX_SMP_STATE_RX_HOG_LO = 1;
localparam CM_APPLY_RX_SMP_STATE_RX_HOG_HI = 1;
localparam CM_APPLY_RX_SMP_STATE_RX_HOG_RESET = 1'h0;
localparam CM_APPLY_RX_SMP_STATE_RX_PRIVATE_LO = 0;
localparam CM_APPLY_RX_SMP_STATE_RX_PRIVATE_HI = 0;
localparam CM_APPLY_RX_SMP_STATE_RX_PRIVATE_RESET = 1'h0;
localparam CM_APPLY_RX_SMP_STATE_USEMASK = 64'h3;
localparam CM_APPLY_RX_SMP_STATE_RO_MASK = 64'h3;
localparam CM_APPLY_RX_SMP_STATE_WO_MASK = 64'h0;
localparam CM_APPLY_RX_SMP_STATE_RESET = 64'h0;

typedef struct packed {
    logic [58:0] reserved0;  // RSVD
    logic  [4:0] PORT;  // RW
} CM_APPLY_MIRROR_PROFILE_TABLE_t;

localparam CM_APPLY_MIRROR_PROFILE_TABLE_REG_STRIDE = 48'h8;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_REG_ENTRIES = 64;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_CR_ADDR = 48'h3200;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_SIZE = 64;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_PORT_LO = 0;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_PORT_HI = 4;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_PORT_RESET = 5'h0;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_USEMASK = 64'h1F;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_RO_MASK = 64'h0;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_WO_MASK = 64'h0;
localparam CM_APPLY_MIRROR_PROFILE_TABLE_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] FRAMES;  // RW/V
} CM_APPLY_DROP_COUNT_t;

localparam CM_APPLY_DROP_COUNT_REG_STRIDE = 48'h8;
localparam CM_APPLY_DROP_COUNT_REG_ENTRIES = 32;
localparam CM_APPLY_DROP_COUNT_CR_ADDR = 48'h3400;
localparam CM_APPLY_DROP_COUNT_SIZE = 64;
localparam CM_APPLY_DROP_COUNT_FRAMES_LO = 0;
localparam CM_APPLY_DROP_COUNT_FRAMES_HI = 47;
localparam CM_APPLY_DROP_COUNT_FRAMES_RESET = 48'h0;
localparam CM_APPLY_DROP_COUNT_USEMASK = 64'hFFFFFFFFFFFF;
localparam CM_APPLY_DROP_COUNT_RO_MASK = 64'h0;
localparam CM_APPLY_DROP_COUNT_WO_MASK = 64'h0;
localparam CM_APPLY_DROP_COUNT_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [15:0] GLORT_MASK;  // RW
    logic [15:0] GLORT;  // RW
} CM_APPLY_LOOPBACK_SUPPRESS_t;

localparam CM_APPLY_LOOPBACK_SUPPRESS_REG_STRIDE = 48'h8;
localparam CM_APPLY_LOOPBACK_SUPPRESS_REG_ENTRIES = 32;
localparam CM_APPLY_LOOPBACK_SUPPRESS_CR_ADDR = 48'h3500;
localparam CM_APPLY_LOOPBACK_SUPPRESS_SIZE = 64;
localparam CM_APPLY_LOOPBACK_SUPPRESS_GLORT_MASK_LO = 16;
localparam CM_APPLY_LOOPBACK_SUPPRESS_GLORT_MASK_HI = 31;
localparam CM_APPLY_LOOPBACK_SUPPRESS_GLORT_MASK_RESET = 16'h0;
localparam CM_APPLY_LOOPBACK_SUPPRESS_GLORT_LO = 0;
localparam CM_APPLY_LOOPBACK_SUPPRESS_GLORT_HI = 15;
localparam CM_APPLY_LOOPBACK_SUPPRESS_GLORT_RESET = 16'hffff;
localparam CM_APPLY_LOOPBACK_SUPPRESS_USEMASK = 64'hFFFFFFFF;
localparam CM_APPLY_LOOPBACK_SUPPRESS_RO_MASK = 64'h0;
localparam CM_APPLY_LOOPBACK_SUPPRESS_WO_MASK = 64'h0;
localparam CM_APPLY_LOOPBACK_SUPPRESS_RESET = 64'hFFFF;

typedef struct packed {
    logic [60:0] reserved0;  // RSVD
    logic  [2:0] JITTER_BITS;  // RW
} CM_APPLY_SOFTDROP_CFG_t;

localparam CM_APPLY_SOFTDROP_CFG_REG_STRIDE = 48'h8;
localparam CM_APPLY_SOFTDROP_CFG_REG_ENTRIES = 8;
localparam CM_APPLY_SOFTDROP_CFG_CR_ADDR = 48'h3600;
localparam CM_APPLY_SOFTDROP_CFG_SIZE = 64;
localparam CM_APPLY_SOFTDROP_CFG_JITTER_BITS_LO = 0;
localparam CM_APPLY_SOFTDROP_CFG_JITTER_BITS_HI = 2;
localparam CM_APPLY_SOFTDROP_CFG_JITTER_BITS_RESET = 3'h0;
localparam CM_APPLY_SOFTDROP_CFG_USEMASK = 64'h7;
localparam CM_APPLY_SOFTDROP_CFG_RO_MASK = 64'h0;
localparam CM_APPLY_SOFTDROP_CFG_WO_MASK = 64'h0;
localparam CM_APPLY_SOFTDROP_CFG_RESET = 64'h0;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [0:0] OVER_LIMIT;  // RO/V
    logic  [7:0] USAGE_OVER_LIMIT;  // RO/V
} CM_APPLY_SOFTDROP_STATE_t;

localparam CM_APPLY_SOFTDROP_STATE_REG_STRIDE = 48'h8;
localparam CM_APPLY_SOFTDROP_STATE_REG_ENTRIES = 8;
localparam CM_APPLY_SOFTDROP_STATE_CR_ADDR = 48'h3640;
localparam CM_APPLY_SOFTDROP_STATE_SIZE = 64;
localparam CM_APPLY_SOFTDROP_STATE_OVER_LIMIT_LO = 8;
localparam CM_APPLY_SOFTDROP_STATE_OVER_LIMIT_HI = 8;
localparam CM_APPLY_SOFTDROP_STATE_OVER_LIMIT_RESET = 1'h0;
localparam CM_APPLY_SOFTDROP_STATE_USAGE_OVER_LIMIT_LO = 0;
localparam CM_APPLY_SOFTDROP_STATE_USAGE_OVER_LIMIT_HI = 7;
localparam CM_APPLY_SOFTDROP_STATE_USAGE_OVER_LIMIT_RESET = 8'h0;
localparam CM_APPLY_SOFTDROP_STATE_USEMASK = 64'h1FF;
localparam CM_APPLY_SOFTDROP_STATE_RO_MASK = 64'h1FF;
localparam CM_APPLY_SOFTDROP_STATE_WO_MASK = 64'h0;
localparam CM_APPLY_SOFTDROP_STATE_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] TRAP_GLORT;  // RW
} CM_APPLY_TRAP_GLORT_t;

localparam CM_APPLY_TRAP_GLORT_REG_STRIDE = 48'h8;
localparam CM_APPLY_TRAP_GLORT_REG_ENTRIES = 16;
localparam [15:0][47:0] CM_APPLY_TRAP_GLORT_CR_ADDR = {48'h36F8, 48'h36F0, 48'h36E8, 48'h36E0, 48'h36D8, 48'h36D0, 48'h36C8, 48'h36C0, 48'h36B8, 48'h36B0, 48'h36A8, 48'h36A0, 48'h3698, 48'h3690, 48'h3688, 48'h3680};
localparam CM_APPLY_TRAP_GLORT_SIZE = 64;
localparam CM_APPLY_TRAP_GLORT_TRAP_GLORT_LO = 0;
localparam CM_APPLY_TRAP_GLORT_TRAP_GLORT_HI = 15;
localparam CM_APPLY_TRAP_GLORT_TRAP_GLORT_RESET = 16'h0;
localparam CM_APPLY_TRAP_GLORT_USEMASK = 64'hFFFF;
localparam CM_APPLY_TRAP_GLORT_RO_MASK = 64'h0;
localparam CM_APPLY_TRAP_GLORT_WO_MASK = 64'h0;
localparam CM_APPLY_TRAP_GLORT_RESET = 64'h0;

typedef struct packed {
    logic [55:0] reserved0;  // RSVD
    logic  [0:0] SMP_7;  // RW
    logic  [0:0] SMP_6;  // RW
    logic  [0:0] SMP_5;  // RW
    logic  [0:0] SMP_4;  // RW
    logic  [0:0] SMP_3;  // RW
    logic  [0:0] SMP_2;  // RW
    logic  [0:0] SMP_1;  // RW
    logic  [0:0] SMP_0;  // RW
} CM_APPLY_TC_TO_SMP_t;

localparam CM_APPLY_TC_TO_SMP_REG_STRIDE = 48'h8;
localparam CM_APPLY_TC_TO_SMP_REG_ENTRIES = 1;
localparam [47:0] CM_APPLY_TC_TO_SMP_CR_ADDR = 48'h3700;
localparam CM_APPLY_TC_TO_SMP_SIZE = 64;
localparam CM_APPLY_TC_TO_SMP_SMP_7_LO = 7;
localparam CM_APPLY_TC_TO_SMP_SMP_7_HI = 7;
localparam CM_APPLY_TC_TO_SMP_SMP_7_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_SMP_6_LO = 6;
localparam CM_APPLY_TC_TO_SMP_SMP_6_HI = 6;
localparam CM_APPLY_TC_TO_SMP_SMP_6_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_SMP_5_LO = 5;
localparam CM_APPLY_TC_TO_SMP_SMP_5_HI = 5;
localparam CM_APPLY_TC_TO_SMP_SMP_5_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_SMP_4_LO = 4;
localparam CM_APPLY_TC_TO_SMP_SMP_4_HI = 4;
localparam CM_APPLY_TC_TO_SMP_SMP_4_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_SMP_3_LO = 3;
localparam CM_APPLY_TC_TO_SMP_SMP_3_HI = 3;
localparam CM_APPLY_TC_TO_SMP_SMP_3_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_SMP_2_LO = 2;
localparam CM_APPLY_TC_TO_SMP_SMP_2_HI = 2;
localparam CM_APPLY_TC_TO_SMP_SMP_2_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_SMP_1_LO = 1;
localparam CM_APPLY_TC_TO_SMP_SMP_1_HI = 1;
localparam CM_APPLY_TC_TO_SMP_SMP_1_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_SMP_0_LO = 0;
localparam CM_APPLY_TC_TO_SMP_SMP_0_HI = 0;
localparam CM_APPLY_TC_TO_SMP_SMP_0_RESET = 1'h0;
localparam CM_APPLY_TC_TO_SMP_USEMASK = 64'hFF;
localparam CM_APPLY_TC_TO_SMP_RO_MASK = 64'h0;
localparam CM_APPLY_TC_TO_SMP_WO_MASK = 64'h0;
localparam CM_APPLY_TC_TO_SMP_RESET = 64'h0;

typedef struct packed {
    logic [62:0] reserved0;  // RSVD
    logic  [0:0] CURRENT;  // RW
} CM_APPLY_MCAST_EPOCH_t;

localparam CM_APPLY_MCAST_EPOCH_REG_STRIDE = 48'h8;
localparam CM_APPLY_MCAST_EPOCH_REG_ENTRIES = 1;
localparam [47:0] CM_APPLY_MCAST_EPOCH_CR_ADDR = 48'h3708;
localparam CM_APPLY_MCAST_EPOCH_SIZE = 64;
localparam CM_APPLY_MCAST_EPOCH_CURRENT_LO = 0;
localparam CM_APPLY_MCAST_EPOCH_CURRENT_HI = 0;
localparam CM_APPLY_MCAST_EPOCH_CURRENT_RESET = 1'h0;
localparam CM_APPLY_MCAST_EPOCH_USEMASK = 64'h1;
localparam CM_APPLY_MCAST_EPOCH_RO_MASK = 64'h0;
localparam CM_APPLY_MCAST_EPOCH_WO_MASK = 64'h0;
localparam CM_APPLY_MCAST_EPOCH_RESET = 64'h0;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [0:0] RXS_7;  // RO/V
    logic  [0:0] RXS_6;  // RO/V
    logic  [0:0] RXS_5;  // RO/V
    logic  [0:0] RXS_4;  // RO/V
    logic  [0:0] RXS_3;  // RO/V
    logic  [0:0] RXS_2;  // RO/V
    logic  [0:0] RXS_1;  // RO/V
    logic  [0:0] RXS_0;  // RO/V
    logic  [0:0] GLOBAL_EX;  // RO/V
} CM_APPLY_STATE_t;

localparam CM_APPLY_STATE_REG_STRIDE = 48'h8;
localparam CM_APPLY_STATE_REG_ENTRIES = 1;
localparam [47:0] CM_APPLY_STATE_CR_ADDR = 48'h3710;
localparam CM_APPLY_STATE_SIZE = 64;
localparam CM_APPLY_STATE_RXS_7_LO = 8;
localparam CM_APPLY_STATE_RXS_7_HI = 8;
localparam CM_APPLY_STATE_RXS_7_RESET = 1'h0;
localparam CM_APPLY_STATE_RXS_6_LO = 7;
localparam CM_APPLY_STATE_RXS_6_HI = 7;
localparam CM_APPLY_STATE_RXS_6_RESET = 1'h0;
localparam CM_APPLY_STATE_RXS_5_LO = 6;
localparam CM_APPLY_STATE_RXS_5_HI = 6;
localparam CM_APPLY_STATE_RXS_5_RESET = 1'h0;
localparam CM_APPLY_STATE_RXS_4_LO = 5;
localparam CM_APPLY_STATE_RXS_4_HI = 5;
localparam CM_APPLY_STATE_RXS_4_RESET = 1'h0;
localparam CM_APPLY_STATE_RXS_3_LO = 4;
localparam CM_APPLY_STATE_RXS_3_HI = 4;
localparam CM_APPLY_STATE_RXS_3_RESET = 1'h0;
localparam CM_APPLY_STATE_RXS_2_LO = 3;
localparam CM_APPLY_STATE_RXS_2_HI = 3;
localparam CM_APPLY_STATE_RXS_2_RESET = 1'h0;
localparam CM_APPLY_STATE_RXS_1_LO = 2;
localparam CM_APPLY_STATE_RXS_1_HI = 2;
localparam CM_APPLY_STATE_RXS_1_RESET = 1'h0;
localparam CM_APPLY_STATE_RXS_0_LO = 1;
localparam CM_APPLY_STATE_RXS_0_HI = 1;
localparam CM_APPLY_STATE_RXS_0_RESET = 1'h0;
localparam CM_APPLY_STATE_GLOBAL_EX_LO = 0;
localparam CM_APPLY_STATE_GLOBAL_EX_HI = 0;
localparam CM_APPLY_STATE_GLOBAL_EX_RESET = 1'h0;
localparam CM_APPLY_STATE_USEMASK = 64'h1FF;
localparam CM_APPLY_STATE_RO_MASK = 64'h1FF;
localparam CM_APPLY_STATE_WO_MASK = 64'h0;
localparam CM_APPLY_STATE_RESET = 64'h0;

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic [23:0] DEST_MASK;  // RW
} CM_APPLY_CPU_TRAP_MASK_t;

localparam CM_APPLY_CPU_TRAP_MASK_REG_STRIDE = 48'h8;
localparam CM_APPLY_CPU_TRAP_MASK_REG_ENTRIES = 1;
localparam [47:0] CM_APPLY_CPU_TRAP_MASK_CR_ADDR = 48'h3718;
localparam CM_APPLY_CPU_TRAP_MASK_SIZE = 64;
localparam CM_APPLY_CPU_TRAP_MASK_DEST_MASK_LO = 0;
localparam CM_APPLY_CPU_TRAP_MASK_DEST_MASK_HI = 23;
localparam CM_APPLY_CPU_TRAP_MASK_DEST_MASK_RESET = 24'h1;
localparam CM_APPLY_CPU_TRAP_MASK_USEMASK = 64'hFFFFFF;
localparam CM_APPLY_CPU_TRAP_MASK_RO_MASK = 64'h0;
localparam CM_APPLY_CPU_TRAP_MASK_WO_MASK = 64'h0;
localparam CM_APPLY_CPU_TRAP_MASK_RESET = 64'h1;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic  [5:0] TRIGGER;  // RW
    logic  [5:0] TTL;  // RW
    logic  [5:0] ICMP;  // RW
    logic  [5:0] ARP_REDIRECT;  // RW
    logic  [5:0] RESERVED_MAC;  // RW
    logic  [5:0] FFU;  // RW
} CM_APPLY_LOG_MIRROR_PROFILE_t;

localparam CM_APPLY_LOG_MIRROR_PROFILE_REG_STRIDE = 48'h8;
localparam CM_APPLY_LOG_MIRROR_PROFILE_REG_ENTRIES = 1;
localparam [47:0] CM_APPLY_LOG_MIRROR_PROFILE_CR_ADDR = 48'h3720;
localparam CM_APPLY_LOG_MIRROR_PROFILE_SIZE = 64;
localparam CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER_LO = 30;
localparam CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER_HI = 35;
localparam CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER_RESET = 6'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_TTL_LO = 24;
localparam CM_APPLY_LOG_MIRROR_PROFILE_TTL_HI = 29;
localparam CM_APPLY_LOG_MIRROR_PROFILE_TTL_RESET = 6'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_ICMP_LO = 18;
localparam CM_APPLY_LOG_MIRROR_PROFILE_ICMP_HI = 23;
localparam CM_APPLY_LOG_MIRROR_PROFILE_ICMP_RESET = 6'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT_LO = 12;
localparam CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT_HI = 17;
localparam CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT_RESET = 6'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC_LO = 6;
localparam CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC_HI = 11;
localparam CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC_RESET = 6'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_FFU_LO = 0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_FFU_HI = 5;
localparam CM_APPLY_LOG_MIRROR_PROFILE_FFU_RESET = 6'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_USEMASK = 64'hFFFFFFFFF;
localparam CM_APPLY_LOG_MIRROR_PROFILE_RO_MASK = 64'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_WO_MASK = 64'h0;
localparam CM_APPLY_LOG_MIRROR_PROFILE_RESET = 64'h0;

typedef struct packed {
    logic [53:0] reserved0;  // RSVD
    logic  [0:0] QUEUE_DEPTH_MODE;  // RW
    logic  [2:0] QUEUE_DEPTH_START_BIT;  // RW
    logic  [0:0] SELECT_COMP;  // RW
    logic  [4:0] SAMPLE_RATE_EXP;  // RW
} CM_APPLY_QCN_CFG_t;

localparam CM_APPLY_QCN_CFG_REG_STRIDE = 48'h8;
localparam CM_APPLY_QCN_CFG_REG_ENTRIES = 1;
localparam CM_APPLY_QCN_CFG_CR_ADDR = 48'h3728;
localparam CM_APPLY_QCN_CFG_SIZE = 64;
localparam CM_APPLY_QCN_CFG_QUEUE_DEPTH_MODE_LO = 9;
localparam CM_APPLY_QCN_CFG_QUEUE_DEPTH_MODE_HI = 9;
localparam CM_APPLY_QCN_CFG_QUEUE_DEPTH_MODE_RESET = 1'h0;
localparam CM_APPLY_QCN_CFG_QUEUE_DEPTH_START_BIT_LO = 6;
localparam CM_APPLY_QCN_CFG_QUEUE_DEPTH_START_BIT_HI = 8;
localparam CM_APPLY_QCN_CFG_QUEUE_DEPTH_START_BIT_RESET = 3'h0;
localparam CM_APPLY_QCN_CFG_SELECT_COMP_LO = 5;
localparam CM_APPLY_QCN_CFG_SELECT_COMP_HI = 5;
localparam CM_APPLY_QCN_CFG_SELECT_COMP_RESET = 1'h0;
localparam CM_APPLY_QCN_CFG_SAMPLE_RATE_EXP_LO = 0;
localparam CM_APPLY_QCN_CFG_SAMPLE_RATE_EXP_HI = 4;
localparam CM_APPLY_QCN_CFG_SAMPLE_RATE_EXP_RESET = 5'h0;
localparam CM_APPLY_QCN_CFG_USEMASK = 64'h3FF;
localparam CM_APPLY_QCN_CFG_RO_MASK = 64'h0;
localparam CM_APPLY_QCN_CFG_WO_MASK = 64'h0;
localparam CM_APPLY_QCN_CFG_RESET = 64'h0;

typedef struct packed {
    CM_APPLY_TRAP_GLORT_t [15:0] CM_APPLY_TRAP_GLORT;
    CM_APPLY_TC_TO_SMP_t  CM_APPLY_TC_TO_SMP;
    CM_APPLY_MCAST_EPOCH_t  CM_APPLY_MCAST_EPOCH;
    CM_APPLY_STATE_t  CM_APPLY_STATE;
    CM_APPLY_CPU_TRAP_MASK_t  CM_APPLY_CPU_TRAP_MASK;
    CM_APPLY_LOG_MIRROR_PROFILE_t  CM_APPLY_LOG_MIRROR_PROFILE;
} mby_ppe_cm_apply_map_registers_t;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

typedef struct packed {
    logic  [0:0] RXS_7;  // RO/V
    logic  [0:0] RXS_6;  // RO/V
    logic  [0:0] RXS_5;  // RO/V
    logic  [0:0] RXS_4;  // RO/V
    logic  [0:0] RXS_3;  // RO/V
    logic  [0:0] RXS_2;  // RO/V
    logic  [0:0] RXS_1;  // RO/V
    logic  [0:0] RXS_0;  // RO/V
    logic  [0:0] GLOBAL_EX;  // RO/V
} new_CM_APPLY_STATE_t;

typedef struct packed {
    new_CM_APPLY_STATE_t  CM_APPLY_STATE;
} mby_ppe_cm_apply_map_new_t;

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_CM_APPLY_TX_SOFTDROP_CFG_t;

typedef logic [7:0] we_CM_APPLY_TX_TC_STATE_t;

typedef logic [7:0] we_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t;

typedef logic [7:0] we_CM_APPLY_RX_SMP_STATE_t;

typedef logic [7:0] we_CM_APPLY_MIRROR_PROFILE_TABLE_t;

typedef logic [7:0] we_CM_APPLY_DROP_COUNT_t;

typedef logic [7:0] we_CM_APPLY_LOOPBACK_SUPPRESS_t;

typedef logic [7:0] we_CM_APPLY_SOFTDROP_CFG_t;

typedef logic [7:0] we_CM_APPLY_SOFTDROP_STATE_t;

typedef logic [7:0] we_CM_APPLY_QCN_CFG_t;

typedef struct packed {
    we_CM_APPLY_TX_SOFTDROP_CFG_t CM_APPLY_TX_SOFTDROP_CFG;
    we_CM_APPLY_TX_TC_STATE_t CM_APPLY_TX_TC_STATE;
    we_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
    we_CM_APPLY_RX_SMP_STATE_t CM_APPLY_RX_SMP_STATE;
    we_CM_APPLY_MIRROR_PROFILE_TABLE_t CM_APPLY_MIRROR_PROFILE_TABLE;
    we_CM_APPLY_DROP_COUNT_t CM_APPLY_DROP_COUNT;
    we_CM_APPLY_LOOPBACK_SUPPRESS_t CM_APPLY_LOOPBACK_SUPPRESS;
    we_CM_APPLY_SOFTDROP_CFG_t CM_APPLY_SOFTDROP_CFG;
    we_CM_APPLY_SOFTDROP_STATE_t CM_APPLY_SOFTDROP_STATE;
    we_CM_APPLY_QCN_CFG_t CM_APPLY_QCN_CFG;
} mby_ppe_cm_apply_map_handcoded_t;

typedef logic [7:0] re_CM_APPLY_TX_SOFTDROP_CFG_t;

typedef logic [7:0] re_CM_APPLY_TX_TC_STATE_t;

typedef logic [7:0] re_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t;

typedef logic [7:0] re_CM_APPLY_RX_SMP_STATE_t;

typedef logic [7:0] re_CM_APPLY_MIRROR_PROFILE_TABLE_t;

typedef logic [7:0] re_CM_APPLY_DROP_COUNT_t;

typedef logic [7:0] re_CM_APPLY_LOOPBACK_SUPPRESS_t;

typedef logic [7:0] re_CM_APPLY_SOFTDROP_CFG_t;

typedef logic [7:0] re_CM_APPLY_SOFTDROP_STATE_t;

typedef logic [7:0] re_CM_APPLY_QCN_CFG_t;

typedef struct packed {
    re_CM_APPLY_TX_SOFTDROP_CFG_t CM_APPLY_TX_SOFTDROP_CFG;
    re_CM_APPLY_TX_TC_STATE_t CM_APPLY_TX_TC_STATE;
    re_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
    re_CM_APPLY_RX_SMP_STATE_t CM_APPLY_RX_SMP_STATE;
    re_CM_APPLY_MIRROR_PROFILE_TABLE_t CM_APPLY_MIRROR_PROFILE_TABLE;
    re_CM_APPLY_DROP_COUNT_t CM_APPLY_DROP_COUNT;
    re_CM_APPLY_LOOPBACK_SUPPRESS_t CM_APPLY_LOOPBACK_SUPPRESS;
    re_CM_APPLY_SOFTDROP_CFG_t CM_APPLY_SOFTDROP_CFG;
    re_CM_APPLY_SOFTDROP_STATE_t CM_APPLY_SOFTDROP_STATE;
    re_CM_APPLY_QCN_CFG_t CM_APPLY_QCN_CFG;
} mby_ppe_cm_apply_map_hc_re_t;

typedef logic handcode_rvalid_CM_APPLY_TX_SOFTDROP_CFG_t;

typedef logic handcode_rvalid_CM_APPLY_TX_TC_STATE_t;

typedef logic handcode_rvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t;

typedef logic handcode_rvalid_CM_APPLY_RX_SMP_STATE_t;

typedef logic handcode_rvalid_CM_APPLY_MIRROR_PROFILE_TABLE_t;

typedef logic handcode_rvalid_CM_APPLY_DROP_COUNT_t;

typedef logic handcode_rvalid_CM_APPLY_LOOPBACK_SUPPRESS_t;

typedef logic handcode_rvalid_CM_APPLY_SOFTDROP_CFG_t;

typedef logic handcode_rvalid_CM_APPLY_SOFTDROP_STATE_t;

typedef logic handcode_rvalid_CM_APPLY_QCN_CFG_t;

typedef struct packed {
    handcode_rvalid_CM_APPLY_TX_SOFTDROP_CFG_t CM_APPLY_TX_SOFTDROP_CFG;
    handcode_rvalid_CM_APPLY_TX_TC_STATE_t CM_APPLY_TX_TC_STATE;
    handcode_rvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
    handcode_rvalid_CM_APPLY_RX_SMP_STATE_t CM_APPLY_RX_SMP_STATE;
    handcode_rvalid_CM_APPLY_MIRROR_PROFILE_TABLE_t CM_APPLY_MIRROR_PROFILE_TABLE;
    handcode_rvalid_CM_APPLY_DROP_COUNT_t CM_APPLY_DROP_COUNT;
    handcode_rvalid_CM_APPLY_LOOPBACK_SUPPRESS_t CM_APPLY_LOOPBACK_SUPPRESS;
    handcode_rvalid_CM_APPLY_SOFTDROP_CFG_t CM_APPLY_SOFTDROP_CFG;
    handcode_rvalid_CM_APPLY_SOFTDROP_STATE_t CM_APPLY_SOFTDROP_STATE;
    handcode_rvalid_CM_APPLY_QCN_CFG_t CM_APPLY_QCN_CFG;
} mby_ppe_cm_apply_map_hc_rvalid_t;

typedef logic handcode_wvalid_CM_APPLY_TX_SOFTDROP_CFG_t;

typedef logic handcode_wvalid_CM_APPLY_TX_TC_STATE_t;

typedef logic handcode_wvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t;

typedef logic handcode_wvalid_CM_APPLY_RX_SMP_STATE_t;

typedef logic handcode_wvalid_CM_APPLY_MIRROR_PROFILE_TABLE_t;

typedef logic handcode_wvalid_CM_APPLY_DROP_COUNT_t;

typedef logic handcode_wvalid_CM_APPLY_LOOPBACK_SUPPRESS_t;

typedef logic handcode_wvalid_CM_APPLY_SOFTDROP_CFG_t;

typedef logic handcode_wvalid_CM_APPLY_SOFTDROP_STATE_t;

typedef logic handcode_wvalid_CM_APPLY_QCN_CFG_t;

typedef struct packed {
    handcode_wvalid_CM_APPLY_TX_SOFTDROP_CFG_t CM_APPLY_TX_SOFTDROP_CFG;
    handcode_wvalid_CM_APPLY_TX_TC_STATE_t CM_APPLY_TX_TC_STATE;
    handcode_wvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
    handcode_wvalid_CM_APPLY_RX_SMP_STATE_t CM_APPLY_RX_SMP_STATE;
    handcode_wvalid_CM_APPLY_MIRROR_PROFILE_TABLE_t CM_APPLY_MIRROR_PROFILE_TABLE;
    handcode_wvalid_CM_APPLY_DROP_COUNT_t CM_APPLY_DROP_COUNT;
    handcode_wvalid_CM_APPLY_LOOPBACK_SUPPRESS_t CM_APPLY_LOOPBACK_SUPPRESS;
    handcode_wvalid_CM_APPLY_SOFTDROP_CFG_t CM_APPLY_SOFTDROP_CFG;
    handcode_wvalid_CM_APPLY_SOFTDROP_STATE_t CM_APPLY_SOFTDROP_STATE;
    handcode_wvalid_CM_APPLY_QCN_CFG_t CM_APPLY_QCN_CFG;
} mby_ppe_cm_apply_map_hc_wvalid_t;

typedef logic handcode_error_CM_APPLY_TX_SOFTDROP_CFG_t;

typedef logic handcode_error_CM_APPLY_TX_TC_STATE_t;

typedef logic handcode_error_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t;

typedef logic handcode_error_CM_APPLY_RX_SMP_STATE_t;

typedef logic handcode_error_CM_APPLY_MIRROR_PROFILE_TABLE_t;

typedef logic handcode_error_CM_APPLY_DROP_COUNT_t;

typedef logic handcode_error_CM_APPLY_LOOPBACK_SUPPRESS_t;

typedef logic handcode_error_CM_APPLY_SOFTDROP_CFG_t;

typedef logic handcode_error_CM_APPLY_SOFTDROP_STATE_t;

typedef logic handcode_error_CM_APPLY_QCN_CFG_t;

typedef struct packed {
    handcode_error_CM_APPLY_TX_SOFTDROP_CFG_t CM_APPLY_TX_SOFTDROP_CFG;
    handcode_error_CM_APPLY_TX_TC_STATE_t CM_APPLY_TX_TC_STATE;
    handcode_error_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
    handcode_error_CM_APPLY_RX_SMP_STATE_t CM_APPLY_RX_SMP_STATE;
    handcode_error_CM_APPLY_MIRROR_PROFILE_TABLE_t CM_APPLY_MIRROR_PROFILE_TABLE;
    handcode_error_CM_APPLY_DROP_COUNT_t CM_APPLY_DROP_COUNT;
    handcode_error_CM_APPLY_LOOPBACK_SUPPRESS_t CM_APPLY_LOOPBACK_SUPPRESS;
    handcode_error_CM_APPLY_SOFTDROP_CFG_t CM_APPLY_SOFTDROP_CFG;
    handcode_error_CM_APPLY_SOFTDROP_STATE_t CM_APPLY_SOFTDROP_STATE;
    handcode_error_CM_APPLY_QCN_CFG_t CM_APPLY_QCN_CFG;
} mby_ppe_cm_apply_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    CM_APPLY_TX_SOFTDROP_CFG_t CM_APPLY_TX_SOFTDROP_CFG;
    CM_APPLY_TX_TC_STATE_t CM_APPLY_TX_TC_STATE;
    CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
    CM_APPLY_RX_SMP_STATE_t CM_APPLY_RX_SMP_STATE;
    CM_APPLY_MIRROR_PROFILE_TABLE_t CM_APPLY_MIRROR_PROFILE_TABLE;
    CM_APPLY_DROP_COUNT_t CM_APPLY_DROP_COUNT;
    CM_APPLY_LOOPBACK_SUPPRESS_t CM_APPLY_LOOPBACK_SUPPRESS;
    CM_APPLY_SOFTDROP_CFG_t CM_APPLY_SOFTDROP_CFG;
    CM_APPLY_SOFTDROP_STATE_t CM_APPLY_SOFTDROP_STATE;
    CM_APPLY_QCN_CFG_t CM_APPLY_QCN_CFG;
} mby_ppe_cm_apply_map_hc_reg_read_t;

typedef struct packed {
    CM_APPLY_TX_SOFTDROP_CFG_t CM_APPLY_TX_SOFTDROP_CFG;
    CM_APPLY_TX_TC_STATE_t CM_APPLY_TX_TC_STATE;
    CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
    CM_APPLY_RX_SMP_STATE_t CM_APPLY_RX_SMP_STATE;
    CM_APPLY_MIRROR_PROFILE_TABLE_t CM_APPLY_MIRROR_PROFILE_TABLE;
    CM_APPLY_DROP_COUNT_t CM_APPLY_DROP_COUNT;
    CM_APPLY_LOOPBACK_SUPPRESS_t CM_APPLY_LOOPBACK_SUPPRESS;
    CM_APPLY_SOFTDROP_CFG_t CM_APPLY_SOFTDROP_CFG;
    CM_APPLY_SOFTDROP_STATE_t CM_APPLY_SOFTDROP_STATE;
    CM_APPLY_QCN_CFG_t CM_APPLY_QCN_CFG;
} mby_ppe_cm_apply_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_cm_apply_map_pkg

`endif // MBY_PPE_CM_APPLY_MAP_PKG_VH
