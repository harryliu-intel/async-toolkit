magic
tech scmos
timestamp 962800458
<< ndiffusion >>
rect 54 24 62 25
rect 54 16 62 21
rect 84 16 92 17
rect 54 8 62 13
rect 84 8 92 13
rect 54 4 62 5
rect 54 -5 62 -4
rect 54 -13 62 -8
rect 84 4 92 5
rect 84 -5 92 -4
rect 175 0 183 1
rect 84 -13 92 -8
rect 175 -4 183 -3
rect 175 -13 183 -12
rect 54 -21 62 -16
rect 84 -17 92 -16
rect 54 -25 62 -24
rect 175 -17 183 -16
<< pdiffusion >>
rect 131 30 141 35
rect 131 29 149 30
rect 131 25 149 26
rect 131 20 137 25
rect 108 16 116 17
rect 137 16 149 17
rect 108 8 116 13
rect 108 4 116 5
rect 108 -5 116 -4
rect 137 8 149 13
rect 137 4 149 5
rect 137 -5 149 -4
rect 199 0 207 1
rect 108 -13 116 -8
rect 137 -13 149 -8
rect 199 -4 207 -3
rect 199 -13 207 -12
rect 108 -17 116 -16
rect 137 -17 149 -16
rect 199 -17 207 -16
<< ntransistor >>
rect 54 21 62 24
rect 54 13 62 16
rect 84 13 92 16
rect 54 5 62 8
rect 84 5 92 8
rect 54 -8 62 -5
rect 84 -8 92 -5
rect 175 -3 183 0
rect 54 -16 62 -13
rect 84 -16 92 -13
rect 175 -16 183 -13
rect 54 -24 62 -21
<< ptransistor >>
rect 131 26 149 29
rect 108 13 116 16
rect 137 13 149 16
rect 108 5 116 8
rect 137 5 149 8
rect 108 -8 116 -5
rect 137 -8 149 -5
rect 199 -3 207 0
rect 108 -16 116 -13
rect 137 -16 149 -13
rect 199 -16 207 -13
<< polysilicon >>
rect 127 26 131 29
rect 149 26 153 29
rect 50 21 54 24
rect 62 21 67 24
rect 50 13 54 16
rect 62 13 84 16
rect 92 13 108 16
rect 116 13 137 16
rect 149 13 153 16
rect 49 5 54 8
rect 62 5 67 8
rect 72 5 84 8
rect 92 5 108 8
rect 116 5 120 8
rect 49 0 52 5
rect 50 -5 52 0
rect 50 -8 54 -5
rect 62 -8 67 -5
rect 72 -13 75 5
rect 125 -5 128 13
rect 133 5 137 8
rect 149 5 154 8
rect 151 0 154 5
rect 151 -5 153 0
rect 80 -8 84 -5
rect 92 -8 108 -5
rect 116 -8 128 -5
rect 133 -8 137 -5
rect 149 -8 153 -5
rect 170 -3 175 0
rect 183 -3 199 0
rect 207 -3 212 0
rect 170 -13 173 -3
rect 209 -13 212 -3
rect 50 -16 54 -13
rect 62 -16 84 -13
rect 92 -16 108 -13
rect 116 -16 137 -13
rect 149 -16 153 -13
rect 170 -16 175 -13
rect 183 -16 199 -13
rect 207 -16 212 -13
rect 50 -24 54 -21
rect 62 -24 66 -21
<< ndcontact >>
rect 54 25 62 33
rect 84 17 92 25
rect 54 -4 62 4
rect 84 -4 92 4
rect 175 1 183 9
rect 175 -12 183 -4
rect 84 -25 92 -17
rect 175 -25 183 -17
rect 54 -33 62 -25
<< pdcontact >>
rect 141 30 149 38
rect 108 17 116 25
rect 137 17 149 25
rect 108 -4 116 4
rect 137 -4 149 4
rect 199 1 207 9
rect 199 -12 207 -4
rect 108 -25 116 -17
rect 137 -25 149 -17
rect 199 -25 207 -17
<< polycontact >>
rect 42 -8 50 0
rect 153 -8 161 0
<< metal1 >>
rect 141 34 149 38
rect 54 25 62 33
rect 141 30 157 34
rect 54 17 92 25
rect 108 17 149 25
rect 153 8 157 30
rect 145 4 157 8
rect 42 -8 50 0
rect 54 -4 149 4
rect 175 1 183 9
rect 199 1 207 9
rect 153 -8 161 0
rect 45 -13 158 -8
rect 175 -12 207 -4
rect 54 -25 92 -17
rect 108 -25 149 -17
rect 175 -25 183 -17
rect 199 -25 207 -17
rect 54 -33 62 -25
<< labels >>
rlabel metal1 112 21 112 21 5 Vdd!
rlabel metal1 112 -21 112 -21 1 Vdd!
rlabel polysilicon 53 14 53 14 3 b
rlabel polysilicon 53 -15 53 -15 3 a
rlabel polysilicon 150 -14 150 -14 7 a
rlabel polysilicon 150 15 150 15 7 b
rlabel metal1 143 21 143 21 5 Vdd!
rlabel metal1 143 -21 143 -21 1 Vdd!
rlabel polysilicon 53 22 53 22 1 _SReset!
rlabel metal1 58 -29 58 -29 1 GND!
rlabel polysilicon 53 -23 53 -23 1 _SReset!
rlabel metal1 157 -4 157 -4 1 x
rlabel metal1 46 -4 46 -4 1 x
rlabel metal1 58 0 58 0 1 _x
rlabel metal1 88 0 88 0 1 _x
rlabel metal1 112 0 112 0 1 _x
rlabel metal1 143 0 143 0 1 _x
rlabel metal1 88 -21 88 -21 1 GND!
rlabel metal1 88 21 88 21 5 GND!
rlabel metal1 58 29 58 29 5 GND!
rlabel ndcontact 179 -8 179 -8 1 x
rlabel pdcontact 203 -8 203 -8 1 x
rlabel pdcontact 203 -21 203 -21 1 Vdd!
rlabel pdcontact 203 5 203 5 5 Vdd!
rlabel ndcontact 179 5 179 5 5 GND!
rlabel polysilicon 174 -2 174 -2 1 _x
rlabel polysilicon 174 -15 174 -15 1 _x
rlabel polysilicon 208 -2 208 -2 1 _x
rlabel polysilicon 208 -15 208 -15 1 _x
rlabel space 169 -26 176 10 7 ^n2
rlabel space 206 -26 213 10 3 ^p2
rlabel ndcontact 179 -21 179 -21 1 GND!
rlabel polysilicon 150 28 150 28 7 _PReset!
rlabel metal1 145 34 145 34 5 _x
rlabel space 41 -34 85 34 7 ^n1
rlabel space 115 -26 162 40 3 ^p1
<< end >>
