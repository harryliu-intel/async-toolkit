module mby_checker(

                   );

`include "mby_sva_include.sv"

endmodule 
