// vim: noai : ts=3 : sw=3 : expandtab : ft=systemverilog

//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors.  The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//=======================================================================
// COPYRIGHT (C)  2012 SYNOPSYS INC.
// This software and the associated documentation are confidential and
// proprietary to Synopsys, Inc. Your use or disclosure of this software
// is subject to the terms and conditions of a written license agreement
// between you, or your company, and Synopsys, Inc. In the event of
// publications, the following notice is applicable:
//
// ALL RIGHTS RESERVED
//
// The entire notice above must be reproduced on all authorized copies.
//
//------------------------------------------------------------------------------
//   Author        : Akshay Kotian
//   Project       : Madison Bay
//------------------------------------------------------------------------------

//Class:    axi_master_directed_sequence
//
// This directed sequence demonstrates the way user can control AXI BFM to
//generate AXI Master transactions.
//This class defines a sequence in which a AXI WRITE followed by a AXI READ
//sequence is generated by assigning values to the transactions rather than
//randomization, and then transmitted using `uvm_send.
//
//Execution phase: main_phase
//Sequencer: Master agent sequencer
//

`ifndef __AXI_MASTER_DIRECTED_SEQUENCE_GUARD
`define __AXI_MASTER_DIRECTED_SEQUENCE_GUARD


`ifndef __INSIDE_SVT_AXI_BFM_PKG__
`error "File is meant to be used only through the svt_axi_bfm_pkg.  Do not include it individually."
`endif

class axi_master_directed_sequence extends svt_axi_master_base_sequence;

    // Parameter that controls the number of transactions that will be generated
    rand int unsigned sequence_length = 10;

    //Constrain the sequence length to a reasonable value
    constraint reasonable_sequence_length {
        sequence_length <= 100;
    }

    //UVM Object Utility macro
    `uvm_object_utils(axi_master_directed_sequence)

    // Class Constructor
    function new(string name="axi_master_directed_sequence");
        super.new(name);
    endfunction

    virtual task body();
        svt_axi_master_transaction write_tran, read_tran;
        bit status;
        `uvm_info("body", "Started running axi_master_directed_sequence..", UVM_LOW)

        super.body();

        status = uvm_config_db #(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
        `uvm_info("body", $sformatf("sequence_length is %0d as a result of %0s.", sequence_length, status ? "config DB" : "randomization"), UVM_LOW);

        // Obtain a handle to the port configuration
        get_port_cfg();

        for(int i = 0; i < sequence_length; i++) begin

            // Set up the write transaction
            `uvm_create(write_tran)
            write_tran.port_cfg     = cfg;
            write_tran.xact_type    = svt_axi_transaction::WRITE;
            write_tran.addr         = 32'h0400_0000 | ('h400 * i);
            write_tran.burst_type   = svt_axi_transaction::INCR;
            write_tran.burst_size   = svt_axi_transaction::BURST_SIZE_32BIT;
            write_tran.atomic_type  = svt_axi_transaction::NORMAL;
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
            write_tran.burst_length = 1;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
            write_tran.burst_length = 2;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
            write_tran.burst_length = 4;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_4
            write_tran.burst_length = 8;
`else
            write_tran.burst_length = 16;
`endif
            write_tran.data         = new[write_tran.burst_length];
            write_tran.wstrb        = new[write_tran.burst_length];
            write_tran.data_user    = new[write_tran.burst_length];
            foreach (write_tran.data[i]) begin
                write_tran.data[i] = i;
            end
            foreach(write_tran.wstrb[i]) begin
                write_tran.wstrb[i] = 4'hf;
            end
            write_tran.wvalid_delay = new[write_tran.burst_length];
            foreach (write_tran.wvalid_delay[i]) begin
                write_tran.wvalid_delay[i]=i;
            end

            // Send the write transaction
            `uvm_send(write_tran)

            // Wait for the write transaction to complete
            get_response(rsp);

            `uvm_info("body", "AXI WRITE transaction completed", UVM_LOW);

            // Set up the read transaction
            `uvm_create(read_tran)
            read_tran.port_cfg     = cfg;
            read_tran.xact_type    = svt_axi_transaction::READ;
            read_tran.addr         = 32'h0400_0000 | ('h400 * i);
            read_tran.burst_type   = svt_axi_transaction::INCR;
            read_tran.burst_size   = svt_axi_transaction::BURST_SIZE_32BIT;
            read_tran.atomic_type  = svt_axi_transaction::NORMAL;
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
            read_tran.burst_length = 1;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
            read_tran.burst_length = 2;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
            read_tran.burst_length = 4;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_4
            read_tran.burst_length = 8;
`else
            read_tran.burst_length = 16;
`endif
            read_tran.rresp        = new[read_tran.burst_length];
            read_tran.data         = new[read_tran.burst_length];
            read_tran.rready_delay = new[read_tran.burst_length];
            read_tran.data_user    = new[read_tran.burst_length];
            foreach (read_tran.rready_delay[i]) begin
                read_tran.rready_delay[i]=i;
            end

            // Send the read transaction
            `uvm_send(read_tran)

            // Wait for the read transaction to complete
            get_response(rsp);

            `uvm_info("body", "AXI READ transaction completed", UVM_LOW);
        end

        `uvm_info("body", "Exiting...", UVM_LOW)
    endtask: body

    task get_port_cfg();
        svt_configuration get_cfg;

        // Obtain a handle to the port configuration
        p_sequencer.get_cfg(get_cfg);
        if (!$cast(cfg, get_cfg)) begin
            `uvm_fatal("body", "Unable to $cast the configuration to a svt_axi_port_configuration class");
        end

    endtask

endclass: axi_master_directed_sequence

`endif // __AXI_MASTER_DIRECTED_SEQUENCE_GUARD


