magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 192 638 198 639
rect 192 632 198 636
rect 192 629 198 630
rect 192 625 194 629
rect 192 624 198 625
rect 192 618 198 622
rect 192 615 198 616
rect 192 610 198 611
rect 192 604 198 608
rect 192 601 198 602
rect 192 597 194 601
rect 192 596 198 597
rect 192 590 198 594
rect 192 587 198 588
<< pdiffusion >>
rect 210 642 220 643
rect 210 639 220 640
rect 218 635 220 639
rect 210 634 220 635
rect 210 631 220 632
rect 210 627 216 631
rect 210 626 220 627
rect 210 623 220 624
rect 218 619 220 623
rect 210 618 220 619
rect 210 615 220 616
rect 210 611 216 615
rect 210 610 220 611
rect 210 607 220 608
rect 218 603 220 607
rect 210 602 220 603
rect 210 599 220 600
rect 210 595 216 599
rect 210 594 220 595
rect 210 591 220 592
rect 218 587 220 591
rect 210 586 220 587
rect 210 583 220 584
<< ntransistor >>
rect 192 636 198 638
rect 192 630 198 632
rect 192 622 198 624
rect 192 616 198 618
rect 192 608 198 610
rect 192 602 198 604
rect 192 594 198 596
rect 192 588 198 590
<< ptransistor >>
rect 210 640 220 642
rect 210 632 220 634
rect 210 624 220 626
rect 210 616 220 618
rect 210 608 220 610
rect 210 600 220 602
rect 210 592 220 594
rect 210 584 220 586
<< polysilicon >>
rect 200 640 210 642
rect 220 640 223 642
rect 200 638 202 640
rect 189 636 192 638
rect 198 636 202 638
rect 206 632 210 634
rect 220 632 223 634
rect 189 630 192 632
rect 198 630 208 632
rect 206 624 210 626
rect 220 624 223 626
rect 189 622 192 624
rect 198 622 208 624
rect 189 616 192 618
rect 198 616 210 618
rect 220 616 223 618
rect 189 608 192 610
rect 198 608 210 610
rect 220 608 223 610
rect 189 602 192 604
rect 198 602 208 604
rect 206 600 210 602
rect 220 600 223 602
rect 189 594 192 596
rect 198 594 208 596
rect 206 592 210 594
rect 220 592 223 594
rect 189 588 192 590
rect 198 588 202 590
rect 200 586 202 588
rect 200 584 210 586
rect 220 584 223 586
<< ndcontact >>
rect 192 639 198 643
rect 194 625 198 629
rect 192 611 198 615
rect 194 597 198 601
rect 192 583 198 587
<< pdcontact >>
rect 210 643 220 647
rect 210 635 218 639
rect 216 627 220 631
rect 210 619 218 623
rect 216 611 220 615
rect 210 603 218 607
rect 216 595 220 599
rect 210 587 218 591
rect 210 579 220 583
<< metal1 >>
rect 210 643 220 647
rect 192 639 198 643
rect 210 635 218 639
rect 210 629 213 635
rect 194 625 213 629
rect 216 627 220 631
rect 210 623 213 625
rect 210 619 218 623
rect 192 611 198 615
rect 210 607 213 619
rect 216 611 220 615
rect 210 603 218 607
rect 210 601 213 603
rect 194 597 213 601
rect 210 591 213 597
rect 216 595 220 599
rect 210 587 218 591
rect 192 583 198 587
rect 210 579 220 583
<< labels >>
rlabel space 189 582 195 644 7 ^n
rlabel polysilicon 191 603 191 603 3 a
rlabel polysilicon 191 609 191 609 3 b
rlabel polysilicon 191 589 191 589 3 a
rlabel polysilicon 191 595 191 595 3 b
rlabel polysilicon 191 623 191 623 3 b
rlabel polysilicon 191 617 191 617 3 a
rlabel polysilicon 191 637 191 637 3 b
rlabel polysilicon 191 631 191 631 3 a
rlabel space 217 578 224 648 3 ^p
rlabel polysilicon 221 641 221 641 3 b
rlabel polysilicon 221 625 221 625 3 b
rlabel polysilicon 221 609 221 609 3 b
rlabel polysilicon 221 593 221 593 3 b
rlabel polysilicon 221 585 221 585 3 a
rlabel polysilicon 221 601 221 601 3 a
rlabel polysilicon 221 617 221 617 3 a
rlabel polysilicon 221 633 221 633 3 a
rlabel ndcontact 196 641 196 641 1 GND!
rlabel ndcontact 196 627 196 627 1 x
rlabel ndcontact 196 613 196 613 1 GND!
rlabel ndcontact 196 599 196 599 1 x
rlabel ndcontact 196 585 196 585 1 GND!
rlabel pdcontact 212 589 212 589 1 x
rlabel pdcontact 212 605 212 605 1 x
rlabel pdcontact 212 621 212 621 1 x
rlabel pdcontact 212 637 212 637 1 x
rlabel pdcontact 218 629 218 629 1 Vdd!
rlabel pdcontact 218 613 218 613 1 Vdd!
rlabel pdcontact 218 597 218 597 1 Vdd!
rlabel pdcontact 218 581 218 581 1 Vdd!
rlabel pdcontact 218 645 218 645 1 Vdd!
<< end >>
