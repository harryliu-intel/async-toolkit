magic
tech scmos
timestamp 988943070
<< nselect >>
rect -34 8 0 63
<< pselect >>
rect 0 -1 46 66
<< ndiffusion >>
rect -28 49 -8 50
rect -28 41 -8 46
rect -28 33 -8 38
rect -28 25 -8 30
rect -28 21 -8 22
<< pdiffusion >>
rect 8 54 40 55
rect 8 50 40 51
rect 28 42 40 50
rect 8 41 40 42
rect 8 37 40 38
rect 8 28 40 29
rect 8 24 40 25
rect 8 13 24 16
rect 8 9 24 10
<< ntransistor >>
rect -28 46 -8 49
rect -28 38 -8 41
rect -28 30 -8 33
rect -28 22 -8 25
<< ptransistor >>
rect 8 51 40 54
rect 8 38 40 41
rect 8 25 40 28
rect 8 10 24 13
<< polysilicon >>
rect 3 51 8 54
rect 40 51 44 54
rect 3 49 6 51
rect -32 46 -28 49
rect -8 46 6 49
rect -32 38 -28 41
rect -8 38 8 41
rect 40 38 44 41
rect -32 30 -28 33
rect -8 30 6 33
rect 3 28 6 30
rect 3 25 8 28
rect 40 25 44 28
rect -32 22 -28 25
rect -8 22 -4 25
rect 4 10 8 13
rect 24 10 28 13
<< ndcontact >>
rect -28 50 -8 58
rect -28 13 -8 21
<< pdcontact >>
rect 8 55 40 63
rect 8 42 28 50
rect 8 29 40 37
rect 8 16 40 24
rect 8 1 24 9
<< metal1 >>
rect -28 50 -8 58
rect 8 55 40 63
rect -16 42 28 50
rect -4 24 4 42
rect 32 37 40 55
rect 8 29 40 37
rect -28 13 -8 21
rect -4 16 40 24
rect 8 1 24 9
<< labels >>
rlabel space -35 -1 -28 66 7 ^n
rlabel space 28 20 47 66 3 ^p
rlabel metal1 -28 13 -8 21 1 GND!|pin|s|0
rlabel metal1 32 29 40 63 1 Vdd!|pin|s|1
rlabel metal1 -4 16 4 50 1 x|pin|s|2
rlabel metal1 -28 50 -8 58 1 x|pin|s|2
rlabel metal1 -16 42 28 50 1 x|pin|s|2
rlabel metal1 -4 16 40 24 1 x|pin|s|2
rlabel polysilicon 40 25 44 28 1 a|pin|w|3|poly
rlabel polysilicon 3 25 7 28 1 a|pin|w|3|poly
rlabel polysilicon -32 30 -28 33 1 a|pin|w|3|poly
rlabel polysilicon -32 38 -28 41 1 b|pin|w|4|poly
rlabel polysilicon 40 38 44 41 1 b|pin|w|4|poly
rlabel polysilicon 40 51 44 54 1 c|pin|w|5|poly
rlabel polysilicon 3 51 7 54 1 c|pin|w|5|poly
rlabel polysilicon -32 46 -28 49 1 c|pin|w|5|poly
rlabel polysilicon -32 22 -28 25 1 _SReset!|pin|w|6|poly
rlabel polysilicon -8 22 -4 25 1 _SReset!|pin|w|6|poly
rlabel polysilicon 4 10 8 13 1 _PReset!|pin|w|7|poly
rlabel polysilicon 24 10 28 13 1 _PReset!|pin|w|7|poly
rlabel metal1 8 55 40 63 1 Vdd!|pin|s|1
rlabel metal1 8 29 40 37 1 Vdd!|pin|s|1
rlabel metal1 8 1 24 9 1 Vdd!|pin|s|0
<< end >>
