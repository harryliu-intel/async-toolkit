// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Mike Jarvis <michael.a.jarvis.com> 
// -- Project Name : MBY 
// -- Description  : mpp (MegaPort Pair) netlist. 
// ------------------------------------------------------------------- 

module TB_MGP

(
  
);
//Input List
logic                   arst_n;                                   //Asynchronous negedge reset     
logic                   cclk;                                     
logic            [7:0]  grp_a0_rx_data_valid;                     
logic            [1:0]  grp_a0_rx_port_num;                       
logic            [7:0]  grp_a1_rx_data_valid;                     
logic            [1:0]  grp_a1_rx_port_num;                       
logic            [7:0]  grp_b0_rx_data_valid;                     
logic            [1:0]  grp_b0_rx_port_num;                       
logic            [7:0]  grp_b1_rx_data_valid;                     
logic            [1:0]  grp_b1_rx_port_num;                       
logic            [7:0]  grp_c0_rx_data_valid;                     
logic            [1:0]  grp_c0_rx_port_num;                       
logic            [7:0]  grp_c1_rx_data_valid;                     
logic            [1:0]  grp_c1_rx_port_num;                       
logic            [7:0]  grp_d0_rx_data_valid;                     
logic            [1:0]  grp_d0_rx_port_num;                       
logic            [7:0]  grp_d1_rx_data_valid;                     
logic            [1:0]  grp_d1_rx_port_num;                       
logic           [19:0]  igr0_vp_cpp_rx_metadata;                  
logic            [7:0]  igr0_vp_rx_data_valid;                    
logic            [7:0]  igr0_vp_rx_ecc;                           
logic            [2:0]  igr0_vp_rx_flow_control_tc;               
logic           [23:0]  igr0_vp_rx_metadata;                      
logic            [1:0]  igr0_vp_rx_port_num;                      
logic           [35:0]  igr0_vp_rx_time_stamp;                    
logic           [19:0]  igr1_vp_cpp_rx_metadata;                  
logic            [7:0]  igr1_vp_rx_data_valid;                    
logic            [7:0]  igr1_vp_rx_ecc;                           
logic            [2:0]  igr1_vp_rx_flow_control_tc;               
logic           [23:0]  igr1_vp_rx_metadata;                      
logic            [1:0]  igr1_vp_rx_port_num;                      
logic           [35:0]  igr1_vp_rx_time_stamp;                    
//edr logic           [31:0]  i_mpp_csr_end;                            // tied in mpp shell 
//edr logic           [31:0]  i_mpp_csr_start;                          // tied in mpp shell  
logic           [23:0]  mpp_dqring_in_0_0;                        
logic           [23:0]  mpp_dqring_in_0_1;                        
logic           [23:0]  mpp_dqring_in_1_0;                        
logic           [23:0]  mpp_dqring_in_1_1;                        
logic           [23:0]  mpp_dqring_in_2_0;                        
logic           [23:0]  mpp_dqring_in_2_1;                        
logic           [23:0]  mpp_dqring_in_3_0;                        
logic           [23:0]  mpp_dqring_in_3_1;                        
logic           [23:0]  mpp_dqring_in_4_0;                        
logic           [23:0]  mpp_dqring_in_4_1;                        
logic           [23:0]  mpp_dqring_in_5_0;                        
logic           [23:0]  mpp_dqring_in_5_1;                        
logic           [23:0]  mpp_dqring_in_6_0;                        
logic           [23:0]  mpp_dqring_in_6_1;                        
logic           [23:0]  mpp_dqring_in_7_0;                        
logic           [23:0]  mpp_dqring_in_7_1;                        
logic           [25:0]  mpp_gpolring_in_0_0;                      
logic           [25:0]  mpp_gpolring_in_0_1;                      
logic           [25:0]  mpp_gpolring_in_1_0;                      
logic           [25:0]  mpp_gpolring_in_1_1;                      
logic           [25:0]  mpp_gpolring_in_2_0;                      
logic           [25:0]  mpp_gpolring_in_2_1;                      
logic           [25:0]  mpp_gpolring_in_3_0;                      
logic           [25:0]  mpp_gpolring_in_3_1;                      
logic           [25:0]  mpp_gpolring_in_4_0;                      
logic           [25:0]  mpp_gpolring_in_4_1;                      
logic           [25:0]  mpp_gpolring_in_5_0;                      
logic           [25:0]  mpp_gpolring_in_5_1;                      
logic           [25:0]  mpp_gpolring_in_6_0;                      
logic           [25:0]  mpp_gpolring_in_6_1;                      
logic           [25:0]  mpp_gpolring_in_7_0;                      
logic           [25:0]  mpp_gpolring_in_7_1;                      
logic          [106:0]  mpp_gpolring_update_in_0;                 
logic          [106:0]  mpp_gpolring_update_in_1;                 
logic           [68:0]  mpp_mctagring_in_0;                       
logic           [68:0]  mpp_mctagring_in_1;                       
logic           [68:0]  mpp_mctagring_in_2;                       
logic           [68:0]  mpp_mctagring_in_3;                       
logic           [33:0]  mpp_mrpodring_in_dn;                      
logic           [33:0]  mpp_mrpodring_in_up;                      
logic                   mpp_mrpodring_stall_in_dn;                
logic                   mpp_mrpodring_stall_in_up;                
logic           [33:0]  mpp_podring_in_dn;                        
logic           [33:0]  mpp_podring_in_up;                        
logic                   mpp_podring_stall_in_dn;                  
logic                   mpp_podring_stall_in_up;                  
logic           [67:0]  mpp_tagring_in_dn_0_0;                    
logic           [67:0]  mpp_tagring_in_dn_0_1;                    
logic           [67:0]  mpp_tagring_in_dn_10_0;                   
logic           [67:0]  mpp_tagring_in_dn_10_1;                   
logic           [67:0]  mpp_tagring_in_dn_11_0;                   
logic           [67:0]  mpp_tagring_in_dn_11_1;                   
logic           [67:0]  mpp_tagring_in_dn_12_0;                   
logic           [67:0]  mpp_tagring_in_dn_12_1;                   
logic           [67:0]  mpp_tagring_in_dn_13_0;                   
logic           [67:0]  mpp_tagring_in_dn_13_1;                   
logic           [67:0]  mpp_tagring_in_dn_14_0;                   
logic           [67:0]  mpp_tagring_in_dn_14_1;                   
logic           [67:0]  mpp_tagring_in_dn_15_0;                   
logic           [67:0]  mpp_tagring_in_dn_15_1;                   
logic           [67:0]  mpp_tagring_in_dn_1_0;                    
logic           [67:0]  mpp_tagring_in_dn_1_1;                    
logic           [67:0]  mpp_tagring_in_dn_2_0;                    
logic           [67:0]  mpp_tagring_in_dn_2_1;                    
logic           [67:0]  mpp_tagring_in_dn_3_0;                    
logic           [67:0]  mpp_tagring_in_dn_3_1;                    
logic           [67:0]  mpp_tagring_in_dn_4_0;                    
logic           [67:0]  mpp_tagring_in_dn_4_1;                    
logic           [67:0]  mpp_tagring_in_dn_5_0;                    
logic           [67:0]  mpp_tagring_in_dn_5_1;                    
logic           [67:0]  mpp_tagring_in_dn_6_0;                    
logic           [67:0]  mpp_tagring_in_dn_6_1;                    
logic           [67:0]  mpp_tagring_in_dn_7_0;                    
logic           [67:0]  mpp_tagring_in_dn_7_1;                    
logic           [67:0]  mpp_tagring_in_dn_8_0;                    
logic           [67:0]  mpp_tagring_in_dn_8_1;                    
logic           [67:0]  mpp_tagring_in_dn_9_0;                    
logic           [67:0]  mpp_tagring_in_dn_9_1;                    
logic           [67:0]  mpp_tagring_in_up_0_0;                    
logic           [67:0]  mpp_tagring_in_up_0_1;                    
logic           [67:0]  mpp_tagring_in_up_10_0;                   
logic           [67:0]  mpp_tagring_in_up_10_1;                   
logic           [67:0]  mpp_tagring_in_up_11_0;                   
logic           [67:0]  mpp_tagring_in_up_11_1;                   
logic           [67:0]  mpp_tagring_in_up_12_0;                   
logic           [67:0]  mpp_tagring_in_up_12_1;                   
logic           [67:0]  mpp_tagring_in_up_13_0;                   
logic           [67:0]  mpp_tagring_in_up_13_1;                   
logic           [67:0]  mpp_tagring_in_up_14_0;                   
logic           [67:0]  mpp_tagring_in_up_14_1;                   
logic           [67:0]  mpp_tagring_in_up_15_0;                   
logic           [67:0]  mpp_tagring_in_up_15_1;                   
logic           [67:0]  mpp_tagring_in_up_1_0;                    
logic           [67:0]  mpp_tagring_in_up_1_1;                    
logic           [67:0]  mpp_tagring_in_up_2_0;                    
logic           [67:0]  mpp_tagring_in_up_2_1;                    
logic           [67:0]  mpp_tagring_in_up_3_0;                    
logic           [67:0]  mpp_tagring_in_up_3_1;                    
logic           [67:0]  mpp_tagring_in_up_4_0;                    
logic           [67:0]  mpp_tagring_in_up_4_1;                    
logic           [67:0]  mpp_tagring_in_up_5_0;                    
logic           [67:0]  mpp_tagring_in_up_5_1;                    
logic           [67:0]  mpp_tagring_in_up_6_0;                    
logic           [67:0]  mpp_tagring_in_up_6_1;                    
logic           [67:0]  mpp_tagring_in_up_7_0;                    
logic           [67:0]  mpp_tagring_in_up_7_1;                    
logic           [67:0]  mpp_tagring_in_up_8_0;                    
logic           [67:0]  mpp_tagring_in_up_8_1;                    
logic           [67:0]  mpp_tagring_in_up_9_0;                    
logic           [67:0]  mpp_tagring_in_up_9_1;                    
//edr logic           [31:0]  i_reqAddr;                                
//edr logic            [7:0]  i_reqID;                                  // from iMC axi 
//edr logic                   i_reqParity;                              // odd parity bit to cover req 
//edr logic                   i_reqValid;                               
//edr logic                   i_reqWr;                                  // '0'= read 
//edr logic           [63:0]  i_reqWrData;                              
logic                   sreset;                                   
logic           [39:0]  grp_d0_rx_time_stamp;           
logic           [63:0]  grp_b0_rx5_data;                
logic           [63:0]  grp_d1_rx3_data;                
logic           [63:0]  grp_d0_rx0_data;                
logic           [39:0]  grp_a1_rx_time_stamp;           
logic           [63:0]  grp_b1_rx3_data;                
logic           [63:0]  grp_c0_rx4_data;                
logic           [63:0]  grp_b1_rx7_data;                
logic           [71:0]  igr1_vp_rx5_data_w_ecc;         
logic           [63:0]  grp_c0_rx7_data;                
logic           [63:0]  grp_c1_rx7_data;                
logic           [63:0]  grp_a1_rx0_data;                
logic           [23:0]  grp_a0_rx_metadata;             
logic           [63:0]  grp_c1_rx3_data;                
logic           [63:0]  grp_d0_rx4_data;                
logic           [63:0]  grp_a1_rx1_data;                
logic           [63:0]  grp_c1_rx6_data;                
logic           [63:0]  grp_c1_rx2_data;                
logic           [63:0]  grp_c0_rx2_data;                
logic           [63:0]  grp_a0_rx5_data;                
logic           [63:0]  grp_c0_rx3_data;                
logic           [71:0]  igr1_vp_rx0_data_w_ecc;         
logic           [71:0]  igr0_vp_rx7_data_w_ecc;         
logic           [63:0]  grp_b1_rx6_data;                
logic           [71:0]  igr1_vp_rx2_data_w_ecc;         
logic           [63:0]  grp_d0_rx3_data;                
logic           [63:0]  grp_a0_rx3_data;                
logic           [63:0]  grp_b1_rx1_data;                
logic           [63:0]  grp_a0_rx6_data;                
logic           [63:0]  grp_c0_rx0_data;                
logic           [63:0]  grp_c0_rx6_data;                
logic           [71:0]  igr0_vp_rx4_data_w_ecc;         
logic           [63:0]  grp_a1_rx6_data;                
logic           [23:0]  grp_c1_rx_metadata;             
logic           [63:0]  grp_a0_rx2_data;                
logic           [63:0]  grp_d0_rx1_data;                
logic           [71:0]  igr1_vp_rx1_data_w_ecc;         
logic           [39:0]  grp_c1_rx_time_stamp;           
logic           [63:0]  grp_a1_rx7_data;                
logic           [63:0]  grp_d1_rx6_data;                
logic           [63:0]  grp_a1_rx3_data;                
logic           [63:0]  grp_a0_rx1_data;                
logic           [63:0]  grp_b0_rx2_data;                
logic           [39:0]  grp_d1_rx_time_stamp;           
logic           [63:0]  grp_d1_rx4_data;                
logic           [63:0]  grp_c1_rx0_data;                
logic           [39:0]  grp_c0_rx_time_stamp;           
logic            [2:0]  mpp_id;                         
logic           [71:0]  igr1_vp_rx7_data_w_ecc;         
logic           [23:0]  grp_b1_rx_metadata;             
logic           [63:0]  grp_b1_rx4_data;                
logic           [63:0]  grp_d1_rx1_data;                
logic           [63:0]  grp_d0_rx5_data;                
logic           [39:0]  grp_b1_rx_time_stamp;           
logic           [63:0]  grp_b0_rx0_data;                
logic           [63:0]  grp_b0_rx6_data;                
logic           [63:0]  grp_d0_rx6_data;                
logic           [63:0]  grp_c1_rx4_data;                
logic           [63:0]  grp_c0_rx5_data;                
logic           [39:0]  grp_a0_rx_time_stamp;           
logic           [63:0]  grp_b1_rx2_data;                
logic           [63:0]  grp_a1_rx2_data;                
logic           [63:0]  grp_c0_rx1_data;                
logic           [63:0]  grp_a0_rx0_data;                
logic           [71:0]  igr1_vp_rx6_data_w_ecc;         
logic           [63:0]  grp_b0_rx7_data;                
logic           [71:0]  igr1_vp_rx3_data_w_ecc;         
logic           [63:0]  grp_b0_rx3_data;                
logic           [23:0]  grp_d1_rx_metadata;             
logic           [23:0]  grp_a1_rx_metadata;             
logic           [63:0]  grp_d0_rx2_data;                
logic           [63:0]  grp_d1_rx2_data;                
logic           [63:0]  grp_d1_rx7_data;                
logic           [23:0]  grp_b0_rx_metadata;             
logic           [23:0]  grp_c0_rx_metadata;             
logic           [23:0]  grp_d0_rx_metadata;             
logic           [63:0]  grp_d0_rx7_data;                
logic           [63:0]  grp_b1_rx0_data;                
logic           [71:0]  igr0_vp_rx0_data_w_ecc;         
logic           [63:0]  grp_c1_rx1_data;                
logic           [39:0]  grp_b0_rx_time_stamp;           
logic           [63:0]  grp_b1_rx5_data;                
logic           [63:0]  grp_d1_rx5_data;                
logic           [63:0]  grp_a0_rx7_data;                
logic           [63:0]  grp_b0_rx1_data;                
logic           [71:0]  igr1_vp_rx4_data_w_ecc;         
logic           [63:0]  grp_d1_rx0_data;                
logic           [63:0]  grp_a0_rx4_data;                
logic           [71:0]  igr0_vp_rx2_data_w_ecc;         
logic           [63:0]  grp_b0_rx4_data;                
logic           [71:0]  igr0_vp_rx6_data_w_ecc;         
logic           [71:0]  igr0_vp_rx1_data_w_ecc;         
logic           [63:0]  grp_c1_rx5_data;                
logic           [71:0]  igr0_vp_rx3_data_w_ecc;         
logic           [71:0]  igr0_vp_rx5_data_w_ecc;         
logic           [63:0]  grp_a1_rx4_data;                
logic           [63:0]  grp_a1_rx5_data;                

//Interface List
logic            ahb0_rxppe_ahb_sel;              // Blasted Interface ahb_rx_ppe_if.ppe ahb0_rxppe
logic            ahb0_rxppe_ahb_wr;              
logic  [shared_pkg::W_MGMT_ADDR-1:0]  ahb0_rxppe_ahb_addr;            
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb0_rxppe_ahb_wr_data;         
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb0_rxppe_ahb_rd_data;         
logic            ahb0_rxppe_ahb_rd_ack;          

logic            ahb0_txppe0_ahb_sel;              // Blasted Interface ahb_rx_ppe_if.ppe ahb0_txppe0
logic            ahb0_txppe0_ahb_wr;             
logic  [shared_pkg::W_MGMT_ADDR-1:0]  ahb0_txppe0_ahb_addr;           
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb0_txppe0_ahb_wr_data;        
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb0_txppe0_ahb_rd_data;        
logic            ahb0_txppe0_ahb_rd_ack;         

logic            ahb0_txppe1_ahb_sel;              // Blasted Interface ahb_rx_ppe_if.ppe ahb0_txppe1
logic            ahb0_txppe1_ahb_wr;             
logic  [shared_pkg::W_MGMT_ADDR-1:0]  ahb0_txppe1_ahb_addr;           
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb0_txppe1_ahb_wr_data;        
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb0_txppe1_ahb_rd_data;        
logic            ahb0_txppe1_ahb_rd_ack;         

logic            ahb1_rxppe_ahb_sel;              // Blasted Interface ahb_rx_ppe_if.ppe ahb1_rxppe
logic            ahb1_rxppe_ahb_wr;              
logic  [shared_pkg::W_MGMT_ADDR-1:0]  ahb1_rxppe_ahb_addr;            
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb1_rxppe_ahb_wr_data;         
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb1_rxppe_ahb_rd_data;         
logic            ahb1_rxppe_ahb_rd_ack;          

logic            ahb1_txppe0_ahb_sel;              // Blasted Interface ahb_rx_ppe_if.ppe ahb1_txppe0
logic            ahb1_txppe0_ahb_wr;             
logic  [shared_pkg::W_MGMT_ADDR-1:0]  ahb1_txppe0_ahb_addr;           
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb1_txppe0_ahb_wr_data;        
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb1_txppe0_ahb_rd_data;        
logic            ahb1_txppe0_ahb_rd_ack;         

logic            ahb1_txppe1_ahb_sel;              // Blasted Interface ahb_rx_ppe_if.ppe ahb1_txppe1
logic            ahb1_txppe1_ahb_wr;             
logic  [shared_pkg::W_MGMT_ADDR-1:0]  ahb1_txppe1_ahb_addr;           
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb1_txppe1_ahb_wr_data;        
logic  [shared_pkg::W_MGMT_DATA64-1:0]  ahb1_txppe1_ahb_rd_data;        
logic            ahb1_txppe1_ahb_rd_ack;         

logic            egr0_ahb_ahb_req_p;              // Blasted Interface egr_ahb_if.egr egr0_ahb
logic  [W_AHB_ADDR-1:0]  egr0_ahb_ahb_addr;              
logic            egr0_ahb_ahb_wr;                
logic  [W_AHB_DATA-1:0]  egr0_ahb_ahb_wr_data;           
logic            egr0_ahb_ahb_ack_p;             
logic  [W_AHB_DATA-1:0]  egr0_ahb_ahb_rd_data;           
logic            egr0_ahb_dfxsignal_in;          
logic            egr0_ahb_dfxsignal_out;         

logic            egr1_ahb_ahb_req_p;              // Blasted Interface egr_ahb_if.egr egr1_ahb
logic  [W_AHB_ADDR-1:0]  egr1_ahb_ahb_addr;              
logic            egr1_ahb_ahb_wr;                
logic  [W_AHB_DATA-1:0]  egr1_ahb_ahb_wr_data;           
logic            egr1_ahb_ahb_ack_p;             
logic  [W_AHB_DATA-1:0]  egr1_ahb_ahb_rd_data;           
logic            egr1_ahb_dfxsignal_in;          
logic            egr1_ahb_dfxsignal_out;         

logic            glb0_rxppe_glb_sync;              // Blasted Interface glb_rx_ppe_if.ppe glb0_rxppe
logic            glb0_rxppe_glb_ack;             

logic            glb0_txppe0_glb_sync;              // Blasted Interface glb_rx_ppe_if.ppe glb0_txppe0
logic            glb0_txppe0_glb_ack;            

logic            glb0_txppe1_glb_sync;              // Blasted Interface glb_rx_ppe_if.ppe glb0_txppe1
logic            glb0_txppe1_glb_ack;            

logic            glb1_rxppe_glb_sync;              // Blasted Interface glb_rx_ppe_if.ppe glb1_rxppe
logic            glb1_rxppe_glb_ack;             

logic            glb1_txppe0_glb_sync;              // Blasted Interface glb_rx_ppe_if.ppe glb1_txppe0
logic            glb1_txppe0_glb_ack;            

logic            glb1_txppe1_glb_sync;              // Blasted Interface glb_rx_ppe_if.ppe glb1_txppe1
logic            glb1_txppe1_glb_ack;            

logic     [1:0]  grp_a0_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_a0
logic            grp_a0_tx_enable;               
logic     [7:0]  grp_a0_tx_data_valid;           
logic     [1:0]  grp_a0_tx_port_num;             
logic            grp_a0_tx_valid_resp;           
logic    [23:0]  grp_a0_tx_metadata;             
logic    [63:0]  grp_a0_tx0_data;                
logic    [63:0]  grp_a0_tx1_data;                
logic    [63:0]  grp_a0_tx2_data;                
logic    [63:0]  grp_a0_tx3_data;                
logic    [63:0]  grp_a0_tx4_data;                
logic    [63:0]  grp_a0_tx5_data;                
logic    [63:0]  grp_a0_tx6_data;                
logic    [63:0]  grp_a0_tx7_data;                
logic     [3:0]  grp_a0_rx_pfc_xoff;             
logic            grp_a0_rx_pfc_tc_sync;          

logic     [1:0]  grp_a1_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_a1
logic            grp_a1_tx_enable;               
logic     [7:0]  grp_a1_tx_data_valid;           
logic     [1:0]  grp_a1_tx_port_num;             
logic            grp_a1_tx_valid_resp;           
logic    [23:0]  grp_a1_tx_metadata;             
logic    [63:0]  grp_a1_tx0_data;                
logic    [63:0]  grp_a1_tx1_data;                
logic    [63:0]  grp_a1_tx2_data;                
logic    [63:0]  grp_a1_tx3_data;                
logic    [63:0]  grp_a1_tx4_data;                
logic    [63:0]  grp_a1_tx5_data;                
logic    [63:0]  grp_a1_tx6_data;                
logic    [63:0]  grp_a1_tx7_data;                
logic     [3:0]  grp_a1_rx_pfc_xoff;             
logic            grp_a1_rx_pfc_tc_sync;          

logic     [1:0]  grp_b0_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_b0
logic            grp_b0_tx_enable;               
logic     [7:0]  grp_b0_tx_data_valid;           
logic     [1:0]  grp_b0_tx_port_num;             
logic            grp_b0_tx_valid_resp;           
logic    [23:0]  grp_b0_tx_metadata;             
logic    [63:0]  grp_b0_tx0_data;                
logic    [63:0]  grp_b0_tx1_data;                
logic    [63:0]  grp_b0_tx2_data;                
logic    [63:0]  grp_b0_tx3_data;                
logic    [63:0]  grp_b0_tx4_data;                
logic    [63:0]  grp_b0_tx5_data;                
logic    [63:0]  grp_b0_tx6_data;                
logic    [63:0]  grp_b0_tx7_data;                
logic     [3:0]  grp_b0_rx_pfc_xoff;             
logic            grp_b0_rx_pfc_tc_sync;          

logic     [1:0]  grp_b1_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_b1
logic            grp_b1_tx_enable;               
logic     [7:0]  grp_b1_tx_data_valid;           
logic     [1:0]  grp_b1_tx_port_num;             
logic            grp_b1_tx_valid_resp;           
logic    [23:0]  grp_b1_tx_metadata;             
logic    [63:0]  grp_b1_tx0_data;                
logic    [63:0]  grp_b1_tx1_data;                
logic    [63:0]  grp_b1_tx2_data;                
logic    [63:0]  grp_b1_tx3_data;                
logic    [63:0]  grp_b1_tx4_data;                
logic    [63:0]  grp_b1_tx5_data;                
logic    [63:0]  grp_b1_tx6_data;                
logic    [63:0]  grp_b1_tx7_data;                
logic     [3:0]  grp_b1_rx_pfc_xoff;             
logic            grp_b1_rx_pfc_tc_sync;          

logic     [1:0]  grp_c0_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_c0
logic            grp_c0_tx_enable;               
logic     [7:0]  grp_c0_tx_data_valid;           
logic     [1:0]  grp_c0_tx_port_num;             
logic            grp_c0_tx_valid_resp;           
logic    [23:0]  grp_c0_tx_metadata;             
logic    [63:0]  grp_c0_tx0_data;                
logic    [63:0]  grp_c0_tx1_data;                
logic    [63:0]  grp_c0_tx2_data;                
logic    [63:0]  grp_c0_tx3_data;                
logic    [63:0]  grp_c0_tx4_data;                
logic    [63:0]  grp_c0_tx5_data;                
logic    [63:0]  grp_c0_tx6_data;                
logic    [63:0]  grp_c0_tx7_data;                
logic     [3:0]  grp_c0_rx_pfc_xoff;             
logic            grp_c0_rx_pfc_tc_sync;          

logic     [1:0]  grp_c1_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_c1
logic            grp_c1_tx_enable;               
logic     [7:0]  grp_c1_tx_data_valid;           
logic     [1:0]  grp_c1_tx_port_num;             
logic            grp_c1_tx_valid_resp;           
logic    [23:0]  grp_c1_tx_metadata;             
logic    [63:0]  grp_c1_tx0_data;                
logic    [63:0]  grp_c1_tx1_data;                
logic    [63:0]  grp_c1_tx2_data;                
logic    [63:0]  grp_c1_tx3_data;                
logic    [63:0]  grp_c1_tx4_data;                
logic    [63:0]  grp_c1_tx5_data;                
logic    [63:0]  grp_c1_tx6_data;                
logic    [63:0]  grp_c1_tx7_data;                
logic     [3:0]  grp_c1_rx_pfc_xoff;             
logic            grp_c1_rx_pfc_tc_sync;          

logic     [1:0]  grp_d0_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_d0
logic            grp_d0_tx_enable;               
logic     [7:0]  grp_d0_tx_data_valid;           
logic     [1:0]  grp_d0_tx_port_num;             
logic            grp_d0_tx_valid_resp;           
logic    [23:0]  grp_d0_tx_metadata;             
logic    [63:0]  grp_d0_tx0_data;                
logic    [63:0]  grp_d0_tx1_data;                
logic    [63:0]  grp_d0_tx2_data;                
logic    [63:0]  grp_d0_tx3_data;                
logic    [63:0]  grp_d0_tx4_data;                
logic    [63:0]  grp_d0_tx5_data;                
logic    [63:0]  grp_d0_tx6_data;                
logic    [63:0]  grp_d0_tx7_data;                
logic     [3:0]  grp_d0_rx_pfc_xoff;             
logic            grp_d0_rx_pfc_tc_sync;          

logic     [1:0]  grp_d1_tx_enable_port_num;              // Blasted Interface egr_epl_if.egr grp_d1
logic            grp_d1_tx_enable;               
logic     [7:0]  grp_d1_tx_data_valid;           
logic     [1:0]  grp_d1_tx_port_num;             
logic            grp_d1_tx_valid_resp;           
logic    [23:0]  grp_d1_tx_metadata;             
logic    [63:0]  grp_d1_tx0_data;                
logic    [63:0]  grp_d1_tx1_data;                
logic    [63:0]  grp_d1_tx2_data;                
logic    [63:0]  grp_d1_tx3_data;                
logic    [63:0]  grp_d1_tx4_data;                
logic    [63:0]  grp_d1_tx5_data;                
logic    [63:0]  grp_d1_tx6_data;                
logic    [63:0]  grp_d1_tx7_data;                
logic     [3:0]  grp_d1_rx_pfc_xoff;             
logic            grp_d1_rx_pfc_tc_sync;          

logic            mim0_rd0_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim0_rd0
logic  [20-1:0]  mim0_rd0_mim_seg_ptr;           
logic   [4-1:0]  mim0_rd0_mim_sema;              
logic   [2-1:0]  mim0_rd0_mim_wd_sel;            
logic  [13-1:0]  mim0_rd0_mim_req_id;            
logic   [1-1:0]  mim0_rd0_mim_rreq_credits;      
logic            mim0_rd0_mim_rrsp_valid;        
logic   [3-1:0]  mim0_rd0_mim_rrsp_dest_block;   
logic  [13-1:0]  mim0_rd0_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim0_rd0_mim_rd_data;           

logic            mim0_rd1_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim0_rd1
logic  [20-1:0]  mim0_rd1_mim_seg_ptr;           
logic   [4-1:0]  mim0_rd1_mim_sema;              
logic   [2-1:0]  mim0_rd1_mim_wd_sel;            
logic  [13-1:0]  mim0_rd1_mim_req_id;            
logic   [1-1:0]  mim0_rd1_mim_rreq_credits;      
logic            mim0_rd1_mim_rrsp_valid;        
logic   [3-1:0]  mim0_rd1_mim_rrsp_dest_block;   
logic  [13-1:0]  mim0_rd1_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim0_rd1_mim_rd_data;           

logic            mim0_rd2_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim0_rd2
logic  [20-1:0]  mim0_rd2_mim_seg_ptr;           
logic   [4-1:0]  mim0_rd2_mim_sema;              
logic   [2-1:0]  mim0_rd2_mim_wd_sel;            
logic  [13-1:0]  mim0_rd2_mim_req_id;            
logic   [1-1:0]  mim0_rd2_mim_rreq_credits;      
logic            mim0_rd2_mim_rrsp_valid;        
logic   [3-1:0]  mim0_rd2_mim_rrsp_dest_block;   
logic  [13-1:0]  mim0_rd2_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim0_rd2_mim_rd_data;           

logic            mim0_wr0_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim0_wr0
logic  [20-1:0]  mim0_wr0_mim_wr_seg_ptr;        
logic   [4-1:0]  mim0_wr0_mim_wr_sema;           
logic   [2-1:0]  mim0_wr0_mim_wr_wd_sel;         
logic  [13-1:0]  mim0_wr0_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim0_wr0_mim_wr_data;           
logic   [1-1:0]  mim0_wr0_mim_wreq_credits;      

logic            mim0_wr1_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim0_wr1
logic  [20-1:0]  mim0_wr1_mim_wr_seg_ptr;        
logic   [4-1:0]  mim0_wr1_mim_wr_sema;           
logic   [2-1:0]  mim0_wr1_mim_wr_wd_sel;         
logic  [13-1:0]  mim0_wr1_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim0_wr1_mim_wr_data;           
logic   [1-1:0]  mim0_wr1_mim_wreq_credits;      

logic            mim0_wr2_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim0_wr2
logic  [20-1:0]  mim0_wr2_mim_wr_seg_ptr;        
logic   [4-1:0]  mim0_wr2_mim_wr_sema;           
logic   [2-1:0]  mim0_wr2_mim_wr_wd_sel;         
logic  [13-1:0]  mim0_wr2_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim0_wr2_mim_wr_data;           
logic   [1-1:0]  mim0_wr2_mim_wreq_credits;      

logic            mim1_rd0_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim1_rd0
logic  [20-1:0]  mim1_rd0_mim_seg_ptr;           
logic   [4-1:0]  mim1_rd0_mim_sema;              
logic   [2-1:0]  mim1_rd0_mim_wd_sel;            
logic  [13-1:0]  mim1_rd0_mim_req_id;            
logic   [1-1:0]  mim1_rd0_mim_rreq_credits;      
logic            mim1_rd0_mim_rrsp_valid;        
logic   [3-1:0]  mim1_rd0_mim_rrsp_dest_block;   
logic  [13-1:0]  mim1_rd0_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim1_rd0_mim_rd_data;           

logic            mim1_rd1_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim1_rd1
logic  [20-1:0]  mim1_rd1_mim_seg_ptr;           
logic   [4-1:0]  mim1_rd1_mim_sema;              
logic   [2-1:0]  mim1_rd1_mim_wd_sel;            
logic  [13-1:0]  mim1_rd1_mim_req_id;            
logic   [1-1:0]  mim1_rd1_mim_rreq_credits;      
logic            mim1_rd1_mim_rrsp_valid;        
logic   [3-1:0]  mim1_rd1_mim_rrsp_dest_block;   
logic  [13-1:0]  mim1_rd1_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim1_rd1_mim_rd_data;           

logic            mim1_rd2_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim1_rd2
logic  [20-1:0]  mim1_rd2_mim_seg_ptr;           
logic   [4-1:0]  mim1_rd2_mim_sema;              
logic   [2-1:0]  mim1_rd2_mim_wd_sel;            
logic  [13-1:0]  mim1_rd2_mim_req_id;            
logic   [1-1:0]  mim1_rd2_mim_rreq_credits;      
logic            mim1_rd2_mim_rrsp_valid;        
logic   [3-1:0]  mim1_rd2_mim_rrsp_dest_block;   
logic  [13-1:0]  mim1_rd2_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim1_rd2_mim_rd_data;           

logic            mim1_wr0_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim1_wr0
logic  [20-1:0]  mim1_wr0_mim_wr_seg_ptr;        
logic   [4-1:0]  mim1_wr0_mim_wr_sema;           
logic   [2-1:0]  mim1_wr0_mim_wr_wd_sel;         
logic  [13-1:0]  mim1_wr0_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim1_wr0_mim_wr_data;           
logic   [1-1:0]  mim1_wr0_mim_wreq_credits;      

logic            mim1_wr1_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim1_wr1
logic  [20-1:0]  mim1_wr1_mim_wr_seg_ptr;        
logic   [4-1:0]  mim1_wr1_mim_wr_sema;           
logic   [2-1:0]  mim1_wr1_mim_wr_wd_sel;         
logic  [13-1:0]  mim1_wr1_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim1_wr1_mim_wr_data;           
logic   [1-1:0]  mim1_wr1_mim_wreq_credits;      

logic            mim1_wr2_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim1_wr2
logic  [20-1:0]  mim1_wr2_mim_wr_seg_ptr;        
logic   [4-1:0]  mim1_wr2_mim_wr_sema;           
logic   [2-1:0]  mim1_wr2_mim_wr_wd_sel;         
logic  [13-1:0]  mim1_wr2_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim1_wr2_mim_wr_data;           
logic   [1-1:0]  mim1_wr2_mim_wreq_credits;      

logic            mim2_rd0_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim2_rd0
logic  [20-1:0]  mim2_rd0_mim_seg_ptr;           
logic   [4-1:0]  mim2_rd0_mim_sema;              
logic   [2-1:0]  mim2_rd0_mim_wd_sel;            
logic  [13-1:0]  mim2_rd0_mim_req_id;            
logic   [1-1:0]  mim2_rd0_mim_rreq_credits;      
logic            mim2_rd0_mim_rrsp_valid;        
logic   [3-1:0]  mim2_rd0_mim_rrsp_dest_block;   
logic  [13-1:0]  mim2_rd0_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim2_rd0_mim_rd_data;           

logic            mim2_rd1_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim2_rd1
logic  [20-1:0]  mim2_rd1_mim_seg_ptr;           
logic   [4-1:0]  mim2_rd1_mim_sema;              
logic   [2-1:0]  mim2_rd1_mim_wd_sel;            
logic  [13-1:0]  mim2_rd1_mim_req_id;            
logic   [1-1:0]  mim2_rd1_mim_rreq_credits;      
logic            mim2_rd1_mim_rrsp_valid;        
logic   [3-1:0]  mim2_rd1_mim_rrsp_dest_block;   
logic  [13-1:0]  mim2_rd1_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim2_rd1_mim_rd_data;           

logic            mim2_rd2_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim2_rd2
logic  [20-1:0]  mim2_rd2_mim_seg_ptr;           
logic   [4-1:0]  mim2_rd2_mim_sema;              
logic   [2-1:0]  mim2_rd2_mim_wd_sel;            
logic  [13-1:0]  mim2_rd2_mim_req_id;            
logic   [1-1:0]  mim2_rd2_mim_rreq_credits;      
logic            mim2_rd2_mim_rrsp_valid;        
logic   [3-1:0]  mim2_rd2_mim_rrsp_dest_block;   
logic  [13-1:0]  mim2_rd2_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim2_rd2_mim_rd_data;           

logic            mim2_wr0_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim2_wr0
logic  [20-1:0]  mim2_wr0_mim_wr_seg_ptr;        
logic   [4-1:0]  mim2_wr0_mim_wr_sema;           
logic   [2-1:0]  mim2_wr0_mim_wr_wd_sel;         
logic  [13-1:0]  mim2_wr0_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim2_wr0_mim_wr_data;           
logic   [1-1:0]  mim2_wr0_mim_wreq_credits;      

logic            mim2_wr1_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim2_wr1
logic  [20-1:0]  mim2_wr1_mim_wr_seg_ptr;        
logic   [4-1:0]  mim2_wr1_mim_wr_sema;           
logic   [2-1:0]  mim2_wr1_mim_wr_wd_sel;         
logic  [13-1:0]  mim2_wr1_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim2_wr1_mim_wr_data;           
logic   [1-1:0]  mim2_wr1_mim_wreq_credits;      

logic            mim2_wr2_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim2_wr2
logic  [20-1:0]  mim2_wr2_mim_wr_seg_ptr;        
logic   [4-1:0]  mim2_wr2_mim_wr_sema;           
logic   [2-1:0]  mim2_wr2_mim_wr_wd_sel;         
logic  [13-1:0]  mim2_wr2_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim2_wr2_mim_wr_data;           
logic   [1-1:0]  mim2_wr2_mim_wreq_credits;      

logic            mim3_rd0_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim3_rd0
logic  [20-1:0]  mim3_rd0_mim_seg_ptr;           
logic   [4-1:0]  mim3_rd0_mim_sema;              
logic   [2-1:0]  mim3_rd0_mim_wd_sel;            
logic  [13-1:0]  mim3_rd0_mim_req_id;            
logic   [1-1:0]  mim3_rd0_mim_rreq_credits;      
logic            mim3_rd0_mim_rrsp_valid;        
logic   [3-1:0]  mim3_rd0_mim_rrsp_dest_block;   
logic  [13-1:0]  mim3_rd0_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim3_rd0_mim_rd_data;           

logic            mim3_rd1_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim3_rd1
logic  [20-1:0]  mim3_rd1_mim_seg_ptr;           
logic   [4-1:0]  mim3_rd1_mim_sema;              
logic   [2-1:0]  mim3_rd1_mim_wd_sel;            
logic  [13-1:0]  mim3_rd1_mim_req_id;            
logic   [1-1:0]  mim3_rd1_mim_rreq_credits;      
logic            mim3_rd1_mim_rrsp_valid;        
logic   [3-1:0]  mim3_rd1_mim_rrsp_dest_block;   
logic  [13-1:0]  mim3_rd1_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim3_rd1_mim_rd_data;           

logic            mim3_rd2_mim_rreq_valid;              // Blasted Interface mim_rd_if.request mim3_rd2
logic  [20-1:0]  mim3_rd2_mim_seg_ptr;           
logic   [4-1:0]  mim3_rd2_mim_sema;              
logic   [2-1:0]  mim3_rd2_mim_wd_sel;            
logic  [13-1:0]  mim3_rd2_mim_req_id;            
logic   [1-1:0]  mim3_rd2_mim_rreq_credits;      
logic            mim3_rd2_mim_rrsp_valid;        
logic   [3-1:0]  mim3_rd2_mim_rrsp_dest_block;   
logic  [13-1:0]  mim3_rd2_mim_rrsp_req_id;       
logic  [W_WORD_BITS-1:0]  mim3_rd2_mim_rd_data;           

logic            mim3_wr0_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim3_wr0
logic  [20-1:0]  mim3_wr0_mim_wr_seg_ptr;        
logic   [4-1:0]  mim3_wr0_mim_wr_sema;           
logic   [2-1:0]  mim3_wr0_mim_wr_wd_sel;         
logic  [13-1:0]  mim3_wr0_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim3_wr0_mim_wr_data;           
logic   [1-1:0]  mim3_wr0_mim_wreq_credits;      

logic            mim3_wr1_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim3_wr1
logic  [20-1:0]  mim3_wr1_mim_wr_seg_ptr;        
logic   [4-1:0]  mim3_wr1_mim_wr_sema;           
logic   [2-1:0]  mim3_wr1_mim_wr_wd_sel;         
logic  [13-1:0]  mim3_wr1_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim3_wr1_mim_wr_data;           
logic   [1-1:0]  mim3_wr1_mim_wreq_credits;      

logic            mim3_wr2_mim_wreq_valid;              // Blasted Interface mim_wr_if.request mim3_wr2
logic  [20-1:0]  mim3_wr2_mim_wr_seg_ptr;        
logic   [4-1:0]  mim3_wr2_mim_wr_sema;           
logic   [2-1:0]  mim3_wr2_mim_wr_wd_sel;         
logic  [13-1:0]  mim3_wr2_mim_wreq_id;           
logic  [W_WORD_BITS-1:0]  mim3_wr2_mim_wr_data;           
logic   [1-1:0]  mim3_wr2_mim_wreq_credits;      


//Logic List
logic                  grp_a0_tx_pfc_tc_sync;                    
logic           [3:0]  grp_a0_tx_pfc_xoff;                       
logic                  grp_a1_tx_pfc_tc_sync;                    
logic           [3:0]  grp_a1_tx_pfc_xoff;                       
logic                  grp_b0_tx_pfc_tc_sync;                    
logic           [3:0]  grp_b0_tx_pfc_xoff;                       
logic                  grp_b1_tx_pfc_tc_sync;                    
logic           [3:0]  grp_b1_tx_pfc_xoff;                       
logic                  grp_c0_tx_pfc_tc_sync;                    
logic           [3:0]  grp_c0_tx_pfc_xoff;                       
logic                  grp_c1_tx_pfc_tc_sync;                    
logic           [3:0]  grp_c1_tx_pfc_xoff;                       
logic                  grp_d0_tx_pfc_tc_sync;                    
logic           [3:0]  grp_d0_tx_pfc_xoff;                       
logic                  grp_d1_tx_pfc_tc_sync;                    
logic           [3:0]  grp_d1_tx_pfc_xoff;                       
logic                  igr0_vp_tx_pfc_xoff;                      //FIXME should this be [1:0] for 2 VP   
logic                  igr1_vp_tx_pfc_xoff;                      //FIXME should this be [1:0] for 2 VP   
logic          [23:0]  mpp_dqring_out_0_0;                       
logic          [23:0]  mpp_dqring_out_0_1;                       
logic          [23:0]  mpp_dqring_out_1_0;                       
logic          [23:0]  mpp_dqring_out_1_1;                       
logic          [23:0]  mpp_dqring_out_2_0;                       
logic          [23:0]  mpp_dqring_out_2_1;                       
logic          [23:0]  mpp_dqring_out_3_0;                       
logic          [23:0]  mpp_dqring_out_3_1;                       
logic          [23:0]  mpp_dqring_out_4_0;                       
logic          [23:0]  mpp_dqring_out_4_1;                       
logic          [23:0]  mpp_dqring_out_5_0;                       
logic          [23:0]  mpp_dqring_out_5_1;                       
logic          [23:0]  mpp_dqring_out_6_0;                       
logic          [23:0]  mpp_dqring_out_6_1;                       
logic          [23:0]  mpp_dqring_out_7_0;                       
logic          [23:0]  mpp_dqring_out_7_1;                       
logic          [25:0]  mpp_gpolring_out_0_0;                     
logic          [25:0]  mpp_gpolring_out_0_1;                     
logic          [25:0]  mpp_gpolring_out_1_0;                     
logic          [25:0]  mpp_gpolring_out_1_1;                     
logic          [25:0]  mpp_gpolring_out_2_0;                     
logic          [25:0]  mpp_gpolring_out_2_1;                     
logic          [25:0]  mpp_gpolring_out_3_0;                     
logic          [25:0]  mpp_gpolring_out_3_1;                     
logic          [25:0]  mpp_gpolring_out_4_0;                     
logic          [25:0]  mpp_gpolring_out_4_1;                     
logic          [25:0]  mpp_gpolring_out_5_0;                     
logic          [25:0]  mpp_gpolring_out_5_1;                     
logic          [25:0]  mpp_gpolring_out_6_0;                     
logic          [25:0]  mpp_gpolring_out_6_1;                     
logic          [25:0]  mpp_gpolring_out_7_0;                     
logic          [25:0]  mpp_gpolring_out_7_1;                     
logic         [106:0]  mpp_gpolring_update_out_0;                
logic         [106:0]  mpp_gpolring_update_out_1;                
logic          [68:0]  mpp_mctagring_out_0;                      
logic          [68:0]  mpp_mctagring_out_1;                      
logic          [68:0]  mpp_mctagring_out_2;                      
logic          [68:0]  mpp_mctagring_out_3;                      
logic          [33:0]  mpp_mrpodring_out_dn;                     
logic          [33:0]  mpp_mrpodring_out_up;                     
logic                  mpp_mrpodring_stall_out_dn;               
logic                  mpp_mrpodring_stall_out_up;               
logic          [33:0]  mpp_podring_out_dn;                       
logic          [33:0]  mpp_podring_out_up;                       
logic                  mpp_podring_stall_out_dn;                 
logic                  mpp_podring_stall_out_up;                 
logic          [67:0]  mpp_tagring_out_dn_0_0;                   
logic          [67:0]  mpp_tagring_out_dn_0_1;                   
logic          [67:0]  mpp_tagring_out_dn_10_0;                  
logic          [67:0]  mpp_tagring_out_dn_10_1;                  
logic          [67:0]  mpp_tagring_out_dn_11_0;                  
logic          [67:0]  mpp_tagring_out_dn_11_1;                  
logic          [67:0]  mpp_tagring_out_dn_12_0;                  
logic          [67:0]  mpp_tagring_out_dn_12_1;                  
logic          [67:0]  mpp_tagring_out_dn_13_0;                  
logic          [67:0]  mpp_tagring_out_dn_13_1;                  
logic          [67:0]  mpp_tagring_out_dn_14_0;                  
logic          [67:0]  mpp_tagring_out_dn_14_1;                  
logic          [67:0]  mpp_tagring_out_dn_15_0;                  
logic          [67:0]  mpp_tagring_out_dn_15_1;                  
logic          [67:0]  mpp_tagring_out_dn_1_0;                   
logic          [67:0]  mpp_tagring_out_dn_1_1;                   
logic          [67:0]  mpp_tagring_out_dn_2_0;                   
logic          [67:0]  mpp_tagring_out_dn_2_1;                   
logic          [67:0]  mpp_tagring_out_dn_3_0;                   
logic          [67:0]  mpp_tagring_out_dn_3_1;                   
logic          [67:0]  mpp_tagring_out_dn_4_0;                   
logic          [67:0]  mpp_tagring_out_dn_4_1;                   
logic          [67:0]  mpp_tagring_out_dn_5_0;                   
logic          [67:0]  mpp_tagring_out_dn_5_1;                   
logic          [67:0]  mpp_tagring_out_dn_6_0;                   
logic          [67:0]  mpp_tagring_out_dn_6_1;                   
logic          [67:0]  mpp_tagring_out_dn_7_0;                   
logic          [67:0]  mpp_tagring_out_dn_7_1;                   
logic          [67:0]  mpp_tagring_out_dn_8_0;                   
logic          [67:0]  mpp_tagring_out_dn_8_1;                   
logic          [67:0]  mpp_tagring_out_dn_9_0;                   
logic          [67:0]  mpp_tagring_out_dn_9_1;                   
logic          [67:0]  mpp_tagring_out_up_0_0;                   
logic          [67:0]  mpp_tagring_out_up_0_1;                   
logic          [67:0]  mpp_tagring_out_up_10_0;                  
logic          [67:0]  mpp_tagring_out_up_10_1;                  
logic          [67:0]  mpp_tagring_out_up_11_0;                  
logic          [67:0]  mpp_tagring_out_up_11_1;                  
logic          [67:0]  mpp_tagring_out_up_12_0;                  
logic          [67:0]  mpp_tagring_out_up_12_1;                  
logic          [67:0]  mpp_tagring_out_up_13_0;                  
logic          [67:0]  mpp_tagring_out_up_13_1;                  
logic          [67:0]  mpp_tagring_out_up_14_0;                  
logic          [67:0]  mpp_tagring_out_up_14_1;                  
logic          [67:0]  mpp_tagring_out_up_15_0;                  
logic          [67:0]  mpp_tagring_out_up_15_1;                  
logic          [67:0]  mpp_tagring_out_up_1_0;                   
logic          [67:0]  mpp_tagring_out_up_1_1;                   
logic          [67:0]  mpp_tagring_out_up_2_0;                   
logic          [67:0]  mpp_tagring_out_up_2_1;                   
logic          [67:0]  mpp_tagring_out_up_3_0;                   
logic          [67:0]  mpp_tagring_out_up_3_1;                   
logic          [67:0]  mpp_tagring_out_up_4_0;                   
logic          [67:0]  mpp_tagring_out_up_4_1;                   
logic          [67:0]  mpp_tagring_out_up_5_0;                   
logic          [67:0]  mpp_tagring_out_up_5_1;                   
logic          [67:0]  mpp_tagring_out_up_6_0;                   
logic          [67:0]  mpp_tagring_out_up_6_1;                   
logic          [67:0]  mpp_tagring_out_up_7_0;                   
logic          [67:0]  mpp_tagring_out_up_7_1;                   
logic          [67:0]  mpp_tagring_out_up_8_0;                   
logic          [67:0]  mpp_tagring_out_up_8_1;                   
logic          [67:0]  mpp_tagring_out_up_9_0;                   
logic          [67:0]  mpp_tagring_out_up_9_1;                    
// collage-pragma translate_off

import mby_egr_pkg::*; 
import mby_igr_pkg::*; 
import mby_gmm_pkg::*; 
egr_mc_table_if                  egr0_mc_table0();
egr_mc_table_if                  egr0_mc_table1();
egr_ppe_stm_if                   egr0_ppestm();
egr_mc_table_if                  egr1_mc_table0();
egr_mc_table_if                  egr1_mc_table1();
egr_ppe_stm_if                   egr1_ppestm();
egr_cmring_if                    egr_cmring();
//edr logic         fifoEmpty;                      
//edr logic         fifoFilled;                     
logic  [23:0] mgp_dqring_dn_0_0;              
logic  [23:0] mgp_dqring_dn_0_1;              
logic  [23:0] mgp_dqring_dn_1_0;              
logic  [23:0] mgp_dqring_dn_1_1;              
logic  [23:0] mgp_dqring_dn_2_0;              
logic  [23:0] mgp_dqring_dn_2_1;              
logic  [23:0] mgp_dqring_dn_3_0;              
logic  [23:0] mgp_dqring_dn_3_1;              
logic  [23:0] mgp_dqring_dn_4_0;              
logic  [23:0] mgp_dqring_dn_4_1;              
logic  [23:0] mgp_dqring_dn_5_0;              
logic  [23:0] mgp_dqring_dn_5_1;              
logic  [23:0] mgp_dqring_dn_6_0;              
logic  [23:0] mgp_dqring_dn_6_1;              
logic  [23:0] mgp_dqring_dn_7_0;              
logic  [23:0] mgp_dqring_dn_7_1;              
logic  [23:0] mgp_dqring_up_0_0;              
logic  [23:0] mgp_dqring_up_0_1;              
logic  [23:0] mgp_dqring_up_1_0;              
logic  [23:0] mgp_dqring_up_1_1;              
logic  [23:0] mgp_dqring_up_2_0;              
logic  [23:0] mgp_dqring_up_2_1;              
logic  [23:0] mgp_dqring_up_3_0;              
logic  [23:0] mgp_dqring_up_3_1;              
logic  [23:0] mgp_dqring_up_4_0;              
logic  [23:0] mgp_dqring_up_4_1;              
logic  [23:0] mgp_dqring_up_5_0;              
logic  [23:0] mgp_dqring_up_5_1;              
logic  [23:0] mgp_dqring_up_6_0;              
logic  [23:0] mgp_dqring_up_6_1;              
logic  [23:0] mgp_dqring_up_7_0;              
logic  [23:0] mgp_dqring_up_7_1;              
logic  [25:0] mgp_gpolring_dn_0_0;            
logic  [25:0] mgp_gpolring_dn_0_1;            
logic  [25:0] mgp_gpolring_dn_1_0;            
logic  [25:0] mgp_gpolring_dn_1_1;            
logic  [25:0] mgp_gpolring_dn_2_0;            
logic  [25:0] mgp_gpolring_dn_2_1;            
logic  [25:0] mgp_gpolring_dn_3_0;            
logic  [25:0] mgp_gpolring_dn_3_1;            
logic  [25:0] mgp_gpolring_dn_4_0;            
logic  [25:0] mgp_gpolring_dn_4_1;            
logic  [25:0] mgp_gpolring_dn_5_0;            
logic  [25:0] mgp_gpolring_dn_5_1;            
logic  [25:0] mgp_gpolring_dn_6_0;            
logic  [25:0] mgp_gpolring_dn_6_1;            
logic  [25:0] mgp_gpolring_dn_7_0;            
logic  [25:0] mgp_gpolring_dn_7_1;            
logic [106:0] mgp_gpolring_update_dn_0;       
logic [106:0] mgp_gpolring_update_dn_1;       
logic  [68:0] mgp_mctagring_dn_0;             
logic  [68:0] mgp_mctagring_dn_1;             
logic  [68:0] mgp_mctagring_dn_2;             
logic  [68:0] mgp_mctagring_dn_3;             
logic  [68:0] mgp_mctagring_up_0;             
logic  [68:0] mgp_mctagring_up_1;             
logic  [68:0] mgp_mctagring_up_2;             
logic  [68:0] mgp_mctagring_up_3;             
logic  [33:0] mgp_mrpodring_dn;               
logic         mgp_mrpodring_stall_dn;         
logic         mgp_mrpodring_stall_up;         
logic  [33:0] mgp_mrpodring_up;               
logic  [33:0] mgp_podring_dn;                 
logic         mgp_podring_stall_dn;           
logic         mgp_podring_stall_up;           
logic  [33:0] mgp_podring_up;                 
logic  [67:0] mgp_tagring_dn_0_0;             
logic  [67:0] mgp_tagring_dn_0_1;             
logic  [67:0] mgp_tagring_dn_10_0;            
logic  [67:0] mgp_tagring_dn_10_1;            
logic  [67:0] mgp_tagring_dn_11_0;            
logic  [67:0] mgp_tagring_dn_11_1;            
logic  [67:0] mgp_tagring_dn_12_0;            
logic  [67:0] mgp_tagring_dn_12_1;            
logic  [67:0] mgp_tagring_dn_13_0;            
logic  [67:0] mgp_tagring_dn_13_1;            
logic  [67:0] mgp_tagring_dn_14_0;            
logic  [67:0] mgp_tagring_dn_14_1;            
logic  [67:0] mgp_tagring_dn_15_0;            
logic  [67:0] mgp_tagring_dn_15_1;            
logic  [67:0] mgp_tagring_dn_1_0;             
logic  [67:0] mgp_tagring_dn_1_1;             
logic  [67:0] mgp_tagring_dn_2_0;             
logic  [67:0] mgp_tagring_dn_2_1;             
logic  [67:0] mgp_tagring_dn_3_0;             
logic  [67:0] mgp_tagring_dn_3_1;             
logic  [67:0] mgp_tagring_dn_4_0;             
logic  [67:0] mgp_tagring_dn_4_1;             
logic  [67:0] mgp_tagring_dn_5_0;             
logic  [67:0] mgp_tagring_dn_5_1;             
logic  [67:0] mgp_tagring_dn_6_0;             
logic  [67:0] mgp_tagring_dn_6_1;             
logic  [67:0] mgp_tagring_dn_7_0;             
logic  [67:0] mgp_tagring_dn_7_1;             
logic  [67:0] mgp_tagring_dn_8_0;             
logic  [67:0] mgp_tagring_dn_8_1;             
logic  [67:0] mgp_tagring_dn_9_0;             
logic  [67:0] mgp_tagring_dn_9_1;             
logic  [67:0] mgp_tagring_up_0_0;             
logic  [67:0] mgp_tagring_up_0_1;             
logic  [67:0] mgp_tagring_up_10_0;            
logic  [67:0] mgp_tagring_up_10_1;            
logic  [67:0] mgp_tagring_up_11_0;            
logic  [67:0] mgp_tagring_up_11_1;            
logic  [67:0] mgp_tagring_up_12_0;            
logic  [67:0] mgp_tagring_up_12_1;            
logic  [67:0] mgp_tagring_up_13_0;            
logic  [67:0] mgp_tagring_up_13_1;            
logic  [67:0] mgp_tagring_up_14_0;            
logic  [67:0] mgp_tagring_up_14_1;            
logic  [67:0] mgp_tagring_up_15_0;            
logic  [67:0] mgp_tagring_up_15_1;            
logic  [67:0] mgp_tagring_up_1_0;             
logic  [67:0] mgp_tagring_up_1_1;             
logic  [67:0] mgp_tagring_up_2_0;             
logic  [67:0] mgp_tagring_up_2_1;             
logic  [67:0] mgp_tagring_up_3_0;             
logic  [67:0] mgp_tagring_up_3_1;             
logic  [67:0] mgp_tagring_up_4_0;             
logic  [67:0] mgp_tagring_up_4_1;             
logic  [67:0] mgp_tagring_up_5_0;             
logic  [67:0] mgp_tagring_up_5_1;             
logic  [67:0] mgp_tagring_up_6_0;             
logic  [67:0] mgp_tagring_up_6_1;             
logic  [67:0] mgp_tagring_up_7_0;             
logic  [67:0] mgp_tagring_up_7_1;             
logic  [67:0] mgp_tagring_up_8_0;             
logic  [67:0] mgp_tagring_up_8_1;             
logic  [67:0] mgp_tagring_up_9_0;             
logic  [67:0] mgp_tagring_up_9_1;             
//edr logic  [63:0] respData;                       
//edr logic   [7:0] respID;                         
//edr logic         respParity;                     
//edr logic         respValid;                      
rx_ppe_ppe_stm0_if               rxppe0_ppestm0();
rx_ppe_ppe_stm1_if               rxppe0_ppestm1();
rx_ppe_ppe_stm0_if               rxppe1_ppestm0();
rx_ppe_ppe_stm1_if               rxppe1_ppestm1();
ahb_rx_ppe_if ahb0_rxppe();
// Blasted Wires for ahb_rx_ppe_if ppe ahb0_rxppe;
    assign ahb0_rxppe.ahb_sel = ahb0_rxppe_ahb_sel;
    assign ahb0_rxppe.ahb_wr = ahb0_rxppe_ahb_wr;
    assign ahb0_rxppe.ahb_addr = ahb0_rxppe_ahb_addr;
    assign ahb0_rxppe.ahb_wr_data = ahb0_rxppe_ahb_wr_data;
    assign ahb0_rxppe_ahb_rd_data = ahb0_rxppe.ahb_rd_data;
    assign ahb0_rxppe_ahb_rd_ack = ahb0_rxppe.ahb_rd_ack;

ahb_rx_ppe_if ahb0_txppe0();
// Blasted Wires for ahb_rx_ppe_if ppe ahb0_txppe0;
    assign ahb0_txppe0.ahb_sel = ahb0_txppe0_ahb_sel;
    assign ahb0_txppe0.ahb_wr = ahb0_txppe0_ahb_wr;
    assign ahb0_txppe0.ahb_addr = ahb0_txppe0_ahb_addr;
    assign ahb0_txppe0.ahb_wr_data = ahb0_txppe0_ahb_wr_data;
    assign ahb0_txppe0_ahb_rd_data = ahb0_txppe0.ahb_rd_data;
    assign ahb0_txppe0_ahb_rd_ack = ahb0_txppe0.ahb_rd_ack;

ahb_rx_ppe_if ahb0_txppe1();
// Blasted Wires for ahb_rx_ppe_if ppe ahb0_txppe1;
    assign ahb0_txppe1.ahb_sel = ahb0_txppe1_ahb_sel;
    assign ahb0_txppe1.ahb_wr = ahb0_txppe1_ahb_wr;
    assign ahb0_txppe1.ahb_addr = ahb0_txppe1_ahb_addr;
    assign ahb0_txppe1.ahb_wr_data = ahb0_txppe1_ahb_wr_data;
    assign ahb0_txppe1_ahb_rd_data = ahb0_txppe1.ahb_rd_data;
    assign ahb0_txppe1_ahb_rd_ack = ahb0_txppe1.ahb_rd_ack;

ahb_rx_ppe_if ahb1_rxppe();
// Blasted Wires for ahb_rx_ppe_if ppe ahb1_rxppe;
    assign ahb1_rxppe.ahb_sel = ahb1_rxppe_ahb_sel;
    assign ahb1_rxppe.ahb_wr = ahb1_rxppe_ahb_wr;
    assign ahb1_rxppe.ahb_addr = ahb1_rxppe_ahb_addr;
    assign ahb1_rxppe.ahb_wr_data = ahb1_rxppe_ahb_wr_data;
    assign ahb1_rxppe_ahb_rd_data = ahb1_rxppe.ahb_rd_data;
    assign ahb1_rxppe_ahb_rd_ack = ahb1_rxppe.ahb_rd_ack;

ahb_rx_ppe_if ahb1_txppe0();
// Blasted Wires for ahb_rx_ppe_if ppe ahb1_txppe0;
    assign ahb1_txppe0.ahb_sel = ahb1_txppe0_ahb_sel;
    assign ahb1_txppe0.ahb_wr = ahb1_txppe0_ahb_wr;
    assign ahb1_txppe0.ahb_addr = ahb1_txppe0_ahb_addr;
    assign ahb1_txppe0.ahb_wr_data = ahb1_txppe0_ahb_wr_data;
    assign ahb1_txppe0_ahb_rd_data = ahb1_txppe0.ahb_rd_data;
    assign ahb1_txppe0_ahb_rd_ack = ahb1_txppe0.ahb_rd_ack;

ahb_rx_ppe_if ahb1_txppe1();
// Blasted Wires for ahb_rx_ppe_if ppe ahb1_txppe1;
    assign ahb1_txppe1.ahb_sel = ahb1_txppe1_ahb_sel;
    assign ahb1_txppe1.ahb_wr = ahb1_txppe1_ahb_wr;
    assign ahb1_txppe1.ahb_addr = ahb1_txppe1_ahb_addr;
    assign ahb1_txppe1.ahb_wr_data = ahb1_txppe1_ahb_wr_data;
    assign ahb1_txppe1_ahb_rd_data = ahb1_txppe1.ahb_rd_data;
    assign ahb1_txppe1_ahb_rd_ack = ahb1_txppe1.ahb_rd_ack;

egr_ahb_if egr0_ahb();
// Blasted Wires for egr_ahb_if egr egr0_ahb;
    assign egr0_ahb.ahb_req_p = egr0_ahb_ahb_req_p;
    assign egr0_ahb.ahb_addr = egr0_ahb_ahb_addr;
    assign egr0_ahb.ahb_wr = egr0_ahb_ahb_wr;
    assign egr0_ahb.ahb_wr_data = egr0_ahb_ahb_wr_data;
    assign egr0_ahb_ahb_ack_p = egr0_ahb.ahb_ack_p;
    assign egr0_ahb_ahb_rd_data = egr0_ahb.ahb_rd_data;
    assign egr0_ahb.dfxsignal_in = egr0_ahb_dfxsignal_in;
    assign egr0_ahb_dfxsignal_out = egr0_ahb.dfxsignal_out;

egr_ahb_if egr1_ahb();
// Blasted Wires for egr_ahb_if egr egr1_ahb;
    assign egr1_ahb.ahb_req_p = egr1_ahb_ahb_req_p;
    assign egr1_ahb.ahb_addr = egr1_ahb_ahb_addr;
    assign egr1_ahb.ahb_wr = egr1_ahb_ahb_wr;
    assign egr1_ahb.ahb_wr_data = egr1_ahb_ahb_wr_data;
    assign egr1_ahb_ahb_ack_p = egr1_ahb.ahb_ack_p;
    assign egr1_ahb_ahb_rd_data = egr1_ahb.ahb_rd_data;
    assign egr1_ahb.dfxsignal_in = egr1_ahb_dfxsignal_in;
    assign egr1_ahb_dfxsignal_out = egr1_ahb.dfxsignal_out;

glb_rx_ppe_if glb0_rxppe();
// Blasted Wires for glb_rx_ppe_if ppe glb0_rxppe;
    assign glb0_rxppe.glb_sync = glb0_rxppe_glb_sync;
    assign glb0_rxppe_glb_ack = glb0_rxppe.glb_ack;

glb_rx_ppe_if glb0_txppe0();
// Blasted Wires for glb_rx_ppe_if ppe glb0_txppe0;
    assign glb0_txppe0.glb_sync = glb0_txppe0_glb_sync;
    assign glb0_txppe0_glb_ack = glb0_txppe0.glb_ack;

glb_rx_ppe_if glb0_txppe1();
// Blasted Wires for glb_rx_ppe_if ppe glb0_txppe1;
    assign glb0_txppe1.glb_sync = glb0_txppe1_glb_sync;
    assign glb0_txppe1_glb_ack = glb0_txppe1.glb_ack;

glb_rx_ppe_if glb1_rxppe();
// Blasted Wires for glb_rx_ppe_if ppe glb1_rxppe;
    assign glb1_rxppe.glb_sync = glb1_rxppe_glb_sync;
    assign glb1_rxppe_glb_ack = glb1_rxppe.glb_ack;

glb_rx_ppe_if glb1_txppe0();
// Blasted Wires for glb_rx_ppe_if ppe glb1_txppe0;
    assign glb1_txppe0.glb_sync = glb1_txppe0_glb_sync;
    assign glb1_txppe0_glb_ack = glb1_txppe0.glb_ack;

glb_rx_ppe_if glb1_txppe1();
// Blasted Wires for glb_rx_ppe_if ppe glb1_txppe1;
    assign glb1_txppe1.glb_sync = glb1_txppe1_glb_sync;
    assign glb1_txppe1_glb_ack = glb1_txppe1.glb_ack;

egr_epl_if grp_a0();
// Blasted Wires for egr_epl_if egr grp_a0;
    assign grp_a0.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_a0_tx_enable_port_num);
    assign grp_a0.tx_enable = epl_tx_enable_t'(grp_a0_tx_enable);
    assign grp_a0_tx_data_valid = grp_a0.tx_data_valid;
    assign grp_a0_tx_port_num = grp_a0.tx_port_num;
    assign grp_a0_tx_valid_resp = grp_a0.tx_valid_resp;
    assign grp_a0_tx_metadata = grp_a0.tx_metadata;
    assign grp_a0_tx0_data = grp_a0.tx0_data;
    assign grp_a0_tx1_data = grp_a0.tx1_data;
    assign grp_a0_tx2_data = grp_a0.tx2_data;
    assign grp_a0_tx3_data = grp_a0.tx3_data;
    assign grp_a0_tx4_data = grp_a0.tx4_data;
    assign grp_a0_tx5_data = grp_a0.tx5_data;
    assign grp_a0_tx6_data = grp_a0.tx6_data;
    assign grp_a0_tx7_data = grp_a0.tx7_data;
    assign grp_a0.rx_pfc_xoff = grp_a0_rx_pfc_xoff;
    assign grp_a0.rx_pfc_tc_sync = grp_a0_rx_pfc_tc_sync;

egr_epl_if grp_a1();
// Blasted Wires for egr_epl_if egr grp_a1;
    assign grp_a1.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_a1_tx_enable_port_num);
    assign grp_a1.tx_enable = epl_tx_enable_t'(grp_a1_tx_enable);
    assign grp_a1_tx_data_valid = grp_a1.tx_data_valid;
    assign grp_a1_tx_port_num = grp_a1.tx_port_num;
    assign grp_a1_tx_valid_resp = grp_a1.tx_valid_resp;
    assign grp_a1_tx_metadata = grp_a1.tx_metadata;
    assign grp_a1_tx0_data = grp_a1.tx0_data;
    assign grp_a1_tx1_data = grp_a1.tx1_data;
    assign grp_a1_tx2_data = grp_a1.tx2_data;
    assign grp_a1_tx3_data = grp_a1.tx3_data;
    assign grp_a1_tx4_data = grp_a1.tx4_data;
    assign grp_a1_tx5_data = grp_a1.tx5_data;
    assign grp_a1_tx6_data = grp_a1.tx6_data;
    assign grp_a1_tx7_data = grp_a1.tx7_data;
    assign grp_a1.rx_pfc_xoff = grp_a1_rx_pfc_xoff;
    assign grp_a1.rx_pfc_tc_sync = grp_a1_rx_pfc_tc_sync;

egr_epl_if grp_b0();
// Blasted Wires for egr_epl_if egr grp_b0;
    assign grp_b0.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_b0_tx_enable_port_num);
    assign grp_b0.tx_enable = epl_tx_enable_t'(grp_b0_tx_enable);
    assign grp_b0_tx_data_valid = grp_b0.tx_data_valid;
    assign grp_b0_tx_port_num = grp_b0.tx_port_num;
    assign grp_b0_tx_valid_resp = grp_b0.tx_valid_resp;
    assign grp_b0_tx_metadata = grp_b0.tx_metadata;
    assign grp_b0_tx0_data = grp_b0.tx0_data;
    assign grp_b0_tx1_data = grp_b0.tx1_data;
    assign grp_b0_tx2_data = grp_b0.tx2_data;
    assign grp_b0_tx3_data = grp_b0.tx3_data;
    assign grp_b0_tx4_data = grp_b0.tx4_data;
    assign grp_b0_tx5_data = grp_b0.tx5_data;
    assign grp_b0_tx6_data = grp_b0.tx6_data;
    assign grp_b0_tx7_data = grp_b0.tx7_data;
    assign grp_b0.rx_pfc_xoff = grp_b0_rx_pfc_xoff;
    assign grp_b0.rx_pfc_tc_sync = grp_b0_rx_pfc_tc_sync;

egr_epl_if grp_b1();
// Blasted Wires for egr_epl_if egr grp_b1;
    assign grp_b1.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_b1_tx_enable_port_num);
    assign grp_b1.tx_enable = epl_tx_enable_t'(grp_b1_tx_enable);
    assign grp_b1_tx_data_valid = grp_b1.tx_data_valid;
    assign grp_b1_tx_port_num = grp_b1.tx_port_num;
    assign grp_b1_tx_valid_resp = grp_b1.tx_valid_resp;
    assign grp_b1_tx_metadata = grp_b1.tx_metadata;
    assign grp_b1_tx0_data = grp_b1.tx0_data;
    assign grp_b1_tx1_data = grp_b1.tx1_data;
    assign grp_b1_tx2_data = grp_b1.tx2_data;
    assign grp_b1_tx3_data = grp_b1.tx3_data;
    assign grp_b1_tx4_data = grp_b1.tx4_data;
    assign grp_b1_tx5_data = grp_b1.tx5_data;
    assign grp_b1_tx6_data = grp_b1.tx6_data;
    assign grp_b1_tx7_data = grp_b1.tx7_data;
    assign grp_b1.rx_pfc_xoff = grp_b1_rx_pfc_xoff;
    assign grp_b1.rx_pfc_tc_sync = grp_b1_rx_pfc_tc_sync;

egr_epl_if grp_c0();
// Blasted Wires for egr_epl_if egr grp_c0;
    assign grp_c0.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_c0_tx_enable_port_num);
    assign grp_c0.tx_enable = epl_tx_enable_t'(grp_c0_tx_enable);
    assign grp_c0_tx_data_valid = grp_c0.tx_data_valid;
    assign grp_c0_tx_port_num = grp_c0.tx_port_num;
    assign grp_c0_tx_valid_resp = grp_c0.tx_valid_resp;
    assign grp_c0_tx_metadata = grp_c0.tx_metadata;
    assign grp_c0_tx0_data = grp_c0.tx0_data;
    assign grp_c0_tx1_data = grp_c0.tx1_data;
    assign grp_c0_tx2_data = grp_c0.tx2_data;
    assign grp_c0_tx3_data = grp_c0.tx3_data;
    assign grp_c0_tx4_data = grp_c0.tx4_data;
    assign grp_c0_tx5_data = grp_c0.tx5_data;
    assign grp_c0_tx6_data = grp_c0.tx6_data;
    assign grp_c0_tx7_data = grp_c0.tx7_data;
    assign grp_c0.rx_pfc_xoff = grp_c0_rx_pfc_xoff;
    assign grp_c0.rx_pfc_tc_sync = grp_c0_rx_pfc_tc_sync;

egr_epl_if grp_c1();
// Blasted Wires for egr_epl_if egr grp_c1;
    assign grp_c1.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_c1_tx_enable_port_num);
    assign grp_c1.tx_enable = epl_tx_enable_t'(grp_c1_tx_enable);
    assign grp_c1_tx_data_valid = grp_c1.tx_data_valid;
    assign grp_c1_tx_port_num = grp_c1.tx_port_num;
    assign grp_c1_tx_valid_resp = grp_c1.tx_valid_resp;
    assign grp_c1_tx_metadata = grp_c1.tx_metadata;
    assign grp_c1_tx0_data = grp_c1.tx0_data;
    assign grp_c1_tx1_data = grp_c1.tx1_data;
    assign grp_c1_tx2_data = grp_c1.tx2_data;
    assign grp_c1_tx3_data = grp_c1.tx3_data;
    assign grp_c1_tx4_data = grp_c1.tx4_data;
    assign grp_c1_tx5_data = grp_c1.tx5_data;
    assign grp_c1_tx6_data = grp_c1.tx6_data;
    assign grp_c1_tx7_data = grp_c1.tx7_data;
    assign grp_c1.rx_pfc_xoff = grp_c1_rx_pfc_xoff;
    assign grp_c1.rx_pfc_tc_sync = grp_c1_rx_pfc_tc_sync;

egr_epl_if grp_d0();
// Blasted Wires for egr_epl_if egr grp_d0;
    assign grp_d0.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_d0_tx_enable_port_num);
    assign grp_d0.tx_enable = epl_tx_enable_t'(grp_d0_tx_enable);
    assign grp_d0_tx_data_valid = grp_d0.tx_data_valid;
    assign grp_d0_tx_port_num = grp_d0.tx_port_num;
    assign grp_d0_tx_valid_resp = grp_d0.tx_valid_resp;
    assign grp_d0_tx_metadata = grp_d0.tx_metadata;
    assign grp_d0_tx0_data = grp_d0.tx0_data;
    assign grp_d0_tx1_data = grp_d0.tx1_data;
    assign grp_d0_tx2_data = grp_d0.tx2_data;
    assign grp_d0_tx3_data = grp_d0.tx3_data;
    assign grp_d0_tx4_data = grp_d0.tx4_data;
    assign grp_d0_tx5_data = grp_d0.tx5_data;
    assign grp_d0_tx6_data = grp_d0.tx6_data;
    assign grp_d0_tx7_data = grp_d0.tx7_data;
    assign grp_d0.rx_pfc_xoff = grp_d0_rx_pfc_xoff;
    assign grp_d0.rx_pfc_tc_sync = grp_d0_rx_pfc_tc_sync;

egr_epl_if grp_d1();
// Blasted Wires for egr_epl_if egr grp_d1;
    assign grp_d1.tx_enable_port_num = epl_tx_enable_port_num_t'(grp_d1_tx_enable_port_num);
    assign grp_d1.tx_enable = epl_tx_enable_t'(grp_d1_tx_enable);
    assign grp_d1_tx_data_valid = grp_d1.tx_data_valid;
    assign grp_d1_tx_port_num = grp_d1.tx_port_num;
    assign grp_d1_tx_valid_resp = grp_d1.tx_valid_resp;
    assign grp_d1_tx_metadata = grp_d1.tx_metadata;
    assign grp_d1_tx0_data = grp_d1.tx0_data;
    assign grp_d1_tx1_data = grp_d1.tx1_data;
    assign grp_d1_tx2_data = grp_d1.tx2_data;
    assign grp_d1_tx3_data = grp_d1.tx3_data;
    assign grp_d1_tx4_data = grp_d1.tx4_data;
    assign grp_d1_tx5_data = grp_d1.tx5_data;
    assign grp_d1_tx6_data = grp_d1.tx6_data;
    assign grp_d1_tx7_data = grp_d1.tx7_data;
    assign grp_d1.rx_pfc_xoff = grp_d1_rx_pfc_xoff;
    assign grp_d1.rx_pfc_tc_sync = grp_d1_rx_pfc_tc_sync;

mim_rd_if mim0_rd0();
// Blasted Wires for mim_rd_if request mim0_rd0;
    assign mim0_rd0_mim_rreq_valid = mim0_rd0.mim_rreq_valid;
    assign mim0_rd0_mim_seg_ptr = mim0_rd0.mim_seg_ptr;
    assign mim0_rd0_mim_sema = mim0_rd0.mim_sema;
    assign mim0_rd0_mim_wd_sel = mim0_rd0.mim_wd_sel;
    assign mim0_rd0_mim_req_id = mim0_rd0.mim_req_id;
    assign mim0_rd0.mim_rreq_credits = mim0_rd0_mim_rreq_credits;
    assign mim0_rd0.mim_rrsp_valid = mim0_rd0_mim_rrsp_valid;
    assign mim0_rd0.mim_rrsp_dest_block = mim0_rd0_mim_rrsp_dest_block;
    assign mim0_rd0.mim_rrsp_req_id = mim0_rd0_mim_rrsp_req_id;
    assign mim0_rd0.mim_rd_data = mim0_rd0_mim_rd_data;

mim_rd_if mim0_rd1();
// Blasted Wires for mim_rd_if request mim0_rd1;
    assign mim0_rd1_mim_rreq_valid = mim0_rd1.mim_rreq_valid;
    assign mim0_rd1_mim_seg_ptr = mim0_rd1.mim_seg_ptr;
    assign mim0_rd1_mim_sema = mim0_rd1.mim_sema;
    assign mim0_rd1_mim_wd_sel = mim0_rd1.mim_wd_sel;
    assign mim0_rd1_mim_req_id = mim0_rd1.mim_req_id;
    assign mim0_rd1.mim_rreq_credits = mim0_rd1_mim_rreq_credits;
    assign mim0_rd1.mim_rrsp_valid = mim0_rd1_mim_rrsp_valid;
    assign mim0_rd1.mim_rrsp_dest_block = mim0_rd1_mim_rrsp_dest_block;
    assign mim0_rd1.mim_rrsp_req_id = mim0_rd1_mim_rrsp_req_id;
    assign mim0_rd1.mim_rd_data = mim0_rd1_mim_rd_data;

mim_rd_if mim0_rd2();
// Blasted Wires for mim_rd_if request mim0_rd2;
    assign mim0_rd2_mim_rreq_valid = mim0_rd2.mim_rreq_valid;
    assign mim0_rd2_mim_seg_ptr = mim0_rd2.mim_seg_ptr;
    assign mim0_rd2_mim_sema = mim0_rd2.mim_sema;
    assign mim0_rd2_mim_wd_sel = mim0_rd2.mim_wd_sel;
    assign mim0_rd2_mim_req_id = mim0_rd2.mim_req_id;
    assign mim0_rd2.mim_rreq_credits = mim0_rd2_mim_rreq_credits;
    assign mim0_rd2.mim_rrsp_valid = mim0_rd2_mim_rrsp_valid;
    assign mim0_rd2.mim_rrsp_dest_block = mim0_rd2_mim_rrsp_dest_block;
    assign mim0_rd2.mim_rrsp_req_id = mim0_rd2_mim_rrsp_req_id;
    assign mim0_rd2.mim_rd_data = mim0_rd2_mim_rd_data;

mim_wr_if mim0_wr0();
// Blasted Wires for mim_wr_if request mim0_wr0;
    assign mim0_wr0_mim_wreq_valid = mim0_wr0.mim_wreq_valid;
    assign mim0_wr0_mim_wr_seg_ptr = mim0_wr0.mim_wr_seg_ptr;
    assign mim0_wr0_mim_wr_sema = mim0_wr0.mim_wr_sema;
    assign mim0_wr0_mim_wr_wd_sel = mim0_wr0.mim_wr_wd_sel;
    assign mim0_wr0_mim_wreq_id = mim0_wr0.mim_wreq_id;
    assign mim0_wr0_mim_wr_data = mim0_wr0.mim_wr_data;
    assign mim0_wr0.mim_wreq_credits = mim0_wr0_mim_wreq_credits;

mim_wr_if mim0_wr1();
// Blasted Wires for mim_wr_if request mim0_wr1;
    assign mim0_wr1_mim_wreq_valid = mim0_wr1.mim_wreq_valid;
    assign mim0_wr1_mim_wr_seg_ptr = mim0_wr1.mim_wr_seg_ptr;
    assign mim0_wr1_mim_wr_sema = mim0_wr1.mim_wr_sema;
    assign mim0_wr1_mim_wr_wd_sel = mim0_wr1.mim_wr_wd_sel;
    assign mim0_wr1_mim_wreq_id = mim0_wr1.mim_wreq_id;
    assign mim0_wr1_mim_wr_data = mim0_wr1.mim_wr_data;
    assign mim0_wr1.mim_wreq_credits = mim0_wr1_mim_wreq_credits;

mim_wr_if mim0_wr2();
// Blasted Wires for mim_wr_if request mim0_wr2;
    assign mim0_wr2_mim_wreq_valid = mim0_wr2.mim_wreq_valid;
    assign mim0_wr2_mim_wr_seg_ptr = mim0_wr2.mim_wr_seg_ptr;
    assign mim0_wr2_mim_wr_sema = mim0_wr2.mim_wr_sema;
    assign mim0_wr2_mim_wr_wd_sel = mim0_wr2.mim_wr_wd_sel;
    assign mim0_wr2_mim_wreq_id = mim0_wr2.mim_wreq_id;
    assign mim0_wr2_mim_wr_data = mim0_wr2.mim_wr_data;
    assign mim0_wr2.mim_wreq_credits = mim0_wr2_mim_wreq_credits;

mim_rd_if mim1_rd0();
// Blasted Wires for mim_rd_if request mim1_rd0;
    assign mim1_rd0_mim_rreq_valid = mim1_rd0.mim_rreq_valid;
    assign mim1_rd0_mim_seg_ptr = mim1_rd0.mim_seg_ptr;
    assign mim1_rd0_mim_sema = mim1_rd0.mim_sema;
    assign mim1_rd0_mim_wd_sel = mim1_rd0.mim_wd_sel;
    assign mim1_rd0_mim_req_id = mim1_rd0.mim_req_id;
    assign mim1_rd0.mim_rreq_credits = mim1_rd0_mim_rreq_credits;
    assign mim1_rd0.mim_rrsp_valid = mim1_rd0_mim_rrsp_valid;
    assign mim1_rd0.mim_rrsp_dest_block = mim1_rd0_mim_rrsp_dest_block;
    assign mim1_rd0.mim_rrsp_req_id = mim1_rd0_mim_rrsp_req_id;
    assign mim1_rd0.mim_rd_data = mim1_rd0_mim_rd_data;

mim_rd_if mim1_rd1();
// Blasted Wires for mim_rd_if request mim1_rd1;
    assign mim1_rd1_mim_rreq_valid = mim1_rd1.mim_rreq_valid;
    assign mim1_rd1_mim_seg_ptr = mim1_rd1.mim_seg_ptr;
    assign mim1_rd1_mim_sema = mim1_rd1.mim_sema;
    assign mim1_rd1_mim_wd_sel = mim1_rd1.mim_wd_sel;
    assign mim1_rd1_mim_req_id = mim1_rd1.mim_req_id;
    assign mim1_rd1.mim_rreq_credits = mim1_rd1_mim_rreq_credits;
    assign mim1_rd1.mim_rrsp_valid = mim1_rd1_mim_rrsp_valid;
    assign mim1_rd1.mim_rrsp_dest_block = mim1_rd1_mim_rrsp_dest_block;
    assign mim1_rd1.mim_rrsp_req_id = mim1_rd1_mim_rrsp_req_id;
    assign mim1_rd1.mim_rd_data = mim1_rd1_mim_rd_data;

mim_rd_if mim1_rd2();
// Blasted Wires for mim_rd_if request mim1_rd2;
    assign mim1_rd2_mim_rreq_valid = mim1_rd2.mim_rreq_valid;
    assign mim1_rd2_mim_seg_ptr = mim1_rd2.mim_seg_ptr;
    assign mim1_rd2_mim_sema = mim1_rd2.mim_sema;
    assign mim1_rd2_mim_wd_sel = mim1_rd2.mim_wd_sel;
    assign mim1_rd2_mim_req_id = mim1_rd2.mim_req_id;
    assign mim1_rd2.mim_rreq_credits = mim1_rd2_mim_rreq_credits;
    assign mim1_rd2.mim_rrsp_valid = mim1_rd2_mim_rrsp_valid;
    assign mim1_rd2.mim_rrsp_dest_block = mim1_rd2_mim_rrsp_dest_block;
    assign mim1_rd2.mim_rrsp_req_id = mim1_rd2_mim_rrsp_req_id;
    assign mim1_rd2.mim_rd_data = mim1_rd2_mim_rd_data;

mim_wr_if mim1_wr0();
// Blasted Wires for mim_wr_if request mim1_wr0;
    assign mim1_wr0_mim_wreq_valid = mim1_wr0.mim_wreq_valid;
    assign mim1_wr0_mim_wr_seg_ptr = mim1_wr0.mim_wr_seg_ptr;
    assign mim1_wr0_mim_wr_sema = mim1_wr0.mim_wr_sema;
    assign mim1_wr0_mim_wr_wd_sel = mim1_wr0.mim_wr_wd_sel;
    assign mim1_wr0_mim_wreq_id = mim1_wr0.mim_wreq_id;
    assign mim1_wr0_mim_wr_data = mim1_wr0.mim_wr_data;
    assign mim1_wr0.mim_wreq_credits = mim1_wr0_mim_wreq_credits;

mim_wr_if mim1_wr1();
// Blasted Wires for mim_wr_if request mim1_wr1;
    assign mim1_wr1_mim_wreq_valid = mim1_wr1.mim_wreq_valid;
    assign mim1_wr1_mim_wr_seg_ptr = mim1_wr1.mim_wr_seg_ptr;
    assign mim1_wr1_mim_wr_sema = mim1_wr1.mim_wr_sema;
    assign mim1_wr1_mim_wr_wd_sel = mim1_wr1.mim_wr_wd_sel;
    assign mim1_wr1_mim_wreq_id = mim1_wr1.mim_wreq_id;
    assign mim1_wr1_mim_wr_data = mim1_wr1.mim_wr_data;
    assign mim1_wr1.mim_wreq_credits = mim1_wr1_mim_wreq_credits;

mim_wr_if mim1_wr2();
// Blasted Wires for mim_wr_if request mim1_wr2;
    assign mim1_wr2_mim_wreq_valid = mim1_wr2.mim_wreq_valid;
    assign mim1_wr2_mim_wr_seg_ptr = mim1_wr2.mim_wr_seg_ptr;
    assign mim1_wr2_mim_wr_sema = mim1_wr2.mim_wr_sema;
    assign mim1_wr2_mim_wr_wd_sel = mim1_wr2.mim_wr_wd_sel;
    assign mim1_wr2_mim_wreq_id = mim1_wr2.mim_wreq_id;
    assign mim1_wr2_mim_wr_data = mim1_wr2.mim_wr_data;
    assign mim1_wr2.mim_wreq_credits = mim1_wr2_mim_wreq_credits;

mim_rd_if mim2_rd0();
// Blasted Wires for mim_rd_if request mim2_rd0;
    assign mim2_rd0_mim_rreq_valid = mim2_rd0.mim_rreq_valid;
    assign mim2_rd0_mim_seg_ptr = mim2_rd0.mim_seg_ptr;
    assign mim2_rd0_mim_sema = mim2_rd0.mim_sema;
    assign mim2_rd0_mim_wd_sel = mim2_rd0.mim_wd_sel;
    assign mim2_rd0_mim_req_id = mim2_rd0.mim_req_id;
    assign mim2_rd0.mim_rreq_credits = mim2_rd0_mim_rreq_credits;
    assign mim2_rd0.mim_rrsp_valid = mim2_rd0_mim_rrsp_valid;
    assign mim2_rd0.mim_rrsp_dest_block = mim2_rd0_mim_rrsp_dest_block;
    assign mim2_rd0.mim_rrsp_req_id = mim2_rd0_mim_rrsp_req_id;
    assign mim2_rd0.mim_rd_data = mim2_rd0_mim_rd_data;

mim_rd_if mim2_rd1();
// Blasted Wires for mim_rd_if request mim2_rd1;
    assign mim2_rd1_mim_rreq_valid = mim2_rd1.mim_rreq_valid;
    assign mim2_rd1_mim_seg_ptr = mim2_rd1.mim_seg_ptr;
    assign mim2_rd1_mim_sema = mim2_rd1.mim_sema;
    assign mim2_rd1_mim_wd_sel = mim2_rd1.mim_wd_sel;
    assign mim2_rd1_mim_req_id = mim2_rd1.mim_req_id;
    assign mim2_rd1.mim_rreq_credits = mim2_rd1_mim_rreq_credits;
    assign mim2_rd1.mim_rrsp_valid = mim2_rd1_mim_rrsp_valid;
    assign mim2_rd1.mim_rrsp_dest_block = mim2_rd1_mim_rrsp_dest_block;
    assign mim2_rd1.mim_rrsp_req_id = mim2_rd1_mim_rrsp_req_id;
    assign mim2_rd1.mim_rd_data = mim2_rd1_mim_rd_data;

mim_rd_if mim2_rd2();
// Blasted Wires for mim_rd_if request mim2_rd2;
    assign mim2_rd2_mim_rreq_valid = mim2_rd2.mim_rreq_valid;
    assign mim2_rd2_mim_seg_ptr = mim2_rd2.mim_seg_ptr;
    assign mim2_rd2_mim_sema = mim2_rd2.mim_sema;
    assign mim2_rd2_mim_wd_sel = mim2_rd2.mim_wd_sel;
    assign mim2_rd2_mim_req_id = mim2_rd2.mim_req_id;
    assign mim2_rd2.mim_rreq_credits = mim2_rd2_mim_rreq_credits;
    assign mim2_rd2.mim_rrsp_valid = mim2_rd2_mim_rrsp_valid;
    assign mim2_rd2.mim_rrsp_dest_block = mim2_rd2_mim_rrsp_dest_block;
    assign mim2_rd2.mim_rrsp_req_id = mim2_rd2_mim_rrsp_req_id;
    assign mim2_rd2.mim_rd_data = mim2_rd2_mim_rd_data;

mim_wr_if mim2_wr0();
// Blasted Wires for mim_wr_if request mim2_wr0;
    assign mim2_wr0_mim_wreq_valid = mim2_wr0.mim_wreq_valid;
    assign mim2_wr0_mim_wr_seg_ptr = mim2_wr0.mim_wr_seg_ptr;
    assign mim2_wr0_mim_wr_sema = mim2_wr0.mim_wr_sema;
    assign mim2_wr0_mim_wr_wd_sel = mim2_wr0.mim_wr_wd_sel;
    assign mim2_wr0_mim_wreq_id = mim2_wr0.mim_wreq_id;
    assign mim2_wr0_mim_wr_data = mim2_wr0.mim_wr_data;
    assign mim2_wr0.mim_wreq_credits = mim2_wr0_mim_wreq_credits;

mim_wr_if mim2_wr1();
// Blasted Wires for mim_wr_if request mim2_wr1;
    assign mim2_wr1_mim_wreq_valid = mim2_wr1.mim_wreq_valid;
    assign mim2_wr1_mim_wr_seg_ptr = mim2_wr1.mim_wr_seg_ptr;
    assign mim2_wr1_mim_wr_sema = mim2_wr1.mim_wr_sema;
    assign mim2_wr1_mim_wr_wd_sel = mim2_wr1.mim_wr_wd_sel;
    assign mim2_wr1_mim_wreq_id = mim2_wr1.mim_wreq_id;
    assign mim2_wr1_mim_wr_data = mim2_wr1.mim_wr_data;
    assign mim2_wr1.mim_wreq_credits = mim2_wr1_mim_wreq_credits;

mim_wr_if mim2_wr2();
// Blasted Wires for mim_wr_if request mim2_wr2;
    assign mim2_wr2_mim_wreq_valid = mim2_wr2.mim_wreq_valid;
    assign mim2_wr2_mim_wr_seg_ptr = mim2_wr2.mim_wr_seg_ptr;
    assign mim2_wr2_mim_wr_sema = mim2_wr2.mim_wr_sema;
    assign mim2_wr2_mim_wr_wd_sel = mim2_wr2.mim_wr_wd_sel;
    assign mim2_wr2_mim_wreq_id = mim2_wr2.mim_wreq_id;
    assign mim2_wr2_mim_wr_data = mim2_wr2.mim_wr_data;
    assign mim2_wr2.mim_wreq_credits = mim2_wr2_mim_wreq_credits;

mim_rd_if mim3_rd0();
// Blasted Wires for mim_rd_if request mim3_rd0;
    assign mim3_rd0_mim_rreq_valid = mim3_rd0.mim_rreq_valid;
    assign mim3_rd0_mim_seg_ptr = mim3_rd0.mim_seg_ptr;
    assign mim3_rd0_mim_sema = mim3_rd0.mim_sema;
    assign mim3_rd0_mim_wd_sel = mim3_rd0.mim_wd_sel;
    assign mim3_rd0_mim_req_id = mim3_rd0.mim_req_id;
    assign mim3_rd0.mim_rreq_credits = mim3_rd0_mim_rreq_credits;
    assign mim3_rd0.mim_rrsp_valid = mim3_rd0_mim_rrsp_valid;
    assign mim3_rd0.mim_rrsp_dest_block = mim3_rd0_mim_rrsp_dest_block;
    assign mim3_rd0.mim_rrsp_req_id = mim3_rd0_mim_rrsp_req_id;
    assign mim3_rd0.mim_rd_data = mim3_rd0_mim_rd_data;

mim_rd_if mim3_rd1();
// Blasted Wires for mim_rd_if request mim3_rd1;
    assign mim3_rd1_mim_rreq_valid = mim3_rd1.mim_rreq_valid;
    assign mim3_rd1_mim_seg_ptr = mim3_rd1.mim_seg_ptr;
    assign mim3_rd1_mim_sema = mim3_rd1.mim_sema;
    assign mim3_rd1_mim_wd_sel = mim3_rd1.mim_wd_sel;
    assign mim3_rd1_mim_req_id = mim3_rd1.mim_req_id;
    assign mim3_rd1.mim_rreq_credits = mim3_rd1_mim_rreq_credits;
    assign mim3_rd1.mim_rrsp_valid = mim3_rd1_mim_rrsp_valid;
    assign mim3_rd1.mim_rrsp_dest_block = mim3_rd1_mim_rrsp_dest_block;
    assign mim3_rd1.mim_rrsp_req_id = mim3_rd1_mim_rrsp_req_id;
    assign mim3_rd1.mim_rd_data = mim3_rd1_mim_rd_data;

mim_rd_if mim3_rd2();
// Blasted Wires for mim_rd_if request mim3_rd2;
    assign mim3_rd2_mim_rreq_valid = mim3_rd2.mim_rreq_valid;
    assign mim3_rd2_mim_seg_ptr = mim3_rd2.mim_seg_ptr;
    assign mim3_rd2_mim_sema = mim3_rd2.mim_sema;
    assign mim3_rd2_mim_wd_sel = mim3_rd2.mim_wd_sel;
    assign mim3_rd2_mim_req_id = mim3_rd2.mim_req_id;
    assign mim3_rd2.mim_rreq_credits = mim3_rd2_mim_rreq_credits;
    assign mim3_rd2.mim_rrsp_valid = mim3_rd2_mim_rrsp_valid;
    assign mim3_rd2.mim_rrsp_dest_block = mim3_rd2_mim_rrsp_dest_block;
    assign mim3_rd2.mim_rrsp_req_id = mim3_rd2_mim_rrsp_req_id;
    assign mim3_rd2.mim_rd_data = mim3_rd2_mim_rd_data;

mim_wr_if mim3_wr0();
// Blasted Wires for mim_wr_if request mim3_wr0;
    assign mim3_wr0_mim_wreq_valid = mim3_wr0.mim_wreq_valid;
    assign mim3_wr0_mim_wr_seg_ptr = mim3_wr0.mim_wr_seg_ptr;
    assign mim3_wr0_mim_wr_sema = mim3_wr0.mim_wr_sema;
    assign mim3_wr0_mim_wr_wd_sel = mim3_wr0.mim_wr_wd_sel;
    assign mim3_wr0_mim_wreq_id = mim3_wr0.mim_wreq_id;
    assign mim3_wr0_mim_wr_data = mim3_wr0.mim_wr_data;
    assign mim3_wr0.mim_wreq_credits = mim3_wr0_mim_wreq_credits;

mim_wr_if mim3_wr1();
// Blasted Wires for mim_wr_if request mim3_wr1;
    assign mim3_wr1_mim_wreq_valid = mim3_wr1.mim_wreq_valid;
    assign mim3_wr1_mim_wr_seg_ptr = mim3_wr1.mim_wr_seg_ptr;
    assign mim3_wr1_mim_wr_sema = mim3_wr1.mim_wr_sema;
    assign mim3_wr1_mim_wr_wd_sel = mim3_wr1.mim_wr_wd_sel;
    assign mim3_wr1_mim_wreq_id = mim3_wr1.mim_wreq_id;
    assign mim3_wr1_mim_wr_data = mim3_wr1.mim_wr_data;
    assign mim3_wr1.mim_wreq_credits = mim3_wr1_mim_wreq_credits;

mim_wr_if mim3_wr2();
// Blasted Wires for mim_wr_if request mim3_wr2;
    assign mim3_wr2_mim_wreq_valid = mim3_wr2.mim_wreq_valid;
    assign mim3_wr2_mim_wr_seg_ptr = mim3_wr2.mim_wr_seg_ptr;
    assign mim3_wr2_mim_wr_sema = mim3_wr2.mim_wr_sema;
    assign mim3_wr2_mim_wr_wd_sel = mim3_wr2.mim_wr_wd_sel;
    assign mim3_wr2_mim_wreq_id = mim3_wr2.mim_wreq_id;
    assign mim3_wr2_mim_wr_data = mim3_wr2.mim_wr_data;
    assign mim3_wr2.mim_wreq_credits = mim3_wr2_mim_wreq_credits;



// module mgp0    from mby_mgp using mgp.map 0
mby_mgp    mgp0(
/* input  logic                     */ .arst_n                     (arst_n),                                     //Asynchronous negedge reset     
/* input  logic                     */ .cclk                       (cclk),                                       
/* input  logic              [23:0] */ .dqring_in_dn_0_0           (mpp_dqring_in_0_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_0_1           (mpp_dqring_in_0_1),                          
/* input  logic              [23:0] */ .dqring_in_dn_1_0           (mpp_dqring_in_1_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_1_1           (mpp_dqring_in_1_1),                          
/* input  logic              [23:0] */ .dqring_in_dn_2_0           (mpp_dqring_in_2_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_2_1           (mpp_dqring_in_2_1),                          
/* input  logic              [23:0] */ .dqring_in_dn_3_0           (mpp_dqring_in_3_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_3_1           (mpp_dqring_in_3_1),                          
/* input  logic              [23:0] */ .dqring_in_dn_4_0           (mpp_dqring_in_4_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_4_1           (mpp_dqring_in_4_1),                          
/* input  logic              [23:0] */ .dqring_in_dn_5_0           (mpp_dqring_in_5_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_5_1           (mpp_dqring_in_5_1),                          
/* input  logic              [23:0] */ .dqring_in_dn_6_0           (mpp_dqring_in_6_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_6_1           (mpp_dqring_in_6_1),                          
/* input  logic              [23:0] */ .dqring_in_dn_7_0           (mpp_dqring_in_7_0),                          
/* input  logic              [23:0] */ .dqring_in_dn_7_1           (mpp_dqring_in_7_1),                          
/* input  logic              [23:0] */ .dqring_in_up_0_0           (mgp_dqring_up_0_0),                          
/* input  logic              [23:0] */ .dqring_in_up_0_1           (mgp_dqring_up_0_1),                          
/* input  logic              [23:0] */ .dqring_in_up_1_0           (mgp_dqring_up_1_0),                          
/* input  logic              [23:0] */ .dqring_in_up_1_1           (mgp_dqring_up_1_1),                          
/* input  logic              [23:0] */ .dqring_in_up_2_0           (mgp_dqring_up_2_0),                          
/* input  logic              [23:0] */ .dqring_in_up_2_1           (mgp_dqring_up_2_1),                          
/* input  logic              [23:0] */ .dqring_in_up_3_0           (mgp_dqring_up_3_0),                          
/* input  logic              [23:0] */ .dqring_in_up_3_1           (mgp_dqring_up_3_1),                          
/* input  logic              [23:0] */ .dqring_in_up_4_0           (mgp_dqring_up_4_0),                          
/* input  logic              [23:0] */ .dqring_in_up_4_1           (mgp_dqring_up_4_1),                          
/* input  logic              [23:0] */ .dqring_in_up_5_0           (mgp_dqring_up_5_0),                          
/* input  logic              [23:0] */ .dqring_in_up_5_1           (mgp_dqring_up_5_1),                          
/* input  logic              [23:0] */ .dqring_in_up_6_0           (mgp_dqring_up_6_0),                          
/* input  logic              [23:0] */ .dqring_in_up_6_1           (mgp_dqring_up_6_1),                          
/* input  logic              [23:0] */ .dqring_in_up_7_0           (mgp_dqring_up_7_0),                          
/* input  logic              [23:0] */ .dqring_in_up_7_1           (mgp_dqring_up_7_1),                          
/* input  logic              [25:0] */ .gpolring_in_dn_0_0         (mpp_gpolring_in_0_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_0_1         (mpp_gpolring_in_0_1),                        
/* input  logic              [25:0] */ .gpolring_in_dn_1_0         (mpp_gpolring_in_1_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_1_1         (mpp_gpolring_in_1_1),                        
/* input  logic              [25:0] */ .gpolring_in_dn_2_0         (mpp_gpolring_in_2_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_2_1         (mpp_gpolring_in_2_1),                        
/* input  logic              [25:0] */ .gpolring_in_dn_3_0         (mpp_gpolring_in_3_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_3_1         (mpp_gpolring_in_3_1),                        
/* input  logic              [25:0] */ .gpolring_in_dn_4_0         (mpp_gpolring_in_4_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_4_1         (mpp_gpolring_in_4_1),                        
/* input  logic              [25:0] */ .gpolring_in_dn_5_0         (mpp_gpolring_in_5_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_5_1         (mpp_gpolring_in_5_1),                        
/* input  logic              [25:0] */ .gpolring_in_dn_6_0         (mpp_gpolring_in_6_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_6_1         (mpp_gpolring_in_6_1),                        
/* input  logic              [25:0] */ .gpolring_in_dn_7_0         (mpp_gpolring_in_7_0),                        
/* input  logic              [25:0] */ .gpolring_in_dn_7_1         (mpp_gpolring_in_7_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_0_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_0_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_1_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_1_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_2_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_2_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_3_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_3_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_4_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_4_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_5_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_5_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_6_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_6_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_7_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_7_1         ({26'b0}),                                    
/* input  logic             [106:0] */ .gpolring_update_in_dn_0    (mpp_gpolring_update_in_0),                   
/* input  logic             [106:0] */ .gpolring_update_in_dn_1    (mpp_gpolring_update_in_1),                   
/* input  logic             [106:0] */ .gpolring_update_in_up_0    ({107'b0}),                                   
/* input  logic             [106:0] */ .gpolring_update_in_up_1    ({107'b0}),                                   
/* input  logic         [0:7][63:0] */ .grp_a_rx_data              ({grp_a0_rx0_data[63:0], grp_a0_rx1_data[63:0], grp_a0_rx2_data[63:0], grp_a0_rx3_data[63:0], grp_a0_rx4_data[63:0], grp_a0_rx5_data[63:0], grp_a0_rx6_data[63:0], grp_a0_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_a_rx_data_valid        (grp_a0_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_a_rx_metadata          ({grp_a0_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_a_rx_port_num          (grp_a0_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_a_rx_time_stamp        ({grp_a0_rx_time_stamp[39:0]}),               
/* input  logic         [0:7][63:0] */ .grp_b_rx_data              ({grp_b0_rx0_data[63:0], grp_b0_rx1_data[63:0], grp_b0_rx2_data[63:0], grp_b0_rx3_data[63:0], grp_b0_rx4_data[63:0], grp_b0_rx5_data[63:0], grp_b0_rx6_data[63:0], grp_b0_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_b_rx_data_valid        (grp_b0_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_b_rx_metadata          ({grp_b0_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_b_rx_port_num          (grp_b0_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_b_rx_time_stamp        ({grp_b0_rx_time_stamp[39:0]}),               
/* input  logic         [0:7][63:0] */ .grp_c_rx_data              ({grp_c0_rx0_data[63:0], grp_c0_rx1_data[63:0], grp_c0_rx2_data[63:0], grp_c0_rx3_data[63:0], grp_c0_rx4_data[63:0], grp_c0_rx5_data[63:0], grp_c0_rx6_data[63:0], grp_c0_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_c_rx_data_valid        (grp_c0_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_c_rx_metadata          ({grp_c0_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_c_rx_port_num          (grp_c0_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_c_rx_time_stamp        ({grp_c0_rx_time_stamp[39:0]}),               
/* input  logic         [0:7][63:0] */ .grp_d_rx_data              ({grp_d0_rx0_data[63:0], grp_d0_rx1_data[63:0], grp_d0_rx2_data[63:0], grp_d0_rx3_data[63:0], grp_d0_rx4_data[63:0], grp_d0_rx5_data[63:0], grp_d0_rx6_data[63:0], grp_d0_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_d_rx_data_valid        (grp_d0_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_d_rx_metadata          ({grp_d0_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_d_rx_port_num          (grp_d0_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_d_rx_time_stamp        ({grp_d0_rx_time_stamp[39:0]}),               
/* input  logic              [19:0] */ .igr_vp_cpp_rx_metadata     (igr0_vp_cpp_rx_metadata),                    
/* input  logic               [7:0] */ .igr_vp_rx_data_valid       (igr0_vp_rx_data_valid),                      
/* input  logic         [0:7][71:0] */ .igr_vp_rx_data_w_ecc       ({igr0_vp_rx0_data_w_ecc[71:0], igr0_vp_rx1_data_w_ecc[71:0], igr0_vp_rx2_data_w_ecc[71:0], igr0_vp_rx3_data_w_ecc[71:0], igr0_vp_rx4_data_w_ecc[71:0], igr0_vp_rx5_data_w_ecc[71:0], igr0_vp_rx6_data_w_ecc[71:0], igr0_vp_rx7_data_w_ecc[71:0]}), 
/* input  logic               [7:0] */ .igr_vp_rx_ecc              (igr0_vp_rx_ecc),                             
/* input  logic               [2:0] */ .igr_vp_rx_flow_control_tc  (igr0_vp_rx_flow_control_tc),                 
/* input  logic              [23:0] */ .igr_vp_rx_metadata         (igr0_vp_rx_metadata),                        
/* input  logic               [1:0] */ .igr_vp_rx_port_num         (igr0_vp_rx_port_num),                        
/* input  logic              [35:0] */ .igr_vp_rx_time_stamp       (igr0_vp_rx_time_stamp),                      
/* input  logic              [68:0] */ .mctagring_in_dn_0          ({69'b0}),                                    
/* input  logic              [68:0] */ .mctagring_in_dn_1          ({69'b0}),                                    
/* input  logic              [68:0] */ .mctagring_in_dn_2          ({69'b0}),                                    
/* input  logic              [68:0] */ .mctagring_in_dn_3          ({69'b0}),                                    
/* input  logic              [68:0] */ .mctagring_in_up_0          (mgp_mctagring_up_0),                         
/* input  logic              [68:0] */ .mctagring_in_up_1          (mgp_mctagring_up_1),                         
/* input  logic              [68:0] */ .mctagring_in_up_2          (mgp_mctagring_up_2),                         
/* input  logic              [68:0] */ .mctagring_in_up_3          (mgp_mctagring_up_3),                         
/* input  logic               [3:0] */ .mgp_id                     ({mpp_id[2:0],1'b0}),                         
/* input  logic              [33:0] */ .mrpodring_in_dn            (mpp_mrpodring_in_dn),                        
/* input  logic              [33:0] */ .mrpodring_in_up            (mgp_mrpodring_up),                           
/* input  logic                     */ .mrpodring_stall_in_dn      (mpp_mrpodring_stall_in_dn),                  
/* input  logic                     */ .mrpodring_stall_in_up      (mgp_mrpodring_stall_up),                     
/* input  logic              [33:0] */ .podring_in_dn              (mpp_podring_in_dn),                          
/* input  logic              [33:0] */ .podring_in_up              (mgp_podring_up),                             
/* input  logic                     */ .podring_stall_in_dn        (mpp_podring_stall_in_dn),                    
/* input  logic                     */ .podring_stall_in_up        (mgp_podring_stall_up),                       
/* input  logic                     */ .sreset                     (sreset),                                     
/* input  logic              [67:0] */ .tagring_in_dn_0_0          (mpp_tagring_in_dn_0_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_0_1          (mpp_tagring_in_dn_0_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_10_0         (mpp_tagring_in_dn_10_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_10_1         (mpp_tagring_in_dn_10_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_11_0         (mpp_tagring_in_dn_11_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_11_1         (mpp_tagring_in_dn_11_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_12_0         (mpp_tagring_in_dn_12_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_12_1         (mpp_tagring_in_dn_12_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_13_0         (mpp_tagring_in_dn_13_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_13_1         (mpp_tagring_in_dn_13_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_14_0         (mpp_tagring_in_dn_14_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_14_1         (mpp_tagring_in_dn_14_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_15_0         (mpp_tagring_in_dn_15_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_15_1         (mpp_tagring_in_dn_15_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_1_0          (mpp_tagring_in_dn_1_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_1_1          (mpp_tagring_in_dn_1_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_2_0          (mpp_tagring_in_dn_2_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_2_1          (mpp_tagring_in_dn_2_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_3_0          (mpp_tagring_in_dn_3_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_3_1          (mpp_tagring_in_dn_3_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_4_0          (mpp_tagring_in_dn_4_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_4_1          (mpp_tagring_in_dn_4_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_5_0          (mpp_tagring_in_dn_5_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_5_1          (mpp_tagring_in_dn_5_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_6_0          (mpp_tagring_in_dn_6_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_6_1          (mpp_tagring_in_dn_6_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_7_0          (mpp_tagring_in_dn_7_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_7_1          (mpp_tagring_in_dn_7_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_8_0          (mpp_tagring_in_dn_8_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_8_1          (mpp_tagring_in_dn_8_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_9_0          (mpp_tagring_in_dn_9_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_9_1          (mpp_tagring_in_dn_9_1),                      
/* input  logic              [67:0] */ .tagring_in_up_0_0          (mgp_tagring_up_0_0),                         
/* input  logic              [67:0] */ .tagring_in_up_0_1          (mgp_tagring_up_0_1),                         
/* input  logic              [67:0] */ .tagring_in_up_10_0         (mgp_tagring_up_10_0),                        
/* input  logic              [67:0] */ .tagring_in_up_10_1         (mgp_tagring_up_10_1),                        
/* input  logic              [67:0] */ .tagring_in_up_11_0         (mgp_tagring_up_11_0),                        
/* input  logic              [67:0] */ .tagring_in_up_11_1         (mgp_tagring_up_11_1),                        
/* input  logic              [67:0] */ .tagring_in_up_12_0         (mgp_tagring_up_12_0),                        
/* input  logic              [67:0] */ .tagring_in_up_12_1         (mgp_tagring_up_12_1),                        
/* input  logic              [67:0] */ .tagring_in_up_13_0         (mgp_tagring_up_13_0),                        
/* input  logic              [67:0] */ .tagring_in_up_13_1         (mgp_tagring_up_13_1),                        
/* input  logic              [67:0] */ .tagring_in_up_14_0         (mgp_tagring_up_14_0),                        
/* input  logic              [67:0] */ .tagring_in_up_14_1         (mgp_tagring_up_14_1),                        
/* input  logic              [67:0] */ .tagring_in_up_15_0         (mgp_tagring_up_15_0),                        
/* input  logic              [67:0] */ .tagring_in_up_15_1         (mgp_tagring_up_15_1),                        
/* input  logic              [67:0] */ .tagring_in_up_1_0          (mgp_tagring_up_1_0),                         
/* input  logic              [67:0] */ .tagring_in_up_1_1          (mgp_tagring_up_1_1),                         
/* input  logic              [67:0] */ .tagring_in_up_2_0          (mgp_tagring_up_2_0),                         
/* input  logic              [67:0] */ .tagring_in_up_2_1          (mgp_tagring_up_2_1),                         
/* input  logic              [67:0] */ .tagring_in_up_3_0          (mgp_tagring_up_3_0),                         
/* input  logic              [67:0] */ .tagring_in_up_3_1          (mgp_tagring_up_3_1),                         
/* input  logic              [67:0] */ .tagring_in_up_4_0          (mgp_tagring_up_4_0),                         
/* input  logic              [67:0] */ .tagring_in_up_4_1          (mgp_tagring_up_4_1),                         
/* input  logic              [67:0] */ .tagring_in_up_5_0          (mgp_tagring_up_5_0),                         
/* input  logic              [67:0] */ .tagring_in_up_5_1          (mgp_tagring_up_5_1),                         
/* input  logic              [67:0] */ .tagring_in_up_6_0          (mgp_tagring_up_6_0),                         
/* input  logic              [67:0] */ .tagring_in_up_6_1          (mgp_tagring_up_6_1),                         
/* input  logic              [67:0] */ .tagring_in_up_7_0          (mgp_tagring_up_7_0),                         
/* input  logic              [67:0] */ .tagring_in_up_7_1          (mgp_tagring_up_7_1),                         
/* input  logic              [67:0] */ .tagring_in_up_8_0          (mgp_tagring_up_8_0),                         
/* input  logic              [67:0] */ .tagring_in_up_8_1          (mgp_tagring_up_8_1),                         
/* input  logic              [67:0] */ .tagring_in_up_9_0          (mgp_tagring_up_9_0),                         
/* input  logic              [67:0] */ .tagring_in_up_9_1          (mgp_tagring_up_9_1),                         
/* Interface ahb_rx_ppe_if.ppe      */ .ahb_rxppe                  (ahb0_rxppe),                                 
/* Interface ahb_rx_ppe_if.ppe      */ .ahb_txppe0                 (ahb0_txppe0),                                
/* Interface ahb_rx_ppe_if.ppe      */ .ahb_txppe1                 (ahb0_txppe1),                                
/* Interface egr_ahb_if.egr         */ .egr_ahb                    (egr0_ahb),                                   
/* Interface egr_cmring_if.egr      */ .egr_cmring                 (egr_cmring),                                 
/* Interface egr_epl_if.egr         */ .egr_epl0                   (grp_a0),                                     
/* Interface egr_epl_if.egr         */ .egr_epl1                   (grp_b0),                                     
/* Interface egr_epl_if.egr         */ .egr_epl2                   (grp_c0),                                     
/* Interface egr_epl_if.egr         */ .egr_epl3                   (grp_d0),                                     
/* Interface egr_mc_table_if.egr    */ .egr_mc_table0              (egr0_mc_table0),                             
/* Interface egr_mc_table_if.egr    */ .egr_mc_table1              (egr0_mc_table1),                             
/* Interface egr_ppe_stm_if.egr     */ .egr_ppestm                 (egr0_ppestm),                                
/* Interface glb_rx_ppe_if.ppe      */ .glb_rxppe                  (glb0_rxppe),                                 
/* Interface glb_rx_ppe_if.ppe      */ .glb_txppe0                 (glb0_txppe0),                                
/* Interface glb_rx_ppe_if.ppe      */ .glb_txppe1                 (glb0_txppe1),                                
/* Interface mim_rd_if.request      */ .mim0_rd0                   (mim0_rd0),                                   
/* Interface mim_rd_if.request      */ .mim0_rd1                   (mim0_rd1),                                   
/* Interface mim_rd_if.request      */ .mim0_rd2                   (mim0_rd2),                                   
/* Interface mim_wr_if.request      */ .mim0_wr0                   (mim0_wr0),                                   
/* Interface mim_wr_if.request      */ .mim0_wr1                   (mim0_wr1),                                   
/* Interface mim_wr_if.request      */ .mim0_wr2                   (mim0_wr2),                                   
/* Interface mim_rd_if.request      */ .mim1_rd0                   (mim1_rd0),                                   
/* Interface mim_rd_if.request      */ .mim1_rd1                   (mim1_rd1),                                   
/* Interface mim_rd_if.request      */ .mim1_rd2                   (mim1_rd2),                                   
/* Interface mim_wr_if.request      */ .mim1_wr0                   (mim1_wr0),                                   
/* Interface mim_wr_if.request      */ .mim1_wr1                   (mim1_wr1),                                   
/* Interface mim_wr_if.request      */ .mim1_wr2                   (mim1_wr2),                                   
/* Interface rx_ppe_ppe_stm0_if.ppe */ .rxppe_ppestm0              (rxppe0_ppestm0),                             
/* Interface rx_ppe_ppe_stm1_if.ppe */ .rxppe_ppestm1              (rxppe0_ppestm1),                             
/* output logic              [23:0] */ .dqring_out_dn_0_0          (mgp_dqring_dn_0_0),                          
/* output logic              [23:0] */ .dqring_out_dn_0_1          (mgp_dqring_dn_0_1),                          
/* output logic              [23:0] */ .dqring_out_dn_1_0          (mgp_dqring_dn_1_0),                          
/* output logic              [23:0] */ .dqring_out_dn_1_1          (mgp_dqring_dn_1_1),                          
/* output logic              [23:0] */ .dqring_out_dn_2_0          (mgp_dqring_dn_2_0),                          
/* output logic              [23:0] */ .dqring_out_dn_2_1          (mgp_dqring_dn_2_1),                          
/* output logic              [23:0] */ .dqring_out_dn_3_0          (mgp_dqring_dn_3_0),                          
/* output logic              [23:0] */ .dqring_out_dn_3_1          (mgp_dqring_dn_3_1),                          
/* output logic              [23:0] */ .dqring_out_dn_4_0          (mgp_dqring_dn_4_0),                          
/* output logic              [23:0] */ .dqring_out_dn_4_1          (mgp_dqring_dn_4_1),                          
/* output logic              [23:0] */ .dqring_out_dn_5_0          (mgp_dqring_dn_5_0),                          
/* output logic              [23:0] */ .dqring_out_dn_5_1          (mgp_dqring_dn_5_1),                          
/* output logic              [23:0] */ .dqring_out_dn_6_0          (mgp_dqring_dn_6_0),                          
/* output logic              [23:0] */ .dqring_out_dn_6_1          (mgp_dqring_dn_6_1),                          
/* output logic              [23:0] */ .dqring_out_dn_7_0          (mgp_dqring_dn_7_0),                          
/* output logic              [23:0] */ .dqring_out_dn_7_1          (mgp_dqring_dn_7_1),                          
/* output logic              [23:0] */ .dqring_out_up_0_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_0_1          (),                                           
/* output logic              [23:0] */ .dqring_out_up_1_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_1_1          (),                                           
/* output logic              [23:0] */ .dqring_out_up_2_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_2_1          (),                                           
/* output logic              [23:0] */ .dqring_out_up_3_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_3_1          (),                                           
/* output logic              [23:0] */ .dqring_out_up_4_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_4_1          (),                                           
/* output logic              [23:0] */ .dqring_out_up_5_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_5_1          (),                                           
/* output logic              [23:0] */ .dqring_out_up_6_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_6_1          (),                                           
/* output logic              [23:0] */ .dqring_out_up_7_0          (),                                           
/* output logic              [23:0] */ .dqring_out_up_7_1          (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_0_0        (mgp_gpolring_dn_0_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_0_1        (mgp_gpolring_dn_0_1),                        
/* output logic              [25:0] */ .gpolring_out_dn_1_0        (mgp_gpolring_dn_1_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_1_1        (mgp_gpolring_dn_1_1),                        
/* output logic              [25:0] */ .gpolring_out_dn_2_0        (mgp_gpolring_dn_2_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_2_1        (mgp_gpolring_dn_2_1),                        
/* output logic              [25:0] */ .gpolring_out_dn_3_0        (mgp_gpolring_dn_3_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_3_1        (mgp_gpolring_dn_3_1),                        
/* output logic              [25:0] */ .gpolring_out_dn_4_0        (mgp_gpolring_dn_4_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_4_1        (mgp_gpolring_dn_4_1),                        
/* output logic              [25:0] */ .gpolring_out_dn_5_0        (mgp_gpolring_dn_5_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_5_1        (mgp_gpolring_dn_5_1),                        
/* output logic              [25:0] */ .gpolring_out_dn_6_0        (mgp_gpolring_dn_6_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_6_1        (mgp_gpolring_dn_6_1),                        
/* output logic              [25:0] */ .gpolring_out_dn_7_0        (mgp_gpolring_dn_7_0),                        
/* output logic              [25:0] */ .gpolring_out_dn_7_1        (mgp_gpolring_dn_7_1),                        
/* output logic              [25:0] */ .gpolring_out_up_0_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_0_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_1_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_1_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_2_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_2_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_3_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_3_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_4_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_4_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_5_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_5_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_6_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_6_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_7_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_7_1        (),                                           
/* output logic             [106:0] */ .gpolring_update_out_dn_0   (mgp_gpolring_update_dn_0),                   
/* output logic             [106:0] */ .gpolring_update_out_dn_1   (mgp_gpolring_update_dn_1),                   
/* output logic             [106:0] */ .gpolring_update_out_up_0   (),                                           
/* output logic             [106:0] */ .gpolring_update_out_up_1   (),                                           
/* output logic                     */ .grp_a_tx_pfc_tc_sync       (grp_a0_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_a_tx_pfc_xoff          (grp_a0_tx_pfc_xoff),                         
/* output logic                     */ .grp_b_tx_pfc_tc_sync       (grp_b0_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_b_tx_pfc_xoff          (grp_b0_tx_pfc_xoff),                         
/* output logic                     */ .grp_c_tx_pfc_tc_sync       (grp_c0_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_c_tx_pfc_xoff          (grp_c0_tx_pfc_xoff),                         
/* output logic                     */ .grp_d_tx_pfc_tc_sync       (grp_d0_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_d_tx_pfc_xoff          (grp_d0_tx_pfc_xoff),                         
/* output logic                     */ .igr_vp_tx_pfc_xoff         (igr0_vp_tx_pfc_xoff),                        //FIXME should this be [1:0] for 2 VP   
/* output logic              [68:0] */ .mctagring_out_dn_0         (mgp_mctagring_dn_0),                         
/* output logic              [68:0] */ .mctagring_out_dn_1         (mgp_mctagring_dn_1),                         
/* output logic              [68:0] */ .mctagring_out_dn_2         (mgp_mctagring_dn_2),                         
/* output logic              [68:0] */ .mctagring_out_dn_3         (mgp_mctagring_dn_3),                         
/* output logic              [68:0] */ .mctagring_out_up_0         (mpp_mctagring_out_0),                        
/* output logic              [68:0] */ .mctagring_out_up_1         (mpp_mctagring_out_1),                        
/* output logic              [68:0] */ .mctagring_out_up_2         (mpp_mctagring_out_2),                        
/* output logic              [68:0] */ .mctagring_out_up_3         (mpp_mctagring_out_3),                        
/* output logic              [33:0] */ .mrpodring_out_dn           (mgp_mrpodring_dn),                           
/* output logic              [33:0] */ .mrpodring_out_up           (mpp_mrpodring_out_up),                       
/* output logic                     */ .mrpodring_stall_out_dn     (mgp_mrpodring_stall_dn),                     
/* output logic                     */ .mrpodring_stall_out_up     (mpp_mrpodring_stall_out_up),                 
/* output logic              [33:0] */ .podring_out_dn             (mgp_podring_dn),                             
/* output logic              [33:0] */ .podring_out_up             (mpp_podring_out_up),                         
/* output logic                     */ .podring_stall_out_dn       (mgp_podring_stall_dn),                       
/* output logic                     */ .podring_stall_out_up       (mpp_podring_stall_out_up),                   
/* output logic              [67:0] */ .tagring_out_dn_0_0         (mgp_tagring_dn_0_0),                         
/* output logic              [67:0] */ .tagring_out_dn_0_1         (mgp_tagring_dn_0_1),                         
/* output logic              [67:0] */ .tagring_out_dn_10_0        (mgp_tagring_dn_10_0),                        
/* output logic              [67:0] */ .tagring_out_dn_10_1        (mgp_tagring_dn_10_1),                        
/* output logic              [67:0] */ .tagring_out_dn_11_0        (mgp_tagring_dn_11_0),                        
/* output logic              [67:0] */ .tagring_out_dn_11_1        (mgp_tagring_dn_11_1),                        
/* output logic              [67:0] */ .tagring_out_dn_12_0        (mgp_tagring_dn_12_0),                        
/* output logic              [67:0] */ .tagring_out_dn_12_1        (mgp_tagring_dn_12_1),                        
/* output logic              [67:0] */ .tagring_out_dn_13_0        (mgp_tagring_dn_13_0),                        
/* output logic              [67:0] */ .tagring_out_dn_13_1        (mgp_tagring_dn_13_1),                        
/* output logic              [67:0] */ .tagring_out_dn_14_0        (mgp_tagring_dn_14_0),                        
/* output logic              [67:0] */ .tagring_out_dn_14_1        (mgp_tagring_dn_14_1),                        
/* output logic              [67:0] */ .tagring_out_dn_15_0        (mgp_tagring_dn_15_0),                        
/* output logic              [67:0] */ .tagring_out_dn_15_1        (mgp_tagring_dn_15_1),                        
/* output logic              [67:0] */ .tagring_out_dn_1_0         (mgp_tagring_dn_1_0),                         
/* output logic              [67:0] */ .tagring_out_dn_1_1         (mgp_tagring_dn_1_1),                         
/* output logic              [67:0] */ .tagring_out_dn_2_0         (mgp_tagring_dn_2_0),                         
/* output logic              [67:0] */ .tagring_out_dn_2_1         (mgp_tagring_dn_2_1),                         
/* output logic              [67:0] */ .tagring_out_dn_3_0         (mgp_tagring_dn_3_0),                         
/* output logic              [67:0] */ .tagring_out_dn_3_1         (mgp_tagring_dn_3_1),                         
/* output logic              [67:0] */ .tagring_out_dn_4_0         (mgp_tagring_dn_4_0),                         
/* output logic              [67:0] */ .tagring_out_dn_4_1         (mgp_tagring_dn_4_1),                         
/* output logic              [67:0] */ .tagring_out_dn_5_0         (mgp_tagring_dn_5_0),                         
/* output logic              [67:0] */ .tagring_out_dn_5_1         (mgp_tagring_dn_5_1),                         
/* output logic              [67:0] */ .tagring_out_dn_6_0         (mgp_tagring_dn_6_0),                         
/* output logic              [67:0] */ .tagring_out_dn_6_1         (mgp_tagring_dn_6_1),                         
/* output logic              [67:0] */ .tagring_out_dn_7_0         (mgp_tagring_dn_7_0),                         
/* output logic              [67:0] */ .tagring_out_dn_7_1         (mgp_tagring_dn_7_1),                         
/* output logic              [67:0] */ .tagring_out_dn_8_0         (mgp_tagring_dn_8_0),                         
/* output logic              [67:0] */ .tagring_out_dn_8_1         (mgp_tagring_dn_8_1),                         
/* output logic              [67:0] */ .tagring_out_dn_9_0         (mgp_tagring_dn_9_0),                         
/* output logic              [67:0] */ .tagring_out_dn_9_1         (mgp_tagring_dn_9_1),                         
/* output logic              [67:0] */ .tagring_out_up_0_0         (mpp_tagring_out_up_0_0),                     
/* output logic              [67:0] */ .tagring_out_up_0_1         (mpp_tagring_out_up_0_1),                     
/* output logic              [67:0] */ .tagring_out_up_10_0        (mpp_tagring_out_up_10_0),                    
/* output logic              [67:0] */ .tagring_out_up_10_1        (mpp_tagring_out_up_10_1),                    
/* output logic              [67:0] */ .tagring_out_up_11_0        (mpp_tagring_out_up_11_0),                    
/* output logic              [67:0] */ .tagring_out_up_11_1        (mpp_tagring_out_up_11_1),                    
/* output logic              [67:0] */ .tagring_out_up_12_0        (mpp_tagring_out_up_12_0),                    
/* output logic              [67:0] */ .tagring_out_up_12_1        (mpp_tagring_out_up_12_1),                    
/* output logic              [67:0] */ .tagring_out_up_13_0        (mpp_tagring_out_up_13_0),                    
/* output logic              [67:0] */ .tagring_out_up_13_1        (mpp_tagring_out_up_13_1),                    
/* output logic              [67:0] */ .tagring_out_up_14_0        (mpp_tagring_out_up_14_0),                    
/* output logic              [67:0] */ .tagring_out_up_14_1        (mpp_tagring_out_up_14_1),                    
/* output logic              [67:0] */ .tagring_out_up_15_0        (mpp_tagring_out_up_15_0),                    
/* output logic              [67:0] */ .tagring_out_up_15_1        (mpp_tagring_out_up_15_1),                    
/* output logic              [67:0] */ .tagring_out_up_1_0         (mpp_tagring_out_up_1_0),                     
/* output logic              [67:0] */ .tagring_out_up_1_1         (mpp_tagring_out_up_1_1),                     
/* output logic              [67:0] */ .tagring_out_up_2_0         (mpp_tagring_out_up_2_0),                     
/* output logic              [67:0] */ .tagring_out_up_2_1         (mpp_tagring_out_up_2_1),                     
/* output logic              [67:0] */ .tagring_out_up_3_0         (mpp_tagring_out_up_3_0),                     
/* output logic              [67:0] */ .tagring_out_up_3_1         (mpp_tagring_out_up_3_1),                     
/* output logic              [67:0] */ .tagring_out_up_4_0         (mpp_tagring_out_up_4_0),                     
/* output logic              [67:0] */ .tagring_out_up_4_1         (mpp_tagring_out_up_4_1),                     
/* output logic              [67:0] */ .tagring_out_up_5_0         (mpp_tagring_out_up_5_0),                     
/* output logic              [67:0] */ .tagring_out_up_5_1         (mpp_tagring_out_up_5_1),                     
/* output logic              [67:0] */ .tagring_out_up_6_0         (mpp_tagring_out_up_6_0),                     
/* output logic              [67:0] */ .tagring_out_up_6_1         (mpp_tagring_out_up_6_1),                     
/* output logic              [67:0] */ .tagring_out_up_7_0         (mpp_tagring_out_up_7_0),                     
/* output logic              [67:0] */ .tagring_out_up_7_1         (mpp_tagring_out_up_7_1),                     
/* output logic              [67:0] */ .tagring_out_up_8_0         (mpp_tagring_out_up_8_0),                     
/* output logic              [67:0] */ .tagring_out_up_8_1         (mpp_tagring_out_up_8_1),                     
/* output logic              [67:0] */ .tagring_out_up_9_0         (mpp_tagring_out_up_9_0),                     
/* output logic              [67:0] */ .tagring_out_up_9_1         (mpp_tagring_out_up_9_1));                     
// End of module mgp0 from mby_mgp


// module mgp1    from mby_mgp using mgp.map 1
mby_mgp    mgp1(
/* input  logic                     */ .arst_n                     (arst_n),                                     //Asynchronous negedge reset     
/* input  logic                     */ .cclk                       (cclk),                                       
/* input  logic              [23:0] */ .dqring_in_dn_0_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_0_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_1_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_1_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_2_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_2_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_3_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_3_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_4_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_4_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_5_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_5_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_6_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_6_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_7_0           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_dn_7_1           ({24'b0}),                                    
/* input  logic              [23:0] */ .dqring_in_up_0_0           (mgp_dqring_dn_0_0),                          
/* input  logic              [23:0] */ .dqring_in_up_0_1           (mgp_dqring_dn_0_1),                          
/* input  logic              [23:0] */ .dqring_in_up_1_0           (mgp_dqring_dn_1_0),                          
/* input  logic              [23:0] */ .dqring_in_up_1_1           (mgp_dqring_dn_1_1),                          
/* input  logic              [23:0] */ .dqring_in_up_2_0           (mgp_dqring_dn_2_0),                          
/* input  logic              [23:0] */ .dqring_in_up_2_1           (mgp_dqring_dn_2_1),                          
/* input  logic              [23:0] */ .dqring_in_up_3_0           (mgp_dqring_dn_3_0),                          
/* input  logic              [23:0] */ .dqring_in_up_3_1           (mgp_dqring_dn_3_1),                          
/* input  logic              [23:0] */ .dqring_in_up_4_0           (mgp_dqring_dn_4_0),                          
/* input  logic              [23:0] */ .dqring_in_up_4_1           (mgp_dqring_dn_4_1),                          
/* input  logic              [23:0] */ .dqring_in_up_5_0           (mgp_dqring_dn_5_0),                          
/* input  logic              [23:0] */ .dqring_in_up_5_1           (mgp_dqring_dn_5_1),                          
/* input  logic              [23:0] */ .dqring_in_up_6_0           (mgp_dqring_dn_6_0),                          
/* input  logic              [23:0] */ .dqring_in_up_6_1           (mgp_dqring_dn_6_1),                          
/* input  logic              [23:0] */ .dqring_in_up_7_0           (mgp_dqring_dn_7_0),                          
/* input  logic              [23:0] */ .dqring_in_up_7_1           (mgp_dqring_dn_7_1),                          
/* input  logic              [25:0] */ .gpolring_in_dn_0_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_0_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_1_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_1_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_2_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_2_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_3_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_3_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_4_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_4_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_5_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_5_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_6_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_6_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_7_0         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_dn_7_1         ({26'b0}),                                    
/* input  logic              [25:0] */ .gpolring_in_up_0_0         (mgp_gpolring_dn_0_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_0_1         (mgp_gpolring_dn_0_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_1_0         (mgp_gpolring_dn_1_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_1_1         (mgp_gpolring_dn_1_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_2_0         (mgp_gpolring_dn_2_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_2_1         (mgp_gpolring_dn_2_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_3_0         (mgp_gpolring_dn_3_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_3_1         (mgp_gpolring_dn_3_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_4_0         (mgp_gpolring_dn_4_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_4_1         (mgp_gpolring_dn_4_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_5_0         (mgp_gpolring_dn_5_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_5_1         (mgp_gpolring_dn_5_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_6_0         (mgp_gpolring_dn_6_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_6_1         (mgp_gpolring_dn_6_1),                        
/* input  logic              [25:0] */ .gpolring_in_up_7_0         (mgp_gpolring_dn_7_0),                        
/* input  logic              [25:0] */ .gpolring_in_up_7_1         (mgp_gpolring_dn_7_1),                        
/* input  logic             [106:0] */ .gpolring_update_in_dn_0    ({107'b0}),                                   
/* input  logic             [106:0] */ .gpolring_update_in_dn_1    ({107'b0}),                                   
/* input  logic             [106:0] */ .gpolring_update_in_up_0    (mgp_gpolring_update_dn_0),                   
/* input  logic             [106:0] */ .gpolring_update_in_up_1    (mgp_gpolring_update_dn_1),                   
/* input  logic         [0:7][63:0] */ .grp_a_rx_data              ({grp_a1_rx0_data[63:0], grp_a1_rx1_data[63:0], grp_a1_rx2_data[63:0], grp_a1_rx3_data[63:0], grp_a1_rx4_data[63:0], grp_a1_rx5_data[63:0], grp_a1_rx6_data[63:0], grp_a1_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_a_rx_data_valid        (grp_a1_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_a_rx_metadata          ({grp_a1_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_a_rx_port_num          (grp_a1_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_a_rx_time_stamp        ({grp_a1_rx_time_stamp[39:0]}),               
/* input  logic         [0:7][63:0] */ .grp_b_rx_data              ({grp_b1_rx0_data[63:0], grp_b1_rx1_data[63:0], grp_b1_rx2_data[63:0], grp_b1_rx3_data[63:0], grp_b1_rx4_data[63:0], grp_b1_rx5_data[63:0], grp_b1_rx6_data[63:0], grp_b1_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_b_rx_data_valid        (grp_b1_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_b_rx_metadata          ({grp_b1_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_b_rx_port_num          (grp_b1_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_b_rx_time_stamp        ({grp_b1_rx_time_stamp[39:0]}),               
/* input  logic         [0:7][63:0] */ .grp_c_rx_data              ({grp_c1_rx0_data[63:0], grp_c1_rx1_data[63:0], grp_c1_rx2_data[63:0], grp_c1_rx3_data[63:0], grp_c1_rx4_data[63:0], grp_c1_rx5_data[63:0], grp_c1_rx6_data[63:0], grp_c1_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_c_rx_data_valid        (grp_c1_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_c_rx_metadata          ({grp_c1_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_c_rx_port_num          (grp_c1_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_c_rx_time_stamp        ({grp_c1_rx_time_stamp[39:0]}),               
/* input  logic         [0:7][63:0] */ .grp_d_rx_data              ({grp_d1_rx0_data[63:0], grp_d1_rx1_data[63:0], grp_d1_rx2_data[63:0], grp_d1_rx3_data[63:0], grp_d1_rx4_data[63:0], grp_d1_rx5_data[63:0], grp_d1_rx6_data[63:0], grp_d1_rx7_data[63:0]}), 
/* input  logic               [7:0] */ .grp_d_rx_data_valid        (grp_d1_rx_data_valid),                       
/* input  logic  [EPL_IGR_MD_MSB:0] */ .grp_d_rx_metadata          ({grp_d1_rx_metadata[23:0]}),                 
/* input  logic               [1:0] */ .grp_d_rx_port_num          (grp_d1_rx_port_num),                         
/* input  logic  [EPL_IGR_TS_MSB:0] */ .grp_d_rx_time_stamp        ({grp_d1_rx_time_stamp[39:0]}),               
/* input  logic              [19:0] */ .igr_vp_cpp_rx_metadata     (igr1_vp_cpp_rx_metadata),                    
/* input  logic               [7:0] */ .igr_vp_rx_data_valid       (igr1_vp_rx_data_valid),                      
/* input  logic         [0:7][71:0] */ .igr_vp_rx_data_w_ecc       ({igr1_vp_rx0_data_w_ecc[71:0], igr1_vp_rx1_data_w_ecc[71:0], igr1_vp_rx2_data_w_ecc[71:0], igr1_vp_rx3_data_w_ecc[71:0], igr1_vp_rx4_data_w_ecc[71:0], igr1_vp_rx5_data_w_ecc[71:0], igr1_vp_rx6_data_w_ecc[71:0], igr1_vp_rx7_data_w_ecc[71:0]}), 
/* input  logic               [7:0] */ .igr_vp_rx_ecc              (igr1_vp_rx_ecc),                             
/* input  logic               [2:0] */ .igr_vp_rx_flow_control_tc  (igr1_vp_rx_flow_control_tc),                 
/* input  logic              [23:0] */ .igr_vp_rx_metadata         (igr1_vp_rx_metadata),                        
/* input  logic               [1:0] */ .igr_vp_rx_port_num         (igr1_vp_rx_port_num),                        
/* input  logic              [35:0] */ .igr_vp_rx_time_stamp       (igr1_vp_rx_time_stamp),                      
/* input  logic              [68:0] */ .mctagring_in_dn_0          (mpp_mctagring_in_0),                         
/* input  logic              [68:0] */ .mctagring_in_dn_1          (mpp_mctagring_in_1),                         
/* input  logic              [68:0] */ .mctagring_in_dn_2          (mpp_mctagring_in_2),                         
/* input  logic              [68:0] */ .mctagring_in_dn_3          (mpp_mctagring_in_3),                         
/* input  logic              [68:0] */ .mctagring_in_up_0          (mgp_mctagring_dn_0),                         
/* input  logic              [68:0] */ .mctagring_in_up_1          (mgp_mctagring_dn_1),                         
/* input  logic              [68:0] */ .mctagring_in_up_2          (mgp_mctagring_dn_2),                         
/* input  logic              [68:0] */ .mctagring_in_up_3          (mgp_mctagring_dn_3),                         
/* input  logic               [3:0] */ .mgp_id                     ({mpp_id[2:0],1'b1}),                         
/* input  logic              [33:0] */ .mrpodring_in_dn            (mpp_mrpodring_in_up),                        
/* input  logic              [33:0] */ .mrpodring_in_up            (mgp_mrpodring_dn),                           
/* input  logic                     */ .mrpodring_stall_in_dn      (mpp_mrpodring_stall_in_up),                  
/* input  logic                     */ .mrpodring_stall_in_up      (mgp_mrpodring_stall_dn),                     
/* input  logic              [33:0] */ .podring_in_dn              (mpp_podring_in_up),                          
/* input  logic              [33:0] */ .podring_in_up              (mgp_podring_dn),                             
/* input  logic                     */ .podring_stall_in_dn        (mpp_podring_stall_in_up),                    
/* input  logic                     */ .podring_stall_in_up        (mgp_podring_stall_dn),                       
/* input  logic                     */ .sreset                     (sreset),                                     
/* input  logic              [67:0] */ .tagring_in_dn_0_0          (mpp_tagring_in_up_0_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_0_1          (mpp_tagring_in_up_0_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_10_0         (mpp_tagring_in_up_10_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_10_1         (mpp_tagring_in_up_10_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_11_0         (mpp_tagring_in_up_11_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_11_1         (mpp_tagring_in_up_11_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_12_0         (mpp_tagring_in_up_12_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_12_1         (mpp_tagring_in_up_12_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_13_0         (mpp_tagring_in_up_13_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_13_1         (mpp_tagring_in_up_13_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_14_0         (mpp_tagring_in_up_14_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_14_1         (mpp_tagring_in_up_14_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_15_0         (mpp_tagring_in_up_15_0),                     
/* input  logic              [67:0] */ .tagring_in_dn_15_1         (mpp_tagring_in_up_15_1),                     
/* input  logic              [67:0] */ .tagring_in_dn_1_0          (mpp_tagring_in_up_1_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_1_1          (mpp_tagring_in_up_1_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_2_0          (mpp_tagring_in_up_2_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_2_1          (mpp_tagring_in_up_2_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_3_0          (mpp_tagring_in_up_3_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_3_1          (mpp_tagring_in_up_3_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_4_0          (mpp_tagring_in_up_4_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_4_1          (mpp_tagring_in_up_4_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_5_0          (mpp_tagring_in_up_5_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_5_1          (mpp_tagring_in_up_5_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_6_0          (mpp_tagring_in_up_6_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_6_1          (mpp_tagring_in_up_6_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_7_0          (mpp_tagring_in_up_7_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_7_1          (mpp_tagring_in_up_7_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_8_0          (mpp_tagring_in_up_8_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_8_1          (mpp_tagring_in_up_8_1),                      
/* input  logic              [67:0] */ .tagring_in_dn_9_0          (mpp_tagring_in_up_9_0),                      
/* input  logic              [67:0] */ .tagring_in_dn_9_1          (mpp_tagring_in_up_9_1),                      
/* input  logic              [67:0] */ .tagring_in_up_0_0          (mgp_tagring_dn_0_0),                         
/* input  logic              [67:0] */ .tagring_in_up_0_1          (mgp_tagring_dn_0_1),                         
/* input  logic              [67:0] */ .tagring_in_up_10_0         (mgp_tagring_dn_10_0),                        
/* input  logic              [67:0] */ .tagring_in_up_10_1         (mgp_tagring_dn_10_1),                        
/* input  logic              [67:0] */ .tagring_in_up_11_0         (mgp_tagring_dn_11_0),                        
/* input  logic              [67:0] */ .tagring_in_up_11_1         (mgp_tagring_dn_11_1),                        
/* input  logic              [67:0] */ .tagring_in_up_12_0         (mgp_tagring_dn_12_0),                        
/* input  logic              [67:0] */ .tagring_in_up_12_1         (mgp_tagring_dn_12_1),                        
/* input  logic              [67:0] */ .tagring_in_up_13_0         (mgp_tagring_dn_13_0),                        
/* input  logic              [67:0] */ .tagring_in_up_13_1         (mgp_tagring_dn_13_1),                        
/* input  logic              [67:0] */ .tagring_in_up_14_0         (mgp_tagring_dn_14_0),                        
/* input  logic              [67:0] */ .tagring_in_up_14_1         (mgp_tagring_dn_14_1),                        
/* input  logic              [67:0] */ .tagring_in_up_15_0         (mgp_tagring_dn_15_0),                        
/* input  logic              [67:0] */ .tagring_in_up_15_1         (mgp_tagring_dn_15_1),                        
/* input  logic              [67:0] */ .tagring_in_up_1_0          (mgp_tagring_dn_1_0),                         
/* input  logic              [67:0] */ .tagring_in_up_1_1          (mgp_tagring_dn_1_1),                         
/* input  logic              [67:0] */ .tagring_in_up_2_0          (mgp_tagring_dn_2_0),                         
/* input  logic              [67:0] */ .tagring_in_up_2_1          (mgp_tagring_dn_2_1),                         
/* input  logic              [67:0] */ .tagring_in_up_3_0          (mgp_tagring_dn_3_0),                         
/* input  logic              [67:0] */ .tagring_in_up_3_1          (mgp_tagring_dn_3_1),                         
/* input  logic              [67:0] */ .tagring_in_up_4_0          (mgp_tagring_dn_4_0),                         
/* input  logic              [67:0] */ .tagring_in_up_4_1          (mgp_tagring_dn_4_1),                         
/* input  logic              [67:0] */ .tagring_in_up_5_0          (mgp_tagring_dn_5_0),                         
/* input  logic              [67:0] */ .tagring_in_up_5_1          (mgp_tagring_dn_5_1),                         
/* input  logic              [67:0] */ .tagring_in_up_6_0          (mgp_tagring_dn_6_0),                         
/* input  logic              [67:0] */ .tagring_in_up_6_1          (mgp_tagring_dn_6_1),                         
/* input  logic              [67:0] */ .tagring_in_up_7_0          (mgp_tagring_dn_7_0),                         
/* input  logic              [67:0] */ .tagring_in_up_7_1          (mgp_tagring_dn_7_1),                         
/* input  logic              [67:0] */ .tagring_in_up_8_0          (mgp_tagring_dn_8_0),                         
/* input  logic              [67:0] */ .tagring_in_up_8_1          (mgp_tagring_dn_8_1),                         
/* input  logic              [67:0] */ .tagring_in_up_9_0          (mgp_tagring_dn_9_0),                         
/* input  logic              [67:0] */ .tagring_in_up_9_1          (mgp_tagring_dn_9_1),                         
/* Interface ahb_rx_ppe_if.ppe      */ .ahb_rxppe                  (ahb1_rxppe),                                 
/* Interface ahb_rx_ppe_if.ppe      */ .ahb_txppe0                 (ahb1_txppe0),                                
/* Interface ahb_rx_ppe_if.ppe      */ .ahb_txppe1                 (ahb1_txppe1),                                
/* Interface egr_ahb_if.egr         */ .egr_ahb                    (egr1_ahb),                                   
/* Interface egr_cmring_if.egr      */ .egr_cmring                 (egr_cmring),                                 
/* Interface egr_epl_if.egr         */ .egr_epl0                   (grp_a1),                                     
/* Interface egr_epl_if.egr         */ .egr_epl1                   (grp_b1),                                     
/* Interface egr_epl_if.egr         */ .egr_epl2                   (grp_c1),                                     
/* Interface egr_epl_if.egr         */ .egr_epl3                   (grp_d1),                                     
/* Interface egr_mc_table_if.egr    */ .egr_mc_table0              (egr1_mc_table0),                             
/* Interface egr_mc_table_if.egr    */ .egr_mc_table1              (egr1_mc_table1),                             
/* Interface egr_ppe_stm_if.egr     */ .egr_ppestm                 (egr1_ppestm),                                
/* Interface glb_rx_ppe_if.ppe      */ .glb_rxppe                  (glb1_rxppe),                                 
/* Interface glb_rx_ppe_if.ppe      */ .glb_txppe0                 (glb1_txppe0),                                
/* Interface glb_rx_ppe_if.ppe      */ .glb_txppe1                 (glb1_txppe1),                                
/* Interface mim_rd_if.request      */ .mim0_rd0                   (mim2_rd0),                                   
/* Interface mim_rd_if.request      */ .mim0_rd1                   (mim2_rd1),                                   
/* Interface mim_rd_if.request      */ .mim0_rd2                   (mim2_rd2),                                   
/* Interface mim_wr_if.request      */ .mim0_wr0                   (mim2_wr0),                                   
/* Interface mim_wr_if.request      */ .mim0_wr1                   (mim2_wr1),                                   
/* Interface mim_wr_if.request      */ .mim0_wr2                   (mim2_wr2),                                   
/* Interface mim_rd_if.request      */ .mim1_rd0                   (mim3_rd0),                                   
/* Interface mim_rd_if.request      */ .mim1_rd1                   (mim3_rd1),                                   
/* Interface mim_rd_if.request      */ .mim1_rd2                   (mim3_rd2),                                   
/* Interface mim_wr_if.request      */ .mim1_wr0                   (mim3_wr0),                                   
/* Interface mim_wr_if.request      */ .mim1_wr1                   (mim3_wr1),                                   
/* Interface mim_wr_if.request      */ .mim1_wr2                   (mim3_wr2),                                   
/* Interface rx_ppe_ppe_stm0_if.ppe */ .rxppe_ppestm0              (rxppe1_ppestm0),                             
/* Interface rx_ppe_ppe_stm1_if.ppe */ .rxppe_ppestm1              (rxppe1_ppestm1),                             
/* output logic              [23:0] */ .dqring_out_dn_0_0          (mgp_dqring_up_0_0),                          
/* output logic              [23:0] */ .dqring_out_dn_0_1          (mgp_dqring_up_0_1),                          
/* output logic              [23:0] */ .dqring_out_dn_1_0          (mgp_dqring_up_1_0),                          
/* output logic              [23:0] */ .dqring_out_dn_1_1          (mgp_dqring_up_1_1),                          
/* output logic              [23:0] */ .dqring_out_dn_2_0          (mgp_dqring_up_2_0),                          
/* output logic              [23:0] */ .dqring_out_dn_2_1          (mgp_dqring_up_2_1),                          
/* output logic              [23:0] */ .dqring_out_dn_3_0          (mgp_dqring_up_3_0),                          
/* output logic              [23:0] */ .dqring_out_dn_3_1          (mgp_dqring_up_3_1),                          
/* output logic              [23:0] */ .dqring_out_dn_4_0          (mgp_dqring_up_4_0),                          
/* output logic              [23:0] */ .dqring_out_dn_4_1          (mgp_dqring_up_4_1),                          
/* output logic              [23:0] */ .dqring_out_dn_5_0          (mgp_dqring_up_5_0),                          
/* output logic              [23:0] */ .dqring_out_dn_5_1          (mgp_dqring_up_5_1),                          
/* output logic              [23:0] */ .dqring_out_dn_6_0          (mgp_dqring_up_6_0),                          
/* output logic              [23:0] */ .dqring_out_dn_6_1          (mgp_dqring_up_6_1),                          
/* output logic              [23:0] */ .dqring_out_dn_7_0          (mgp_dqring_up_7_0),                          
/* output logic              [23:0] */ .dqring_out_dn_7_1          (mgp_dqring_up_7_1),                          
/* output logic              [23:0] */ .dqring_out_up_0_0          (mpp_dqring_out_0_0),                         
/* output logic              [23:0] */ .dqring_out_up_0_1          (mpp_dqring_out_0_1),                         
/* output logic              [23:0] */ .dqring_out_up_1_0          (mpp_dqring_out_1_0),                         
/* output logic              [23:0] */ .dqring_out_up_1_1          (mpp_dqring_out_1_1),                         
/* output logic              [23:0] */ .dqring_out_up_2_0          (mpp_dqring_out_2_0),                         
/* output logic              [23:0] */ .dqring_out_up_2_1          (mpp_dqring_out_2_1),                         
/* output logic              [23:0] */ .dqring_out_up_3_0          (mpp_dqring_out_3_0),                         
/* output logic              [23:0] */ .dqring_out_up_3_1          (mpp_dqring_out_3_1),                         
/* output logic              [23:0] */ .dqring_out_up_4_0          (mpp_dqring_out_4_0),                         
/* output logic              [23:0] */ .dqring_out_up_4_1          (mpp_dqring_out_4_1),                         
/* output logic              [23:0] */ .dqring_out_up_5_0          (mpp_dqring_out_5_0),                         
/* output logic              [23:0] */ .dqring_out_up_5_1          (mpp_dqring_out_5_1),                         
/* output logic              [23:0] */ .dqring_out_up_6_0          (mpp_dqring_out_6_0),                         
/* output logic              [23:0] */ .dqring_out_up_6_1          (mpp_dqring_out_6_1),                         
/* output logic              [23:0] */ .dqring_out_up_7_0          (mpp_dqring_out_7_0),                         
/* output logic              [23:0] */ .dqring_out_up_7_1          (mpp_dqring_out_7_1),                         
/* output logic              [25:0] */ .gpolring_out_dn_0_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_0_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_1_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_1_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_2_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_2_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_3_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_3_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_4_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_4_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_5_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_5_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_6_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_6_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_7_0        (),                                           
/* output logic              [25:0] */ .gpolring_out_dn_7_1        (),                                           
/* output logic              [25:0] */ .gpolring_out_up_0_0        (mpp_gpolring_out_0_0),                       
/* output logic              [25:0] */ .gpolring_out_up_0_1        (mpp_gpolring_out_0_1),                       
/* output logic              [25:0] */ .gpolring_out_up_1_0        (mpp_gpolring_out_1_0),                       
/* output logic              [25:0] */ .gpolring_out_up_1_1        (mpp_gpolring_out_1_1),                       
/* output logic              [25:0] */ .gpolring_out_up_2_0        (mpp_gpolring_out_2_0),                       
/* output logic              [25:0] */ .gpolring_out_up_2_1        (mpp_gpolring_out_2_1),                       
/* output logic              [25:0] */ .gpolring_out_up_3_0        (mpp_gpolring_out_3_0),                       
/* output logic              [25:0] */ .gpolring_out_up_3_1        (mpp_gpolring_out_3_1),                       
/* output logic              [25:0] */ .gpolring_out_up_4_0        (mpp_gpolring_out_4_0),                       
/* output logic              [25:0] */ .gpolring_out_up_4_1        (mpp_gpolring_out_4_1),                       
/* output logic              [25:0] */ .gpolring_out_up_5_0        (mpp_gpolring_out_5_0),                       
/* output logic              [25:0] */ .gpolring_out_up_5_1        (mpp_gpolring_out_5_1),                       
/* output logic              [25:0] */ .gpolring_out_up_6_0        (mpp_gpolring_out_6_0),                       
/* output logic              [25:0] */ .gpolring_out_up_6_1        (mpp_gpolring_out_6_1),                       
/* output logic              [25:0] */ .gpolring_out_up_7_0        (mpp_gpolring_out_7_0),                       
/* output logic              [25:0] */ .gpolring_out_up_7_1        (mpp_gpolring_out_7_1),                       
/* output logic             [106:0] */ .gpolring_update_out_dn_0   (),                                           
/* output logic             [106:0] */ .gpolring_update_out_dn_1   (),                                           
/* output logic             [106:0] */ .gpolring_update_out_up_0   (mpp_gpolring_update_out_0),                  
/* output logic             [106:0] */ .gpolring_update_out_up_1   (mpp_gpolring_update_out_1),                  
/* output logic                     */ .grp_a_tx_pfc_tc_sync       (grp_a1_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_a_tx_pfc_xoff          (grp_a1_tx_pfc_xoff),                         
/* output logic                     */ .grp_b_tx_pfc_tc_sync       (grp_b1_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_b_tx_pfc_xoff          (grp_b1_tx_pfc_xoff),                         
/* output logic                     */ .grp_c_tx_pfc_tc_sync       (grp_c1_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_c_tx_pfc_xoff          (grp_c1_tx_pfc_xoff),                         
/* output logic                     */ .grp_d_tx_pfc_tc_sync       (grp_d1_tx_pfc_tc_sync),                      
/* output logic               [3:0] */ .grp_d_tx_pfc_xoff          (grp_d1_tx_pfc_xoff),                         
/* output logic                     */ .igr_vp_tx_pfc_xoff         (igr1_vp_tx_pfc_xoff),                        //FIXME should this be [1:0] for 2 VP   
/* output logic              [68:0] */ .mctagring_out_dn_0         (mgp_mctagring_up_0),                         
/* output logic              [68:0] */ .mctagring_out_dn_1         (mgp_mctagring_up_1),                         
/* output logic              [68:0] */ .mctagring_out_dn_2         (mgp_mctagring_up_2),                         
/* output logic              [68:0] */ .mctagring_out_dn_3         (mgp_mctagring_up_3),                         
/* output logic              [68:0] */ .mctagring_out_up_0         (),                                           
/* output logic              [68:0] */ .mctagring_out_up_1         (),                                           
/* output logic              [68:0] */ .mctagring_out_up_2         (),                                           
/* output logic              [68:0] */ .mctagring_out_up_3         (),                                           
/* output logic              [33:0] */ .mrpodring_out_dn           (mgp_mrpodring_up),                           
/* output logic              [33:0] */ .mrpodring_out_up           (mpp_mrpodring_out_dn),                       
/* output logic                     */ .mrpodring_stall_out_dn     (mgp_mrpodring_stall_up),                     
/* output logic                     */ .mrpodring_stall_out_up     (mpp_mrpodring_stall_out_dn),                 
/* output logic              [33:0] */ .podring_out_dn             (mgp_podring_up),                             
/* output logic              [33:0] */ .podring_out_up             (mpp_podring_out_dn),                         
/* output logic                     */ .podring_stall_out_dn       (mgp_podring_stall_up),                       
/* output logic                     */ .podring_stall_out_up       (mpp_podring_stall_out_dn),                   
/* output logic              [67:0] */ .tagring_out_dn_0_0         (mgp_tagring_up_0_0),                         
/* output logic              [67:0] */ .tagring_out_dn_0_1         (mgp_tagring_up_0_1),                         
/* output logic              [67:0] */ .tagring_out_dn_10_0        (mgp_tagring_up_10_0),                        
/* output logic              [67:0] */ .tagring_out_dn_10_1        (mgp_tagring_up_10_1),                        
/* output logic              [67:0] */ .tagring_out_dn_11_0        (mgp_tagring_up_11_0),                        
/* output logic              [67:0] */ .tagring_out_dn_11_1        (mgp_tagring_up_11_1),                        
/* output logic              [67:0] */ .tagring_out_dn_12_0        (mgp_tagring_up_12_0),                        
/* output logic              [67:0] */ .tagring_out_dn_12_1        (mgp_tagring_up_12_1),                        
/* output logic              [67:0] */ .tagring_out_dn_13_0        (mgp_tagring_up_13_0),                        
/* output logic              [67:0] */ .tagring_out_dn_13_1        (mgp_tagring_up_13_1),                        
/* output logic              [67:0] */ .tagring_out_dn_14_0        (mgp_tagring_up_14_0),                        
/* output logic              [67:0] */ .tagring_out_dn_14_1        (mgp_tagring_up_14_1),                        
/* output logic              [67:0] */ .tagring_out_dn_15_0        (mgp_tagring_up_15_0),                        
/* output logic              [67:0] */ .tagring_out_dn_15_1        (mgp_tagring_up_15_1),                        
/* output logic              [67:0] */ .tagring_out_dn_1_0         (mgp_tagring_up_1_0),                         
/* output logic              [67:0] */ .tagring_out_dn_1_1         (mgp_tagring_up_1_1),                         
/* output logic              [67:0] */ .tagring_out_dn_2_0         (mgp_tagring_up_2_0),                         
/* output logic              [67:0] */ .tagring_out_dn_2_1         (mgp_tagring_up_2_1),                         
/* output logic              [67:0] */ .tagring_out_dn_3_0         (mgp_tagring_up_3_0),                         
/* output logic              [67:0] */ .tagring_out_dn_3_1         (mgp_tagring_up_3_1),                         
/* output logic              [67:0] */ .tagring_out_dn_4_0         (mgp_tagring_up_4_0),                         
/* output logic              [67:0] */ .tagring_out_dn_4_1         (mgp_tagring_up_4_1),                         
/* output logic              [67:0] */ .tagring_out_dn_5_0         (mgp_tagring_up_5_0),                         
/* output logic              [67:0] */ .tagring_out_dn_5_1         (mgp_tagring_up_5_1),                         
/* output logic              [67:0] */ .tagring_out_dn_6_0         (mgp_tagring_up_6_0),                         
/* output logic              [67:0] */ .tagring_out_dn_6_1         (mgp_tagring_up_6_1),                         
/* output logic              [67:0] */ .tagring_out_dn_7_0         (mgp_tagring_up_7_0),                         
/* output logic              [67:0] */ .tagring_out_dn_7_1         (mgp_tagring_up_7_1),                         
/* output logic              [67:0] */ .tagring_out_dn_8_0         (mgp_tagring_up_8_0),                         
/* output logic              [67:0] */ .tagring_out_dn_8_1         (mgp_tagring_up_8_1),                         
/* output logic              [67:0] */ .tagring_out_dn_9_0         (mgp_tagring_up_9_0),                         
/* output logic              [67:0] */ .tagring_out_dn_9_1         (mgp_tagring_up_9_1),                         
/* output logic              [67:0] */ .tagring_out_up_0_0         (mpp_tagring_out_dn_0_0),                     
/* output logic              [67:0] */ .tagring_out_up_0_1         (mpp_tagring_out_dn_0_1),                     
/* output logic              [67:0] */ .tagring_out_up_10_0        (mpp_tagring_out_dn_10_0),                    
/* output logic              [67:0] */ .tagring_out_up_10_1        (mpp_tagring_out_dn_10_1),                    
/* output logic              [67:0] */ .tagring_out_up_11_0        (mpp_tagring_out_dn_11_0),                    
/* output logic              [67:0] */ .tagring_out_up_11_1        (mpp_tagring_out_dn_11_1),                    
/* output logic              [67:0] */ .tagring_out_up_12_0        (mpp_tagring_out_dn_12_0),                    
/* output logic              [67:0] */ .tagring_out_up_12_1        (mpp_tagring_out_dn_12_1),                    
/* output logic              [67:0] */ .tagring_out_up_13_0        (mpp_tagring_out_dn_13_0),                    
/* output logic              [67:0] */ .tagring_out_up_13_1        (mpp_tagring_out_dn_13_1),                    
/* output logic              [67:0] */ .tagring_out_up_14_0        (mpp_tagring_out_dn_14_0),                    
/* output logic              [67:0] */ .tagring_out_up_14_1        (mpp_tagring_out_dn_14_1),                    
/* output logic              [67:0] */ .tagring_out_up_15_0        (mpp_tagring_out_dn_15_0),                    
/* output logic              [67:0] */ .tagring_out_up_15_1        (mpp_tagring_out_dn_15_1),                    
/* output logic              [67:0] */ .tagring_out_up_1_0         (mpp_tagring_out_dn_1_0),                     
/* output logic              [67:0] */ .tagring_out_up_1_1         (mpp_tagring_out_dn_1_1),                     
/* output logic              [67:0] */ .tagring_out_up_2_0         (mpp_tagring_out_dn_2_0),                     
/* output logic              [67:0] */ .tagring_out_up_2_1         (mpp_tagring_out_dn_2_1),                     
/* output logic              [67:0] */ .tagring_out_up_3_0         (mpp_tagring_out_dn_3_0),                     
/* output logic              [67:0] */ .tagring_out_up_3_1         (mpp_tagring_out_dn_3_1),                     
/* output logic              [67:0] */ .tagring_out_up_4_0         (mpp_tagring_out_dn_4_0),                     
/* output logic              [67:0] */ .tagring_out_up_4_1         (mpp_tagring_out_dn_4_1),                     
/* output logic              [67:0] */ .tagring_out_up_5_0         (mpp_tagring_out_dn_5_0),                     
/* output logic              [67:0] */ .tagring_out_up_5_1         (mpp_tagring_out_dn_5_1),                     
/* output logic              [67:0] */ .tagring_out_up_6_0         (mpp_tagring_out_dn_6_0),                     
/* output logic              [67:0] */ .tagring_out_up_6_1         (mpp_tagring_out_dn_6_1),                     
/* output logic              [67:0] */ .tagring_out_up_7_0         (mpp_tagring_out_dn_7_0),                     
/* output logic              [67:0] */ .tagring_out_up_7_1         (mpp_tagring_out_dn_7_1),                     
/* output logic              [67:0] */ .tagring_out_up_8_0         (mpp_tagring_out_dn_8_0),                     
/* output logic              [67:0] */ .tagring_out_up_8_1         (mpp_tagring_out_dn_8_1),                     
/* output logic              [67:0] */ .tagring_out_up_9_0         (mpp_tagring_out_dn_9_0),                     
/* output logic              [67:0] */ .tagring_out_up_9_1         (mpp_tagring_out_dn_9_1));                     
// End of module mgp1 from mby_mgp


// module ppestm    from ppe_stm_top using ppestm.map 
ppe_stm_top    ppestm(
/* input  logic                       */ .cclk                       (cclk),                                       
/* input  logic                [98:0] */ .i_ibus_ctrl                (),                                           
/* input  logic                       */ .reset                      (sreset),                                     
/* Interface egr_ppe_stm_if.stm       */ .egr_ppe_stm_if0            (egr0_ppestm),                                
/* Interface egr_ppe_stm_if.stm       */ .egr_ppe_stm_if1            (egr1_ppestm),                                
/* Interface egr_mc_table_if.mc_table */ .mc_table_if0_0             (egr0_mc_table0),                             
/* Interface egr_mc_table_if.mc_table */ .mc_table_if0_1             (egr0_mc_table1),                             
/* Interface egr_mc_table_if.mc_table */ .mc_table_if1_0             (egr1_mc_table0),                             
/* Interface egr_mc_table_if.mc_table */ .mc_table_if1_1             (egr1_mc_table1),                             
/* Interface rx_ppe_ppe_stm0_if.stm   */ .rx_ppe_ppe_stm0_if0        (rxppe0_ppestm0),                             
/* Interface rx_ppe_ppe_stm0_if.stm   */ .rx_ppe_ppe_stm0_if1        (rxppe1_ppestm0),                             
/* Interface rx_ppe_ppe_stm1_if.stm   */ .rx_ppe_ppe_stm1_if0        (rxppe0_ppestm1),                             
/* Interface rx_ppe_ppe_stm1_if.stm   */ .rx_ppe_ppe_stm1_if1        (rxppe1_ppestm1),                             
/* output logic                [66:0] */ .o_ibus_resp                ());                                           
// End of module ppestm from ppe_stm_top



// module mpp_csr_shim    from mby_mpp_csr_shim using mpp_csr_shim.map 
//mby_mpp_csr_shim    mpp_csr_shim(
//* input  logic         */ .cclk                       (cclk),                                       // mby core clock 
//* input  logic         */ .reset                      (sreset),                                     // mby core reset 
//* input  logic  [31:0] */ .i_mpp_csr_start            (i_mpp_csr_start),                            // tied in mpp shell  
//* input  logic  [31:0] */ .i_mpp_csr_end              (i_mpp_csr_end),                              // tied in mpp shell 
//* input  logic         */ .i_reqValid                 (i_reqValid),                                 
//* input  logic  [31:0] */ .i_reqAddr                  (i_reqAddr),                                  
//* input  logic         */ .i_reqWr                    (i_reqWr),                                    // '0'= read 
//* input  logic  [63:0] */ .i_reqWrData                (i_reqWrData),                                
//* input  logic   [7:0] */ .i_reqID                    (i_reqID),                                    // from iMC axi 
//* input  logic         */ .i_reqParity                (i_reqParity),                                // odd parity bit to cover req 
//* input  logic         */ .i_respValid                (respValid),                                  
//* input  logic  [63:0] */ .i_respData                 (respData),                                   
//* input  logic   [7:0] */ .i_respID                   (respID),                                     // same as reqID 
//* input  logic         */ .i_respParity               (respParity),                                 // parity bit to cover neighbor resp 
//* output logic         */ .o_respValid                (respValid),                                  
//* output logic  [63:0] */ .o_respData                 (respData),                                   
//* output logic   [7:0] */ .o_respID                   (respID),                                     
//* output logic         */ .o_respParity               (respParity),                                 
//* input  logic         */ .i_fifoFilled               (fifoFilled),                                 
//* input  logic         */ .i_fifoEmpty                (fifoEmpty),                                  
//* output logic         */ .o_fifoFilled               (fifoFilled),                                 
//* output logic         */ .o_fifoEmpty                (fifoEmpty),                                  
//* output logic         */ .o_reqValid_rTable          (),                                           
//* output logic         */ .o_reqValid_m0              (),                                           
//* output logic         */ .o_reqValid_m1              (),                                           
//* output logic  [24:0] */ .o_reqAddr                  (),                                           
//* output logic         */ .o_reqWr                    (),                                           
//* output logic  [63:0] */ .o_reqWrData                (),                                           
//* input  logic         */ .i_igrAck_m0                (1'b0),                                       
//* input  logic  [63:0] */ .i_igrData_m0               (64'b0),                                      
//* input  logic         */ .i_egrAck_m0                (1'b0),                                       
//* input  logic  [63:0] */ .i_egrData_m0               (64'b0),                                      
//* input  logic         */ .i_rxppeAck_m0              (1'b0),                                       
//* input  logic  [63:0] */ .i_rxppeData_m0             (64'b0),                                      
//* input  logic         */ .i_txppe0Ack_m0             (1'b0),                                       // one mgp has two txppes
//* input  logic  [63:0] */ .i_txppe0Data_m0            (64'b0),                                      
//* input  logic         */ .i_txppe1Ack_m0             (1'b0),                                       
//* input  logic  [63:0] */ .i_txppe1Data_m0            (64'b0),                                      
//* input  logic         */ .i_igrAck_m1                (1'b0),                                       
//* input  logic  [63:0] */ .i_igrData_m1               (64'b0),                                      
//* input  logic         */ .i_egrAck_m1                (1'b0),                                       
//* input  logic  [63:0] */ .i_egrData_m1               (64'b0),                                      
//* input  logic         */ .i_rxppeAck_m1              (1'b0),                                       
//* input  logic  [63:0] */ .i_rxppeData_m1             (64'b0),                                      
//* input  logic         */ .i_txppe0Ack_m1             (1'b0),                                       // one mgp has two txppes
//* input  logic  [63:0] */ .i_txppe0Data_m1            (64'b0),                                      
//* input  logic         */ .i_txppe1Ack_m1             (1'b0),                                       
//* input  logic  [63:0] */ .i_txppe1Data_m1            (64'b0),                                      
//* input  logic         */ .i_rTableAck                (1'b0),                                       // serves as both write ack and read ack
//* input  logic  [63:0] */ .i_rTableData               (64'b0));                                      
// End of module mpp_csr_shim from mby_mpp_csr_shim


// collage-pragma translate_on

endmodule // mby_mpp
