magic
tech scmos
timestamp 965420547
<< ndiffusion >>
rect -33 70 -21 71
rect 1 70 9 71
rect -33 62 -21 67
rect -33 58 -21 59
rect -33 50 -31 58
rect -33 49 -21 50
rect 1 62 9 67
rect 1 58 9 59
rect 1 49 9 50
rect -33 41 -21 46
rect 1 41 9 46
rect -33 37 -21 38
rect -33 29 -31 37
rect -23 29 -21 37
rect 1 37 9 38
rect -33 28 -21 29
rect 1 28 9 29
rect -33 22 -21 25
rect -31 18 -21 22
rect 1 20 9 25
rect 1 16 9 17
rect 1 7 9 8
rect 1 -1 9 4
rect 1 -5 9 -4
<< pdiffusion >>
rect 25 70 33 71
rect 54 70 72 71
rect 25 62 33 67
rect 54 62 72 67
rect 25 58 33 59
rect 25 49 33 50
rect 25 41 33 46
rect 54 58 72 59
rect 70 50 72 58
rect 54 49 72 50
rect 54 41 72 46
rect 25 37 33 38
rect 25 28 33 29
rect 54 37 72 38
rect 70 29 72 37
rect 54 28 72 29
rect 25 20 33 25
rect 25 16 33 17
rect 25 7 33 8
rect 54 24 72 25
rect 54 19 64 24
rect 25 -1 33 4
rect 25 -5 33 -4
<< ntransistor >>
rect -33 67 -21 70
rect 1 67 9 70
rect -33 59 -21 62
rect 1 59 9 62
rect -33 46 -21 49
rect 1 46 9 49
rect -33 38 -21 41
rect 1 38 9 41
rect -33 25 -21 28
rect 1 25 9 28
rect 1 17 9 20
rect 1 4 9 7
rect 1 -4 9 -1
<< ptransistor >>
rect 25 67 33 70
rect 54 67 72 70
rect 25 59 33 62
rect 54 59 72 62
rect 25 46 33 49
rect 54 46 72 49
rect 25 38 33 41
rect 54 38 72 41
rect 25 25 33 28
rect 54 25 72 28
rect 25 17 33 20
rect 25 4 33 7
rect 25 -4 33 -1
<< polysilicon >>
rect -37 67 -33 70
rect -21 67 1 70
rect 9 67 25 70
rect 33 67 54 70
rect 72 67 76 70
rect -35 59 -33 62
rect -21 59 -16 62
rect -38 49 -35 54
rect -11 54 -8 67
rect -3 59 1 62
rect 9 59 25 62
rect 33 59 45 62
rect 50 59 54 62
rect 72 59 74 62
rect -38 46 -33 49
rect -21 46 -16 49
rect -3 46 1 49
rect 9 46 25 49
rect 33 46 37 49
rect 42 41 45 59
rect 74 49 77 54
rect 50 46 54 49
rect 72 46 77 49
rect -37 38 -33 41
rect -21 38 1 41
rect 9 38 25 41
rect 33 38 54 41
rect 72 38 76 41
rect -37 25 -33 28
rect -21 25 -19 28
rect 37 33 45 38
rect -3 25 1 28
rect 9 25 25 28
rect 33 25 37 28
rect 50 25 54 28
rect 72 25 77 28
rect -3 17 1 20
rect 9 17 25 20
rect 33 17 37 20
rect -11 -1 -8 12
rect 42 7 45 25
rect 74 12 77 25
rect -3 4 1 7
rect 9 4 25 7
rect 33 4 45 7
rect -11 -4 1 -1
rect 9 -4 25 -1
rect 33 -4 37 -1
<< ndcontact >>
rect -33 71 -21 79
rect 1 71 9 79
rect -31 50 -21 58
rect 1 50 9 58
rect -31 29 -23 37
rect 1 29 9 37
rect -39 14 -31 22
rect 1 8 9 16
rect 1 -13 9 -5
<< pdcontact >>
rect 25 71 33 79
rect 54 71 72 79
rect 25 50 33 58
rect 54 50 70 58
rect 25 29 33 37
rect 54 29 70 37
rect 25 8 33 16
rect 64 16 72 24
rect 25 -13 33 -5
<< polycontact >>
rect -43 54 -35 62
rect -11 46 -3 54
rect 74 54 82 62
rect -19 25 -11 33
rect 37 25 45 33
rect -11 12 -3 20
rect 69 4 77 12
<< metal1 >>
rect -33 71 9 79
rect 25 71 72 79
rect -39 62 78 66
rect -43 54 -35 62
rect -39 22 -35 54
rect -31 54 -21 58
rect -31 50 -15 54
rect -31 29 -23 37
rect -39 14 -31 22
rect -27 -5 -23 29
rect -19 33 -15 50
rect -11 46 -3 54
rect 1 50 70 58
rect 74 54 82 62
rect -19 25 -11 33
rect -19 8 -15 25
rect -7 20 -3 46
rect 1 29 9 37
rect -11 12 -3 20
rect 13 16 21 50
rect 29 37 58 41
rect 25 29 33 37
rect 37 25 45 33
rect 54 29 70 37
rect 74 24 78 54
rect 64 17 78 24
rect 64 16 72 17
rect 1 12 33 16
rect 1 8 77 12
rect -19 4 5 8
rect 27 6 77 8
rect 69 4 77 6
rect -27 -13 9 -5
rect 25 -13 33 -5
<< labels >>
rlabel metal1 5 54 5 54 1 x
rlabel metal1 5 75 5 75 5 GND!
rlabel metal1 29 54 29 54 1 x
rlabel metal1 29 75 29 75 5 Vdd!
rlabel metal1 29 33 29 33 1 Vdd!
rlabel metal1 5 12 5 12 1 x
rlabel metal1 29 12 29 12 1 x
rlabel metal1 5 -9 5 -9 1 GND!
rlabel metal1 29 -9 29 -9 1 Vdd!
rlabel metal1 5 33 5 33 1 GND!
rlabel metal1 63 75 63 75 5 Vdd!
rlabel metal1 62 54 62 54 5 x
rlabel metal1 62 33 62 33 1 Vdd!
rlabel metal1 41 29 41 29 1 b
rlabel space -43 -14 8 80 7 ^n
rlabel space 26 -15 83 80 3 ^p
rlabel metal1 -7 16 -7 16 1 a
rlabel metal1 -7 50 -7 50 1 a
rlabel metal1 -26 54 -26 54 1 x
rlabel metal1 -27 75 -27 75 5 GND!
rlabel metal1 -27 33 -27 33 1 GND!
rlabel metal1 73 8 73 8 1 x
<< end >>
