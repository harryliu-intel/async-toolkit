magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 11 59 15 60
rect 11 53 15 57
rect 29 53 33 54
rect 11 47 15 51
rect -3 39 1 44
rect 11 44 15 45
rect 11 39 15 40
rect 29 47 33 51
rect 29 44 33 45
rect 29 39 33 40
rect -3 34 1 37
rect 11 33 15 37
rect 29 33 33 37
rect 11 27 15 31
rect 29 30 33 31
rect 11 24 15 25
<< pdiffusion >>
rect 45 53 49 54
rect 63 53 69 54
rect 78 53 90 54
rect 45 47 49 51
rect 63 47 69 51
rect 78 50 90 51
rect 78 47 86 50
rect 45 44 49 45
rect 45 39 49 40
rect 45 33 49 37
rect 63 44 69 45
rect 67 40 69 44
rect 63 39 69 40
rect 82 39 85 42
rect 63 33 69 37
rect 79 35 85 39
rect 45 30 49 31
rect 63 30 69 31
rect 79 30 85 33
<< ntransistor >>
rect 11 57 15 59
rect 11 51 15 53
rect 29 51 33 53
rect 11 45 15 47
rect 29 45 33 47
rect -3 37 1 39
rect 11 37 15 39
rect 29 37 33 39
rect 11 31 15 33
rect 29 31 33 33
rect 11 25 15 27
<< ptransistor >>
rect 45 51 49 53
rect 63 51 69 53
rect 78 51 90 53
rect 45 45 49 47
rect 63 45 69 47
rect 45 37 49 39
rect 63 37 69 39
rect 79 33 85 35
rect 45 31 49 33
rect 63 31 69 33
<< polysilicon >>
rect 8 57 11 59
rect 15 57 18 59
rect 8 51 11 53
rect 15 51 29 53
rect 33 51 45 53
rect 49 51 63 53
rect 69 51 72 53
rect 75 51 78 53
rect 90 51 93 53
rect 8 45 11 47
rect 15 45 18 47
rect 8 43 9 45
rect 7 39 9 43
rect 21 39 23 51
rect 26 45 29 47
rect 33 45 45 47
rect 49 45 57 47
rect 60 45 63 47
rect 69 45 73 47
rect -5 37 -3 39
rect 1 37 4 39
rect 7 37 11 39
rect 15 37 18 39
rect 21 37 29 39
rect 33 37 45 39
rect 49 37 52 39
rect 55 33 57 45
rect 71 43 73 45
rect 60 37 63 39
rect 69 37 73 39
rect 76 33 79 35
rect 85 33 87 35
rect 8 31 11 33
rect 15 31 29 33
rect 33 31 45 33
rect 49 31 63 33
rect 69 31 72 33
rect 8 25 11 27
rect 15 25 18 27
<< ndcontact >>
rect 11 60 15 64
rect 29 54 33 58
rect -3 44 1 48
rect 11 40 15 44
rect 29 40 33 44
rect -3 30 1 34
rect 29 26 33 30
rect 11 20 15 24
<< pdcontact >>
rect 45 54 49 58
rect 63 54 69 58
rect 78 54 90 58
rect 86 46 90 50
rect 45 40 49 44
rect 63 40 67 44
rect 78 39 82 43
rect 45 26 49 30
rect 63 26 69 30
rect 79 26 85 30
<< polycontact >>
rect -9 37 -5 41
rect 4 43 8 47
rect 71 39 75 43
rect 87 33 91 37
<< metal1 >>
rect 11 58 15 64
rect 11 54 33 58
rect 45 54 90 58
rect -3 47 1 48
rect 5 47 74 50
rect -3 44 8 47
rect 4 43 8 44
rect -9 40 -5 41
rect 11 40 67 44
rect -9 37 15 40
rect 63 36 67 40
rect 71 43 74 47
rect 86 46 90 50
rect 71 39 82 43
rect 87 37 90 46
rect 87 36 91 37
rect -3 30 1 34
rect 63 33 91 36
rect -3 26 33 30
rect 45 26 85 30
rect 11 20 15 26
<< labels >>
rlabel polysilicon 70 52 70 52 1 b
rlabel polysilicon 70 32 70 32 1 a
rlabel polysilicon 10 52 10 52 3 b
rlabel polysilicon 10 32 10 32 1 a
rlabel polysilicon 10 58 10 58 1 _SReset!
rlabel polysilicon 10 26 10 26 1 _SReset!
rlabel polysilicon 91 52 91 52 1 _PReset!
rlabel space 48 25 94 59 3 ^p
rlabel space -10 19 30 65 7 ^n
rlabel pdcontact 65 42 65 42 1 x
rlabel pdcontact 66 28 66 28 1 Vdd!
rlabel pdcontact 66 56 66 56 1 Vdd!
rlabel ndcontact 31 42 31 42 1 x
rlabel pdcontact 47 42 47 42 1 x
rlabel pdcontact 47 28 47 28 1 Vdd!
rlabel pdcontact 47 56 47 56 1 Vdd!
rlabel ndcontact 13 62 13 62 5 GND!
rlabel ndcontact 13 22 13 22 1 GND!
rlabel pdcontact 84 56 84 56 5 Vdd!
rlabel pdcontact 88 48 88 48 7 x
rlabel ndcontact 31 56 31 56 5 GND!
rlabel ndcontact 31 28 31 28 1 GND!
rlabel ndcontact 13 42 13 42 1 x
rlabel ndcontact -1 32 -1 32 1 GND!
rlabel polycontact -7 39 -7 39 3 x
rlabel pdcontact 82 28 82 28 3 Vdd!
rlabel polycontact 89 35 89 35 7 x
<< end >>
