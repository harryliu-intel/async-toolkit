magic
tech scmos
timestamp 982685480
<< nselect >>
rect -60 -815 0 -691
<< pselect >>
rect 0 -837 73 -668
<< ndiffusion >>
rect -28 -705 -8 -704
rect -28 -713 -8 -708
rect -28 -721 -8 -716
rect -28 -729 -8 -724
rect -28 -737 -8 -732
rect -28 -745 -8 -740
rect -28 -749 -8 -748
rect -28 -758 -8 -757
rect -28 -766 -8 -761
rect -28 -774 -8 -769
rect -28 -782 -8 -777
rect -28 -790 -8 -785
rect -28 -798 -8 -793
rect -28 -802 -8 -801
<< pdiffusion >>
rect 15 -680 41 -679
rect 15 -684 41 -683
rect 28 -692 41 -684
rect 15 -693 41 -692
rect 15 -697 41 -696
rect 15 -706 41 -705
rect 15 -710 41 -709
rect 28 -718 41 -710
rect 15 -719 41 -718
rect 15 -723 41 -722
rect 15 -732 41 -731
rect 15 -736 41 -735
rect 28 -744 41 -736
rect 15 -745 41 -744
rect 15 -749 41 -748
rect 15 -758 41 -757
rect 15 -762 41 -761
rect 28 -770 41 -762
rect 15 -771 41 -770
rect 15 -775 41 -774
rect 15 -784 41 -783
rect 15 -788 41 -787
rect 28 -796 41 -788
rect 15 -797 41 -796
rect 15 -801 41 -800
rect 15 -810 41 -809
rect 15 -814 41 -813
rect 28 -822 41 -814
rect 15 -823 41 -822
rect 15 -827 41 -826
<< ntransistor >>
rect -28 -708 -8 -705
rect -28 -716 -8 -713
rect -28 -724 -8 -721
rect -28 -732 -8 -729
rect -28 -740 -8 -737
rect -28 -748 -8 -745
rect -28 -761 -8 -758
rect -28 -769 -8 -766
rect -28 -777 -8 -774
rect -28 -785 -8 -782
rect -28 -793 -8 -790
rect -28 -801 -8 -798
<< ptransistor >>
rect 15 -683 41 -680
rect 15 -696 41 -693
rect 15 -709 41 -706
rect 15 -722 41 -719
rect 15 -735 41 -732
rect 15 -748 41 -745
rect 15 -761 41 -758
rect 15 -774 41 -771
rect 15 -787 41 -784
rect 15 -800 41 -797
rect 15 -813 41 -810
rect 15 -826 41 -823
<< polysilicon >>
rect -6 -683 15 -680
rect 41 -683 53 -680
rect -6 -705 -3 -683
rect 50 -686 53 -683
rect -32 -708 -28 -705
rect -8 -708 -3 -705
rect 10 -696 15 -693
rect 41 -696 45 -693
rect 10 -706 13 -696
rect 2 -709 15 -706
rect 41 -709 45 -706
rect 2 -713 5 -709
rect -44 -716 -28 -713
rect -8 -716 5 -713
rect 10 -721 15 -719
rect -32 -724 -28 -721
rect -8 -722 15 -721
rect 41 -722 65 -719
rect -8 -724 13 -722
rect -32 -732 -28 -729
rect -8 -732 13 -729
rect 10 -735 15 -732
rect 41 -735 45 -732
rect -52 -740 -28 -737
rect -8 -740 -4 -737
rect -32 -748 -28 -745
rect -8 -748 15 -745
rect 41 -748 45 -745
rect -32 -761 -28 -758
rect -8 -761 15 -758
rect 41 -761 53 -758
rect -40 -769 -28 -766
rect -8 -769 -4 -766
rect 10 -774 15 -771
rect 41 -774 53 -771
rect -32 -777 -28 -774
rect -8 -777 13 -774
rect -32 -785 -28 -782
rect -8 -784 13 -782
rect -8 -785 15 -784
rect 10 -787 15 -785
rect 41 -787 45 -784
rect -48 -793 -28 -790
rect -8 -793 5 -790
rect 2 -797 5 -793
rect -32 -801 -28 -798
rect -8 -801 -3 -798
rect 2 -800 15 -797
rect 41 -800 45 -797
rect -6 -823 -3 -801
rect 10 -810 13 -800
rect 10 -813 15 -810
rect 41 -813 45 -810
rect -6 -826 15 -823
rect 41 -826 45 -823
<< ndcontact >>
rect -28 -704 -8 -696
rect -28 -757 -8 -749
rect -28 -810 -8 -802
<< pdcontact >>
rect 15 -679 41 -671
rect 15 -692 28 -684
rect 15 -705 41 -697
rect 15 -718 28 -710
rect 15 -731 41 -723
rect 15 -744 28 -736
rect 15 -757 41 -749
rect 15 -770 28 -762
rect 15 -783 41 -775
rect 15 -796 28 -788
rect 15 -809 41 -801
rect 15 -822 28 -814
rect 15 -835 41 -827
<< polycontact >>
rect 50 -694 58 -686
rect -52 -721 -44 -713
rect 65 -722 73 -714
rect 45 -735 53 -727
rect -60 -745 -52 -737
rect -40 -753 -32 -745
rect -48 -769 -40 -761
rect 53 -765 61 -757
rect 53 -779 61 -771
rect -56 -793 -48 -785
rect 45 -792 53 -784
rect -40 -806 -32 -798
<< metal1 >>
rect 15 -673 41 -671
rect 27 -679 41 -673
rect -27 -696 -9 -691
rect -4 -692 28 -684
rect -28 -704 -8 -696
rect -4 -710 4 -692
rect 33 -697 41 -679
rect 50 -694 61 -686
rect 15 -705 41 -697
rect -52 -721 -44 -713
rect -60 -745 -52 -737
rect -56 -785 -52 -745
rect -48 -761 -44 -721
rect -4 -718 28 -710
rect -4 -736 4 -718
rect 33 -723 41 -705
rect 15 -724 41 -723
rect 27 -730 41 -724
rect 15 -731 41 -730
rect -4 -744 28 -736
rect -40 -753 -32 -745
rect -4 -749 4 -744
rect 33 -749 41 -731
rect -48 -769 -40 -761
rect -56 -793 -48 -785
rect -36 -798 -32 -753
rect -28 -757 4 -749
rect 15 -757 41 -749
rect -40 -806 -32 -798
rect -4 -762 4 -757
rect -4 -770 28 -762
rect -4 -788 4 -770
rect 33 -775 41 -757
rect 27 -781 41 -775
rect 15 -783 41 -781
rect -4 -796 28 -788
rect -28 -810 -8 -802
rect -27 -817 -9 -810
rect -4 -814 4 -796
rect 33 -801 41 -783
rect 45 -735 53 -727
rect 45 -784 49 -735
rect 57 -757 61 -694
rect 53 -765 61 -757
rect 65 -722 73 -714
rect 65 -771 69 -722
rect 53 -775 69 -771
rect 53 -779 61 -775
rect 45 -792 53 -784
rect 15 -809 41 -801
rect -4 -822 28 -814
rect 33 -827 41 -809
rect 15 -829 41 -827
rect 27 -835 41 -829
<< m2contact >>
rect 9 -679 27 -673
rect -27 -691 -9 -685
rect 9 -730 27 -724
rect 9 -781 27 -775
rect -27 -823 -9 -817
rect 9 -835 27 -829
<< m3contact >>
rect 9 -679 27 -673
rect -27 -691 -9 -685
rect 9 -730 27 -724
rect 9 -781 27 -775
rect -27 -823 -9 -817
rect 9 -835 27 -829
<< metal3 >>
rect -27 -837 -9 -668
rect 9 -837 27 -668
<< labels >>
rlabel metal1 -48 -769 -44 -713 1 e
rlabel metal1 -36 -806 -32 -745 1 a
rlabel metal1 -56 -793 -52 -737 3 b
rlabel space -62 -820 -28 -686 7 ^n
rlabel metal1 45 -792 49 -727 1 c
rlabel metal1 65 -775 69 -714 1 d
rlabel metal1 57 -765 61 -686 1 f
rlabel space 28 -837 74 -668 3 ^p
rlabel metal3 -27 -837 -9 -668 1 GND!|pin|s|0
rlabel metal1 -28 -704 -8 -696 1 GND!|pin|s|0
rlabel metal1 -28 -810 -8 -802 1 GND!|pin|s|0
rlabel metal1 -27 -823 -9 -802 1 GND!|pin|s|0
rlabel metal1 -27 -704 -9 -685 1 GND!|pin|s|0
rlabel metal3 9 -837 27 -668 1 Vdd!|pin|s|1
rlabel metal1 15 -679 41 -671 1 Vdd!|pin|s|1
rlabel metal1 15 -705 41 -697 1 Vdd!|pin|s|1
rlabel metal1 15 -731 41 -723 1 Vdd!|pin|s|1
rlabel metal1 15 -757 41 -749 1 Vdd!|pin|s|1
rlabel metal1 15 -783 41 -775 1 Vdd!|pin|s|1
rlabel metal1 15 -809 41 -801 1 Vdd!|pin|s|1
rlabel metal1 15 -835 41 -827 1 Vdd!|pin|s|1
rlabel metal1 33 -835 41 -671 1 Vdd!|pin|s|1
rlabel metal1 -4 -822 4 -684 1 x|pin|s|2
rlabel metal1 -4 -692 28 -684 1 x|pin|s|2
rlabel metal1 -4 -718 28 -710 1 x|pin|s|2
rlabel metal1 -4 -744 28 -736 1 x|pin|s|2
rlabel metal1 -28 -757 4 -749 1 x|pin|s|2
rlabel metal1 -4 -770 28 -762 1 x|pin|s|2
rlabel metal1 -4 -796 28 -788 1 x|pin|s|2
rlabel metal1 -4 -822 28 -814 1 x|pin|s|2
<< end >>
