magic
tech scmos
timestamp 965071348
<< ndiffusion >>
rect 41 112 49 113
rect 11 96 27 97
rect 41 104 49 109
rect 41 96 49 101
rect 11 88 27 93
rect 41 88 49 93
rect 11 84 27 85
rect 11 76 19 84
rect 11 75 27 76
rect 41 84 49 85
rect 41 75 49 76
rect 11 67 27 72
rect 41 67 49 72
rect 11 63 27 64
rect 41 59 49 64
rect 41 51 49 56
rect 17 41 19 46
rect 41 47 49 48
rect 27 41 33 46
rect 17 40 33 41
rect 17 36 33 37
rect 17 28 19 36
rect 17 27 33 28
rect 17 23 33 24
<< pdiffusion >>
rect 72 127 98 128
rect 103 127 115 128
rect 72 123 98 124
rect 94 115 98 123
rect 72 114 98 115
rect 103 123 115 124
rect 111 115 115 123
rect 103 114 115 115
rect 72 110 98 111
rect 72 102 80 110
rect 72 101 98 102
rect 103 110 115 111
rect 103 102 107 110
rect 103 101 115 102
rect 72 97 98 98
rect 94 89 98 97
rect 72 88 98 89
rect 103 97 115 98
rect 111 89 115 97
rect 103 88 115 89
rect 72 84 98 85
rect 94 76 98 84
rect 72 75 98 76
rect 103 84 115 85
rect 103 76 107 84
rect 103 75 115 76
rect 72 71 98 72
rect 94 63 98 71
rect 72 62 98 63
rect 103 71 115 72
rect 111 63 115 71
rect 103 62 115 63
rect 72 58 98 59
rect 72 50 80 58
rect 72 49 98 50
rect 103 58 115 59
rect 103 50 107 58
rect 103 49 115 50
rect 72 45 98 46
rect 94 37 98 45
rect 72 36 98 37
rect 103 45 115 46
rect 111 37 115 45
rect 103 36 115 37
rect 72 32 98 33
rect 72 30 82 32
rect 65 25 82 30
rect 65 22 77 25
rect 103 32 115 33
rect 103 24 107 32
rect 103 22 115 24
rect 65 18 77 19
rect 103 18 115 19
<< ntransistor >>
rect 41 109 49 112
rect 41 101 49 104
rect 11 93 27 96
rect 41 93 49 96
rect 11 85 27 88
rect 41 85 49 88
rect 11 72 27 75
rect 41 72 49 75
rect 11 64 27 67
rect 41 64 49 67
rect 41 56 49 59
rect 41 48 49 51
rect 17 37 33 40
rect 17 24 33 27
<< ptransistor >>
rect 72 124 98 127
rect 103 124 115 127
rect 72 111 98 114
rect 103 111 115 114
rect 72 98 98 101
rect 103 98 115 101
rect 72 85 98 88
rect 103 85 115 88
rect 72 72 98 75
rect 103 72 115 75
rect 72 59 98 62
rect 103 59 115 62
rect 72 46 98 49
rect 103 46 115 49
rect 72 33 98 36
rect 103 33 115 36
rect 65 19 77 22
rect 103 19 115 22
<< polysilicon >>
rect 51 124 72 127
rect 98 124 103 127
rect 115 124 119 127
rect 51 112 54 124
rect 29 109 41 112
rect 49 109 54 112
rect 59 111 72 114
rect 98 111 103 114
rect 115 111 119 114
rect 29 96 32 109
rect 59 104 62 111
rect 37 101 41 104
rect 49 101 62 104
rect 67 98 72 101
rect 98 98 103 101
rect 115 98 119 101
rect 67 96 70 98
rect 7 93 11 96
rect 27 93 32 96
rect 37 93 41 96
rect 49 93 70 96
rect 7 85 11 88
rect 27 85 41 88
rect 49 85 72 88
rect 98 85 103 88
rect 115 85 119 88
rect 7 72 11 75
rect 27 72 41 75
rect 49 72 72 75
rect 98 72 103 75
rect 115 72 119 75
rect 7 64 11 67
rect 27 64 32 67
rect 37 64 41 67
rect 49 64 70 67
rect 29 51 32 64
rect 67 62 70 64
rect 67 59 72 62
rect 98 59 103 62
rect 115 59 119 62
rect 37 56 41 59
rect 49 56 62 59
rect 29 48 41 51
rect 49 48 54 51
rect 15 37 17 40
rect 33 37 37 40
rect 51 36 54 48
rect 59 49 62 56
rect 59 46 72 49
rect 98 46 103 49
rect 115 46 119 49
rect 51 33 72 36
rect 98 33 103 36
rect 115 33 119 36
rect 13 24 17 27
rect 33 24 53 27
rect 61 19 65 22
rect 77 19 81 22
rect 91 20 103 22
rect 94 19 103 20
rect 115 19 119 22
<< ndcontact >>
rect 41 113 49 121
rect 11 97 27 105
rect 19 76 27 84
rect 41 76 49 84
rect 11 55 27 63
rect 19 41 27 49
rect 41 39 49 47
rect 19 28 33 36
rect 17 15 33 23
<< pdcontact >>
rect 72 128 98 136
rect 103 128 115 136
rect 72 115 94 123
rect 103 115 111 123
rect 80 102 98 110
rect 107 102 115 110
rect 72 89 94 97
rect 103 89 111 97
rect 72 76 94 84
rect 107 76 115 84
rect 72 63 94 71
rect 103 63 111 71
rect 80 50 98 58
rect 107 50 115 58
rect 72 37 94 45
rect 103 37 111 45
rect 82 24 98 32
rect 107 24 115 32
rect 65 10 77 18
rect 103 10 115 18
<< polycontact >>
rect 7 32 15 40
rect 53 19 61 27
rect 86 12 94 20
<< metal1 >>
rect 72 128 98 136
rect 103 132 115 136
rect 103 128 119 132
rect 41 113 49 121
rect 72 115 94 123
rect 103 119 111 123
rect 98 115 111 119
rect 11 97 27 105
rect 72 97 76 115
rect 98 110 103 115
rect 115 110 119 128
rect 80 102 103 110
rect 107 102 119 110
rect 98 97 103 102
rect 11 63 15 97
rect 72 89 94 97
rect 98 89 111 97
rect 19 76 63 84
rect 72 76 94 84
rect 11 55 27 63
rect 19 41 27 55
rect 55 58 63 76
rect 98 71 103 89
rect 115 84 119 102
rect 107 76 119 84
rect 72 63 94 71
rect 98 63 111 71
rect 7 32 15 40
rect 41 36 49 47
rect 11 23 15 32
rect 19 28 49 36
rect 55 27 61 50
rect 72 45 76 63
rect 98 58 103 63
rect 115 58 119 76
rect 88 50 103 58
rect 107 50 119 58
rect 98 45 103 50
rect 72 37 94 45
rect 98 41 111 45
rect 103 37 111 41
rect 115 32 119 50
rect 11 19 33 23
rect 53 19 61 27
rect 82 24 103 32
rect 107 28 119 32
rect 107 24 115 28
rect 17 15 49 19
rect 65 17 77 18
rect 86 17 94 20
rect 65 15 94 17
rect 45 12 94 15
rect 98 18 103 24
rect 45 11 77 12
rect 65 10 77 11
rect 98 10 115 18
<< m2contact >>
rect 55 50 63 58
rect 80 50 88 58
<< metal2 >>
rect 55 50 88 58
<< labels >>
rlabel metal1 76 132 76 132 5 Vdd!
rlabel metal1 76 80 76 80 1 Vdd!
rlabel metal1 45 43 45 43 1 GND!
rlabel metal1 45 117 45 117 5 GND!
rlabel metal1 45 80 45 80 1 x
rlabel metal1 23 80 23 80 1 x
rlabel metal1 111 14 111 14 1 Vdd!
rlabel polysilicon 116 34 116 34 1 _a0
rlabel polysilicon 116 47 116 47 1 _b0
rlabel polysilicon 116 60 116 60 1 _b1
rlabel polysilicon 116 73 116 73 1 _a1
rlabel polysilicon 116 86 116 86 1 _b0
rlabel polysilicon 116 99 116 99 1 _a0
rlabel polysilicon 116 112 116 112 1 _a1
rlabel polysilicon 116 125 116 125 1 _b1
rlabel metal1 90 28 90 28 1 Vdd!
rlabel metal1 26 32 26 32 1 GND!
rlabel m2contact 84 54 84 54 5 x
rlabel metal1 84 106 84 106 1 x
rlabel space 85 9 120 40 3 ^p
rlabel space 89 41 120 137 3 ^p
rlabel space 6 44 42 122 7 ^n
rlabel space 6 14 38 43 7 ^n
<< end >>
