magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect 62 77 70 78
rect 62 69 70 74
rect 62 61 70 66
rect 62 53 70 58
rect 62 49 70 50
rect 62 40 70 41
rect 62 32 70 37
rect 62 24 70 29
rect 62 16 70 21
rect 62 12 70 13
<< pdiffusion >>
rect 86 84 110 85
rect 86 80 110 81
rect 94 75 110 80
rect 86 71 94 72
rect 86 67 94 68
rect 86 58 94 59
rect 86 54 94 55
rect 86 45 94 46
rect 86 41 94 42
rect 86 32 94 33
rect 86 28 94 29
rect 86 19 94 20
rect 86 15 94 16
rect 86 6 94 7
rect 86 2 94 3
<< ntransistor >>
rect 62 74 70 77
rect 62 66 70 69
rect 62 58 70 61
rect 62 50 70 53
rect 62 37 70 40
rect 62 29 70 32
rect 62 21 70 24
rect 62 13 70 16
<< ptransistor >>
rect 86 81 110 84
rect 86 68 94 71
rect 86 55 94 58
rect 86 42 94 45
rect 86 29 94 32
rect 86 16 94 19
rect 86 3 94 6
<< polysilicon >>
rect 82 81 86 84
rect 110 81 114 84
rect 58 74 62 77
rect 70 74 74 77
rect 81 69 86 71
rect 58 66 62 69
rect 70 68 86 69
rect 94 68 98 71
rect 70 66 84 68
rect 58 58 62 61
rect 70 58 84 61
rect 81 55 86 58
rect 94 55 98 58
rect 58 50 62 53
rect 70 50 74 53
rect 81 42 86 45
rect 94 42 98 45
rect 81 40 84 42
rect 58 37 62 40
rect 70 37 84 40
rect 58 29 62 32
rect 70 29 86 32
rect 94 29 98 32
rect 58 21 62 24
rect 70 21 84 24
rect 81 19 84 21
rect 81 16 86 19
rect 94 16 98 19
rect 58 13 62 16
rect 70 13 74 16
rect 81 6 84 16
rect 81 3 86 6
rect 94 3 98 6
<< ndcontact >>
rect 62 78 70 86
rect 62 41 70 49
rect 62 4 70 12
<< pdcontact >>
rect 86 85 110 93
rect 86 72 94 80
rect 86 59 94 67
rect 86 46 94 54
rect 86 33 94 41
rect 86 20 94 28
rect 86 7 94 15
rect 86 -6 94 2
<< metal1 >>
rect 62 78 70 86
rect 74 85 110 93
rect 74 67 82 85
rect 86 72 94 80
rect 74 59 94 67
rect 74 49 82 59
rect 62 41 82 49
rect 86 46 94 54
rect 74 33 94 41
rect 74 15 82 33
rect 86 20 94 28
rect 62 4 70 12
rect 74 7 94 15
rect 86 -6 94 2
<< labels >>
rlabel metal1 90 -2 90 -2 1 Vdd!
rlabel metal1 90 76 90 76 5 Vdd!
rlabel metal1 90 63 90 63 1 x
rlabel metal1 90 50 90 50 5 Vdd!
rlabel metal1 90 37 90 37 5 x
rlabel metal1 90 24 90 24 1 Vdd!
rlabel metal1 90 11 90 11 1 x
rlabel metal1 90 89 90 89 5 x
rlabel polysilicon 61 51 61 51 3 a
rlabel metal1 66 45 66 45 5 x
rlabel polysilicon 61 22 61 22 3 a
rlabel metal1 66 82 66 82 5 GND!
rlabel metal1 66 8 66 8 1 GND!
rlabel polysilicon 61 75 61 75 1 _SReset!
rlabel polysilicon 61 14 61 14 1 _SReset!
rlabel polysilicon 95 56 95 56 3 b
rlabel polysilicon 95 43 95 43 3 c
rlabel polysilicon 95 30 95 30 3 b
rlabel polysilicon 95 69 95 69 3 c
rlabel polysilicon 61 30 61 30 1 b
rlabel polysilicon 61 59 61 59 1 b
rlabel polysilicon 61 67 61 67 1 c
rlabel polysilicon 61 38 61 38 1 c
rlabel polysilicon 95 17 95 17 1 a
rlabel polysilicon 95 4 95 4 1 a
rlabel space 57 4 62 86 7 ^n
rlabel space 94 -6 99 73 3 ^p
rlabel polysilicon 111 82 111 82 7 _PReset!
<< end >>
