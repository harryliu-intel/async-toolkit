magic
tech scmos
timestamp 988943070
use l_c2 l_c2_0
timestamp 988943070
transform 1 0 -1196 0 1 481
box -74 -15 78 82
use l_c2_rhi l_c2_rhi_0
timestamp 988943070
transform 1 0 -974 0 1 580
box -74 -57 78 72
use l_c2_phi l_c2_phi_0
timestamp 988943070
transform 1 0 -730 0 1 471
box -75 40 79 140
use m_c2 m_c2_0
timestamp 988943070
transform 1 0 -1196 0 1 77
box -86 314 94 369
use m_c2_rhi m_c2_rhi_0
timestamp 988943070
transform 1 0 -974 0 1 421
box -88 15 94 86
use s_c2 s_c2_0
timestamp 988943070
transform 1 0 -1196 0 1 58
box -35 283 35 318
use s_c2_rhi s_c2_rhi_0
timestamp 988943070
transform 1 0 -974 0 1 332
box -50 11 62 96
use m_c2_phi m_c2_phi_0
timestamp 988943070
transform 1 0 -730 0 1 605
box -88 -181 94 -110
use m_2and2c2 m_2and2c2_0
timestamp 988943070
transform 1 0 -511 0 1 417
box -77 8 83 139
use m_2and2c2_rhi m_2and2c2_rhi_0
timestamp 988943070
transform 1 0 -299 0 1 432
box -82 29 90 175
use s_c2_phi s_c2_phi_0
timestamp 988943070
transform 1 0 -730 0 1 258
box -50 82 62 155
use s_2and2c2 s_2and2c2_0
timestamp 988943070
transform 1 0 -511 0 1 252
box -61 89 47 154
use s_2and2c2_rhi s_2and2c2_rhi_0
timestamp 988943070
transform 1 0 -299 0 1 318
box -63 23 62 132
use m_and2c2 m_and2c2_0
timestamp 988943070
transform 1 0 -93 0 1 385
box -64 28 79 142
use m_and2c2_rhi m_and2c2_rhi_0
timestamp 988943070
transform 1 0 108 0 1 404
box -72 36 85 163
use s_and2c2 s_and2c2_0
timestamp 988943070
transform 1 0 -93 0 1 -206
box -61 547 47 604
use s_and2c2_rhi s_and2c2_rhi_0
timestamp 988943070
transform 1 0 108 0 1 -164
box -63 505 62 603
<< end >>
