///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cgrp_b_nested_map_pkg.vh                           
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_CGRP_B_NESTED_MAP_PKG_VH
`define MBY_PPE_CGRP_B_NESTED_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_cgrp_b_nested_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_cgrp_b_nested_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_cgrp_b_nested_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_cgrp_b_nested_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [43:0] reserved0;  // RSVD
    logic [19:0] PTR;  // RW
    logic [11:0] reserved1;  // RSVD
    logic  [3:0] SELECT_4;  // RW
    logic  [3:0] SELECT_3;  // RW
    logic  [3:0] SELECT_2;  // RW
    logic  [3:0] SELECT_1;  // RW
    logic  [3:0] SELECT_0;  // RW
    logic [31:0] MASK;  // RW
} EM_HASH_LOOKUP_t;

localparam EM_HASH_LOOKUP_REG_STRIDE = 48'h10;
localparam EM_HASH_LOOKUP_REG_ENTRIES = 8192;
localparam EM_HASH_LOOKUP_CR_ADDR = 48'h0;
localparam EM_HASH_LOOKUP_SIZE = 128;
localparam EM_HASH_LOOKUP_PTR_LO = 64;
localparam EM_HASH_LOOKUP_PTR_HI = 83;
localparam EM_HASH_LOOKUP_PTR_RESET = 20'h0;
localparam EM_HASH_LOOKUP_SELECT_4_LO = 48;
localparam EM_HASH_LOOKUP_SELECT_4_HI = 51;
localparam EM_HASH_LOOKUP_SELECT_4_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_3_LO = 44;
localparam EM_HASH_LOOKUP_SELECT_3_HI = 47;
localparam EM_HASH_LOOKUP_SELECT_3_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_2_LO = 40;
localparam EM_HASH_LOOKUP_SELECT_2_HI = 43;
localparam EM_HASH_LOOKUP_SELECT_2_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_1_LO = 36;
localparam EM_HASH_LOOKUP_SELECT_1_HI = 39;
localparam EM_HASH_LOOKUP_SELECT_1_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_0_LO = 32;
localparam EM_HASH_LOOKUP_SELECT_0_HI = 35;
localparam EM_HASH_LOOKUP_SELECT_0_RESET = 4'h0;
localparam EM_HASH_LOOKUP_MASK_LO = 0;
localparam EM_HASH_LOOKUP_MASK_HI = 31;
localparam EM_HASH_LOOKUP_MASK_RESET = 32'h0;
localparam EM_HASH_LOOKUP_USEMASK = 128'hFFFFF000FFFFFFFFFFFFF;
localparam EM_HASH_LOOKUP_RO_MASK = 128'h0;
localparam EM_HASH_LOOKUP_WO_MASK = 128'h0;
localparam EM_HASH_LOOKUP_RESET = 128'h0;

typedef struct packed {
    logic [23:0] reserved0;  // RSVD
    logic  [7:0] KEY_TOP_INVERT;  // RW
    logic [31:0] KEY_INVERT;  // RW
    logic [23:0] reserved1;  // RSVD
    logic  [7:0] KEY_TOP;  // RW
    logic [31:0] KEY;  // RW
} WCM_TCAM_t;

localparam WCM_TCAM_REG_STRIDE = 48'h10;
localparam WCM_TCAM_REG_ENTRIES = 1024;
localparam WCM_TCAM_REGFILE_STRIDE = 48'h4000;
localparam WCM_TCAM_REGFILE_ENTRIES = 20;
localparam WCM_TCAM_CR_ADDR = 48'h80000;
localparam WCM_TCAM_SIZE = 128;
localparam WCM_TCAM_KEY_TOP_INVERT_LO = 96;
localparam WCM_TCAM_KEY_TOP_INVERT_HI = 103;
localparam WCM_TCAM_KEY_TOP_INVERT_RESET = 8'hff;
localparam WCM_TCAM_KEY_INVERT_LO = 64;
localparam WCM_TCAM_KEY_INVERT_HI = 95;
localparam WCM_TCAM_KEY_INVERT_RESET = 32'hffffffff;
localparam WCM_TCAM_KEY_TOP_LO = 32;
localparam WCM_TCAM_KEY_TOP_HI = 39;
localparam WCM_TCAM_KEY_TOP_RESET = 8'hff;
localparam WCM_TCAM_KEY_LO = 0;
localparam WCM_TCAM_KEY_HI = 31;
localparam WCM_TCAM_KEY_RESET = 32'hffffffff;
localparam WCM_TCAM_USEMASK = 128'hFFFFFFFFFF000000FFFFFFFFFF;
localparam WCM_TCAM_RO_MASK = 128'h0;
localparam WCM_TCAM_WO_MASK = 128'h0;
localparam WCM_TCAM_RESET = 128'hFFFFFFFFFF000000FFFFFFFFFF;

typedef struct packed {
    logic [31:0] ACTION1;  // RW
    logic [31:0] ACTION0;  // RW
} WCM_ACTION_t;

localparam WCM_ACTION_REG_STRIDE = 48'h8;
localparam WCM_ACTION_REG_ENTRIES = 1024;
localparam WCM_ACTION_REGFILE_STRIDE = 48'h2000;
localparam WCM_ACTION_REGFILE_ENTRIES = 24;
localparam WCM_ACTION_CR_ADDR = 48'h100000;
localparam WCM_ACTION_SIZE = 64;
localparam WCM_ACTION_ACTION1_LO = 32;
localparam WCM_ACTION_ACTION1_HI = 63;
localparam WCM_ACTION_ACTION1_RESET = 32'h0;
localparam WCM_ACTION_ACTION0_LO = 0;
localparam WCM_ACTION_ACTION0_HI = 31;
localparam WCM_ACTION_ACTION0_RESET = 32'h0;
localparam WCM_ACTION_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam WCM_ACTION_RO_MASK = 64'h0;
localparam WCM_ACTION_WO_MASK = 64'h0;
localparam WCM_ACTION_RESET = 64'h0;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [15:0] CHUNK_MASK;  // RW
    logic  [0:0] START_COMPARE;  // RW
    logic  [0:0] START_SET;  // RW
    logic  [5:0] SELECT_TOP;  // RW
    logic  [6:0] SELECT0;  // RW
    logic  [6:0] SELECT1;  // RW
    logic  [6:0] SELECT2;  // RW
    logic  [6:0] SELECT3;  // RW
} WCM_TCAM_CFG_t;

localparam WCM_TCAM_CFG_REG_STRIDE = 48'h8;
localparam WCM_TCAM_CFG_REG_ENTRIES = 64;
localparam WCM_TCAM_CFG_REGFILE_STRIDE = 48'h200;
localparam WCM_TCAM_CFG_REGFILE_ENTRIES = 20;
localparam WCM_TCAM_CFG_CR_ADDR = 48'h130000;
localparam WCM_TCAM_CFG_SIZE = 64;
localparam WCM_TCAM_CFG_CHUNK_MASK_LO = 36;
localparam WCM_TCAM_CFG_CHUNK_MASK_HI = 51;
localparam WCM_TCAM_CFG_CHUNK_MASK_RESET = 16'hffff;
localparam WCM_TCAM_CFG_START_COMPARE_LO = 35;
localparam WCM_TCAM_CFG_START_COMPARE_HI = 35;
localparam WCM_TCAM_CFG_START_COMPARE_RESET = 1'h1;
localparam WCM_TCAM_CFG_START_SET_LO = 34;
localparam WCM_TCAM_CFG_START_SET_HI = 34;
localparam WCM_TCAM_CFG_START_SET_RESET = 1'h1;
localparam WCM_TCAM_CFG_SELECT_TOP_LO = 28;
localparam WCM_TCAM_CFG_SELECT_TOP_HI = 33;
localparam WCM_TCAM_CFG_SELECT_TOP_RESET = 6'h0;
localparam WCM_TCAM_CFG_SELECT0_LO = 21;
localparam WCM_TCAM_CFG_SELECT0_HI = 27;
localparam WCM_TCAM_CFG_SELECT0_RESET = 7'h0;
localparam WCM_TCAM_CFG_SELECT1_LO = 14;
localparam WCM_TCAM_CFG_SELECT1_HI = 20;
localparam WCM_TCAM_CFG_SELECT1_RESET = 7'h0;
localparam WCM_TCAM_CFG_SELECT2_LO = 7;
localparam WCM_TCAM_CFG_SELECT2_HI = 13;
localparam WCM_TCAM_CFG_SELECT2_RESET = 7'h0;
localparam WCM_TCAM_CFG_SELECT3_LO = 0;
localparam WCM_TCAM_CFG_SELECT3_HI = 6;
localparam WCM_TCAM_CFG_SELECT3_RESET = 7'h0;
localparam WCM_TCAM_CFG_USEMASK = 64'hFFFFFFFFFFFFF;
localparam WCM_TCAM_CFG_RO_MASK = 64'h0;
localparam WCM_TCAM_CFG_WO_MASK = 64'h0;
localparam WCM_TCAM_CFG_RESET = 64'hFFFFC00000000;

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic [23:0] ENABLE;  // RW
} WCM_ACTION_CFG_EN_t;

localparam WCM_ACTION_CFG_EN_REG_STRIDE = 48'h8;
localparam WCM_ACTION_CFG_EN_REG_ENTRIES = 64;
localparam WCM_ACTION_CFG_EN_CR_ADDR = 48'h132800;
localparam WCM_ACTION_CFG_EN_SIZE = 64;
localparam WCM_ACTION_CFG_EN_ENABLE_LO = 0;
localparam WCM_ACTION_CFG_EN_ENABLE_HI = 23;
localparam WCM_ACTION_CFG_EN_ENABLE_RESET = 1'h0;
localparam WCM_ACTION_CFG_EN_USEMASK = 64'hFFFFFF;
localparam WCM_ACTION_CFG_EN_RO_MASK = 64'h0;
localparam WCM_ACTION_CFG_EN_WO_MASK = 64'h0;
localparam WCM_ACTION_CFG_EN_RESET = 64'h0;

typedef struct packed {
    logic  [3:0] reserved0;  // RSVD
    logic [59:0] INDEX;  // RW
} IDX_t;

localparam IDX_REG_STRIDE = 48'h8;
localparam IDX_REG_ENTRIES = 2;
localparam WCM_ACTION_CFG_REGFILE_STRIDE = 48'h10;
localparam WCM_ACTION_CFG_REGFILE_ENTRIES = 64;
localparam IDX_CR_ADDR = 48'h132C00;
localparam IDX_SIZE = 64;
localparam IDX_INDEX_LO = 0;
localparam IDX_INDEX_HI = 59;
localparam IDX_INDEX_RESET = 'h0;
localparam IDX_USEMASK = 64'hFFFFFFFFFFFFFFF;
localparam IDX_RO_MASK = 64'h0;
localparam IDX_WO_MASK = 64'h0;
localparam IDX_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic  [3:0] HASH_ENTRY_RAM_C_ERR;  // RW/1C/V
    logic  [3:0] HASH_ENTRY_RAM_U_ERR;  // RW/1C/V
    logic  [2:0] FGHASH_ERR;  // RW/1C/V
    logic  [2:0] FGRP_ERR;  // RW/1C/V
    logic  [0:0] TCAM_SWEEP_ERR;  // RW/1C/V
    logic  [0:0] FCMN_SHELL_CTRL_ERR;  // RW/1C/V
} WCM_IP_t;

localparam WCM_IP_REG_STRIDE = 48'h8;
localparam WCM_IP_REG_ENTRIES = 1;
localparam [47:0] WCM_IP_CR_ADDR = 48'h133000;
localparam WCM_IP_SIZE = 64;
localparam WCM_IP_HASH_ENTRY_RAM_C_ERR_LO = 12;
localparam WCM_IP_HASH_ENTRY_RAM_C_ERR_HI = 15;
localparam WCM_IP_HASH_ENTRY_RAM_C_ERR_RESET = 4'h0;
localparam WCM_IP_HASH_ENTRY_RAM_U_ERR_LO = 8;
localparam WCM_IP_HASH_ENTRY_RAM_U_ERR_HI = 11;
localparam WCM_IP_HASH_ENTRY_RAM_U_ERR_RESET = 4'h0;
localparam WCM_IP_FGHASH_ERR_LO = 5;
localparam WCM_IP_FGHASH_ERR_HI = 7;
localparam WCM_IP_FGHASH_ERR_RESET = 3'h0;
localparam WCM_IP_FGRP_ERR_LO = 2;
localparam WCM_IP_FGRP_ERR_HI = 4;
localparam WCM_IP_FGRP_ERR_RESET = 3'h0;
localparam WCM_IP_TCAM_SWEEP_ERR_LO = 1;
localparam WCM_IP_TCAM_SWEEP_ERR_HI = 1;
localparam WCM_IP_TCAM_SWEEP_ERR_RESET = 1'h0;
localparam WCM_IP_FCMN_SHELL_CTRL_ERR_LO = 0;
localparam WCM_IP_FCMN_SHELL_CTRL_ERR_HI = 0;
localparam WCM_IP_FCMN_SHELL_CTRL_ERR_RESET = 1'h0;
localparam WCM_IP_USEMASK = 64'hFFFF;
localparam WCM_IP_RO_MASK = 64'h0;
localparam WCM_IP_WO_MASK = 64'h0;
localparam WCM_IP_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic  [3:0] HASH_ENTRY_RAM_C_ERR;  // RW
    logic  [3:0] HASH_ENTRY_RAM_U_ERR;  // RW
    logic  [2:0] FGHASH_ERR;  // RW
    logic  [2:0] FGRP_ERR;  // RW
    logic  [0:0] TCAM_SWEEP_ERR;  // RW
    logic  [0:0] FCMN_SHELL_CTRL_ERR;  // RW
} WCM_IM_t;

localparam WCM_IM_REG_STRIDE = 48'h8;
localparam WCM_IM_REG_ENTRIES = 1;
localparam [47:0] WCM_IM_CR_ADDR = 48'h133008;
localparam WCM_IM_SIZE = 64;
localparam WCM_IM_HASH_ENTRY_RAM_C_ERR_LO = 12;
localparam WCM_IM_HASH_ENTRY_RAM_C_ERR_HI = 15;
localparam WCM_IM_HASH_ENTRY_RAM_C_ERR_RESET = 4'h0;
localparam WCM_IM_HASH_ENTRY_RAM_U_ERR_LO = 8;
localparam WCM_IM_HASH_ENTRY_RAM_U_ERR_HI = 11;
localparam WCM_IM_HASH_ENTRY_RAM_U_ERR_RESET = 4'h0;
localparam WCM_IM_FGHASH_ERR_LO = 5;
localparam WCM_IM_FGHASH_ERR_HI = 7;
localparam WCM_IM_FGHASH_ERR_RESET = 3'h0;
localparam WCM_IM_FGRP_ERR_LO = 2;
localparam WCM_IM_FGRP_ERR_HI = 4;
localparam WCM_IM_FGRP_ERR_RESET = 3'h0;
localparam WCM_IM_TCAM_SWEEP_ERR_LO = 1;
localparam WCM_IM_TCAM_SWEEP_ERR_HI = 1;
localparam WCM_IM_TCAM_SWEEP_ERR_RESET = 1'h0;
localparam WCM_IM_FCMN_SHELL_CTRL_ERR_LO = 0;
localparam WCM_IM_FCMN_SHELL_CTRL_ERR_HI = 0;
localparam WCM_IM_FCMN_SHELL_CTRL_ERR_RESET = 1'h0;
localparam WCM_IM_USEMASK = 64'hFFFF;
localparam WCM_IM_RO_MASK = 64'h0;
localparam WCM_IM_WO_MASK = 64'h0;
localparam WCM_IM_RESET = 64'h0;

typedef struct packed {
    WCM_IP_t  WCM_IP;
    WCM_IM_t  WCM_IM;
} mby_ppe_cgrp_b_nested_map_registers_t;

// ===================================================
// load

typedef struct packed {
    logic  [0:0] HASH_ENTRY_RAM_C_ERR;  // RW/1C/V
    logic  [0:0] HASH_ENTRY_RAM_U_ERR;  // RW/1C/V
    logic  [0:0] FGHASH_ERR;  // RW/1C/V
    logic  [0:0] FGRP_ERR;  // RW/1C/V
    logic  [0:0] TCAM_SWEEP_ERR;  // RW/1C/V
    logic  [0:0] FCMN_SHELL_CTRL_ERR;  // RW/1C/V
} load_WCM_IP_t;

typedef struct packed {
    load_WCM_IP_t  WCM_IP;
} mby_ppe_cgrp_b_nested_map_load_t;

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

typedef struct packed {
    logic  [3:0] HASH_ENTRY_RAM_C_ERR;  // RW/1C/V
    logic  [3:0] HASH_ENTRY_RAM_U_ERR;  // RW/1C/V
    logic  [2:0] FGHASH_ERR;  // RW/1C/V
    logic  [2:0] FGRP_ERR;  // RW/1C/V
    logic  [0:0] TCAM_SWEEP_ERR;  // RW/1C/V
    logic  [0:0] FCMN_SHELL_CTRL_ERR;  // RW/1C/V
} new_WCM_IP_t;

typedef struct packed {
    new_WCM_IP_t  WCM_IP;
} mby_ppe_cgrp_b_nested_map_new_t;

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [15:0] we_EM_HASH_LOOKUP_t;

typedef logic [15:0] we_WCM_TCAM_t;

typedef logic [7:0] we_WCM_ACTION_t;

typedef logic [7:0] we_WCM_TCAM_CFG_t;

typedef logic [7:0] we_WCM_ACTION_CFG_EN_t;

typedef logic [7:0] we_IDX_t;

typedef struct packed {
    we_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    we_WCM_TCAM_t WCM_TCAM;
    we_WCM_ACTION_t WCM_ACTION;
    we_WCM_TCAM_CFG_t WCM_TCAM_CFG;
    we_WCM_ACTION_CFG_EN_t WCM_ACTION_CFG_EN;
    we_IDX_t IDX;
} mby_ppe_cgrp_b_nested_map_handcoded_t;

typedef logic [15:0] re_EM_HASH_LOOKUP_t;

typedef logic [15:0] re_WCM_TCAM_t;

typedef logic [7:0] re_WCM_ACTION_t;

typedef logic [7:0] re_WCM_TCAM_CFG_t;

typedef logic [7:0] re_WCM_ACTION_CFG_EN_t;

typedef logic [7:0] re_IDX_t;

typedef struct packed {
    re_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    re_WCM_TCAM_t WCM_TCAM;
    re_WCM_ACTION_t WCM_ACTION;
    re_WCM_TCAM_CFG_t WCM_TCAM_CFG;
    re_WCM_ACTION_CFG_EN_t WCM_ACTION_CFG_EN;
    re_IDX_t IDX;
} mby_ppe_cgrp_b_nested_map_hc_re_t;

typedef logic handcode_rvalid_EM_HASH_LOOKUP_t;

typedef logic handcode_rvalid_WCM_TCAM_t;

typedef logic handcode_rvalid_WCM_ACTION_t;

typedef logic handcode_rvalid_WCM_TCAM_CFG_t;

typedef logic handcode_rvalid_WCM_ACTION_CFG_EN_t;

typedef logic handcode_rvalid_IDX_t;

typedef struct packed {
    handcode_rvalid_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    handcode_rvalid_WCM_TCAM_t WCM_TCAM;
    handcode_rvalid_WCM_ACTION_t WCM_ACTION;
    handcode_rvalid_WCM_TCAM_CFG_t WCM_TCAM_CFG;
    handcode_rvalid_WCM_ACTION_CFG_EN_t WCM_ACTION_CFG_EN;
    handcode_rvalid_IDX_t IDX;
} mby_ppe_cgrp_b_nested_map_hc_rvalid_t;

typedef logic handcode_wvalid_EM_HASH_LOOKUP_t;

typedef logic handcode_wvalid_WCM_TCAM_t;

typedef logic handcode_wvalid_WCM_ACTION_t;

typedef logic handcode_wvalid_WCM_TCAM_CFG_t;

typedef logic handcode_wvalid_WCM_ACTION_CFG_EN_t;

typedef logic handcode_wvalid_IDX_t;

typedef struct packed {
    handcode_wvalid_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    handcode_wvalid_WCM_TCAM_t WCM_TCAM;
    handcode_wvalid_WCM_ACTION_t WCM_ACTION;
    handcode_wvalid_WCM_TCAM_CFG_t WCM_TCAM_CFG;
    handcode_wvalid_WCM_ACTION_CFG_EN_t WCM_ACTION_CFG_EN;
    handcode_wvalid_IDX_t IDX;
} mby_ppe_cgrp_b_nested_map_hc_wvalid_t;

typedef logic handcode_error_EM_HASH_LOOKUP_t;

typedef logic handcode_error_WCM_TCAM_t;

typedef logic handcode_error_WCM_ACTION_t;

typedef logic handcode_error_WCM_TCAM_CFG_t;

typedef logic handcode_error_WCM_ACTION_CFG_EN_t;

typedef logic handcode_error_IDX_t;

typedef struct packed {
    handcode_error_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    handcode_error_WCM_TCAM_t WCM_TCAM;
    handcode_error_WCM_ACTION_t WCM_ACTION;
    handcode_error_WCM_TCAM_CFG_t WCM_TCAM_CFG;
    handcode_error_WCM_ACTION_CFG_EN_t WCM_ACTION_CFG_EN;
    handcode_error_IDX_t IDX;
} mby_ppe_cgrp_b_nested_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    WCM_TCAM_t WCM_TCAM;
    WCM_ACTION_t WCM_ACTION;
    WCM_TCAM_CFG_t WCM_TCAM_CFG;
    WCM_ACTION_CFG_EN_t WCM_ACTION_CFG_EN;
    IDX_t IDX;
} mby_ppe_cgrp_b_nested_map_hc_reg_read_t;

typedef struct packed {
    EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    WCM_TCAM_t WCM_TCAM;
    WCM_ACTION_t WCM_ACTION;
    WCM_TCAM_CFG_t WCM_TCAM_CFG;
    WCM_ACTION_CFG_EN_t WCM_ACTION_CFG_EN;
    IDX_t IDX;
} mby_ppe_cgrp_b_nested_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_cgrp_b_nested_map_pkg

`endif // MBY_PPE_CGRP_B_NESTED_MAP_PKG_VH
