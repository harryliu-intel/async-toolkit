// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

module write_ecc
  (
input  logic [34-1:0] i_data,

output logic [34-1:0] o_data
,output logic [7-1:0] o_chk
  );
logic  xor0000;
logic  xor0001;
logic  xor0002;
logic  xor0003;
logic  xor0004;
logic  xor0005;
logic  xor0006;
logic  xor0007;
logic  xor0008;
logic  xor0009;
logic  xor0010;
logic  xor0011;
logic  xor0012;
logic  xor0013;
logic  xor0014;
logic  xor0015;
logic  xor0016;
logic  xor0017;
logic  xor0018;
logic  xor0019;
logic  xor0020;
logic  xor0021;
logic  xor0022;
logic  xor0023;
logic  xor0024;
logic  xor0025;
logic  xor0026;
logic  xor0027;
logic  xor0028;
logic  xor0029;
logic  xor0030;
logic  xor0031;
logic  xor0032;
logic  xor0033;
logic  xor0034;
logic  xor0035;
logic  xor0036;
logic  xor0037;
logic  xor0038;
logic  xor0039;
logic  xor0040;
logic  xor0041;
logic  xor0042;
logic  xor0043;
logic  xor0044;
logic  xor0045;
logic  xor0046;
logic  xor0047;
logic  xor0048;
logic  xor0049;
logic  xor0050;
logic[5:-1] ecc_parity;
logic[40:0] input_data;
assign xor0000 = (input_data[0001]^input_data[0000]^input_data[0003]^input_data[0002]); 
assign xor0001 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); 
assign xor0002 = (input_data[0009]^input_data[0008]^input_data[0011]^input_data[0010]); 
assign xor0003 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); 
assign xor0004 = (input_data[0019]^input_data[0018]^input_data[0017]^input_data[0016]); 
assign xor0005 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); 
assign xor0006 = (input_data[0025]^input_data[0024]^input_data[0027]^input_data[0026]); 
assign xor0007 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); 
assign xor0008 = (input_data[0035]^input_data[0034]^input_data[0033]^input_data[0032]); 
assign xor0009 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); 
assign xor0010 = input_data[0040];
assign xor0011 = (input_data[0005]^input_data[0007]^input_data[0001]^input_data[0003]); 
assign xor0012 = (input_data[0009]^input_data[0015]^input_data[0011]^input_data[0013]); 
assign xor0013 = (input_data[0019]^input_data[0017]^input_data[0021]^input_data[0023]); 
assign xor0014 = (input_data[0025]^input_data[0027]^input_data[0031]^input_data[0029]); 
assign xor0015 = (input_data[0035]^input_data[0037]^input_data[0033]^input_data[0039]); 
assign xor0016 = (input_data[0007]^input_data[0006]^input_data[0003]^input_data[0002]); 
assign xor0017 = (input_data[0015]^input_data[0014]^input_data[0011]^input_data[0010]); 
assign xor0018 = (input_data[0019]^input_data[0018]^input_data[0023]^input_data[0022]); 
assign xor0019 = (input_data[0027]^input_data[0031]^input_data[0030]^input_data[0026]); 
assign xor0020 = (input_data[0035]^input_data[0034]^input_data[0039]^input_data[0038]); 
assign xor0021 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); 
assign xor0022 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); 
assign xor0023 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); 
assign xor0024 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); 
assign xor0025 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); 
assign xor0026 = (xor0013^xor0014^xor0011^xor0012); 
assign xor0027 = xor0015;
assign xor0028 = (xor0027^xor0026); 
assign xor0029 = (xor0017^xor0018^xor0016^xor0019); 
assign xor0030 = xor0020;
assign xor0031 = (xor0030^xor0029); 
assign xor0032 = (xor0023^xor0024^xor0021^xor0022); 
assign xor0033 = xor0025;
assign xor0034 = (xor0033^xor0032); 
assign xor0035 = (xor0002^xor0010^xor0006^xor0022); 
assign xor0036 = xor0024;
assign xor0037 = (xor0035^xor0036); 
assign xor0038 = (xor0036^xor0023^xor0006^xor0004); 
assign xor0039 = (xor0010^xor0008^xor0033); 
assign xor0040 = (xor0002^xor0000^xor0021^xor0022); 
assign xor0041 = xor0038;
assign xor0042 = (xor0040^xor0041); 
assign xor0043 = (input_data[0009]^input_data[0005]^input_data[0006]^input_data[0003]); 
assign xor0044 = (input_data[0015]^input_data[0017]^input_data[0010]^input_data[0012]); 
assign xor0045 = (input_data[0018]^input_data[0024]^input_data[0020]^input_data[0023]); 
assign xor0046 = (input_data[0027]^input_data[0030]^input_data[0033]^input_data[0029]); 
assign xor0047 = (input_data[0034]^input_data[0036]^input_data[0039]); 
assign xor0048 = (xor0045^xor0010^xor0043^xor0044); 
assign xor0049 = (xor0046^xor0047); 
assign xor0050 = (xor0048^xor0049); 
assign ecc_parity[-1] = xor0050;
assign ecc_parity[0] = xor0028;
assign ecc_parity[1] = xor0031;
assign ecc_parity[2] = xor0034;
assign ecc_parity[3] = xor0037;
assign ecc_parity[4] = xor0038;
assign ecc_parity[5] = xor0039;
assign input_data[0] = '0;
assign o_chk     [0] = ecc_parity[0-1];
assign input_data[1] = '0;
assign o_chk     [1] = ecc_parity[1-1];
assign input_data[2] = '0;
assign o_chk     [2] = ecc_parity[2-1];
assign input_data[3] = i_data   [0];
assign o_data    [0] = i_data   [0];
assign input_data[4] = '0;
assign o_chk     [3] = ecc_parity[3-1];
assign input_data[5] = i_data   [1];
assign o_data    [1] = i_data   [1];
assign input_data[6] = i_data   [2];
assign o_data    [2] = i_data   [2];
assign input_data[7] = i_data   [3];
assign o_data    [3] = i_data   [3];
assign input_data[8] = '0;
assign o_chk     [4] = ecc_parity[4-1];
assign input_data[9] = i_data   [4];
assign o_data    [4] = i_data   [4];
assign input_data[10] = i_data   [5];
assign o_data    [5] = i_data   [5];
assign input_data[11] = i_data   [6];
assign o_data    [6] = i_data   [6];
assign input_data[12] = i_data   [7];
assign o_data    [7] = i_data   [7];
assign input_data[13] = i_data   [8];
assign o_data    [8] = i_data   [8];
assign input_data[14] = i_data   [9];
assign o_data    [9] = i_data   [9];
assign input_data[15] = i_data   [10];
assign o_data    [10] = i_data   [10];
assign input_data[16] = '0;
assign o_chk     [5] = ecc_parity[5-1];
assign input_data[17] = i_data   [11];
assign o_data    [11] = i_data   [11];
assign input_data[18] = i_data   [12];
assign o_data    [12] = i_data   [12];
assign input_data[19] = i_data   [13];
assign o_data    [13] = i_data   [13];
assign input_data[20] = i_data   [14];
assign o_data    [14] = i_data   [14];
assign input_data[21] = i_data   [15];
assign o_data    [15] = i_data   [15];
assign input_data[22] = i_data   [16];
assign o_data    [16] = i_data   [16];
assign input_data[23] = i_data   [17];
assign o_data    [17] = i_data   [17];
assign input_data[24] = i_data   [18];
assign o_data    [18] = i_data   [18];
assign input_data[25] = i_data   [19];
assign o_data    [19] = i_data   [19];
assign input_data[26] = i_data   [20];
assign o_data    [20] = i_data   [20];
assign input_data[27] = i_data   [21];
assign o_data    [21] = i_data   [21];
assign input_data[28] = i_data   [22];
assign o_data    [22] = i_data   [22];
assign input_data[29] = i_data   [23];
assign o_data    [23] = i_data   [23];
assign input_data[30] = i_data   [24];
assign o_data    [24] = i_data   [24];
assign input_data[31] = i_data   [25];
assign o_data    [25] = i_data   [25];
assign input_data[32] = '0;
assign o_chk     [6] = ecc_parity[6-1];
assign input_data[33] = i_data   [26];
assign o_data    [26] = i_data   [26];
assign input_data[34] = i_data   [27];
assign o_data    [27] = i_data   [27];
assign input_data[35] = i_data   [28];
assign o_data    [28] = i_data   [28];
assign input_data[36] = i_data   [29];
assign o_data    [29] = i_data   [29];
assign input_data[37] = i_data   [30];
assign o_data    [30] = i_data   [30];
assign input_data[38] = i_data   [31];
assign o_data    [31] = i_data   [31];
assign input_data[39] = i_data   [32];
assign o_data    [32] = i_data   [32];
assign input_data[40] = i_data   [33];
assign o_data    [33] = i_data   [33];
endmodule
