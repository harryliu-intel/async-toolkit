///
///  INTEL CONFIDENTIAL
///
///  Copyright 2017 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
// ---------------------------------------------------------------------------------------------------------------------
// -- Author : Jim McCormick <jim.mccormick@intel.com>
// -- Project Name : ??? 
// -- Description  : This file drives DUT reset 
// ---------------------------------------------------------------------------------------------------------------------

`ifndef SYSTEM_DRIVER_SV
`define SYSTEM_DRIVER_SV

class system_driver;

    virtual gcm_dut_if dut_if;

    string name;

    function new(virtual gcm_dut_if dut_if, configuration cfg);

        this.dut_if = dut_if;

        name = "System Driver";

    endfunction

    // Reset system
    task reset();
        dut_if.reset_n = 1;
        repeat (50) @(posedge dut_if.cclk);
        dut_if.reset_n = 0;
        repeat (50) @(posedge dut_if.cclk);
    endtask

endclass

`endif // SYSTEM_DRIVER_SV
