// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

//----------------------------------------------------------------------------------
// Package: mby_mgp_bfm_pkg
//
// Shared testbench environment components, objects and other definintions.
//-----------------------------------------------------------------------------------
package mby_mgp_bfm_pkg;

   `include "uvm_macros.svh"
   import uvm_pkg::*;
   import shdv_base_pkg::*;
    
   `include "mby_mgp_defines.svh"
   `include "mby_mgp_bfm_cfg.sv"
   `include "mby_mgp_req_seq_item.sv"
   `include "mby_mgp_req_seqr.sv"
   `include "mby_mgp_mem_crdt_io.sv"
   `include "mby_mgp_flow_ctrl.sv"
   `include "mby_mgp_req_drv.sv"
   `include "mby_mgp_req_mon.sv"
   `include "mby_mgp_req_agent.sv"
   `include "mby_mgp_req_agent_cfg.sv"
   `include "mby_mgp_bfm.sv"

endpackage
