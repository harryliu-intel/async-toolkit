magic
tech scmos
timestamp 965420787
<< ndiffusion >>
rect 91 128 103 129
rect 130 128 138 129
rect 91 120 103 125
rect 130 120 138 125
rect 91 112 103 117
rect 130 116 138 117
rect 91 108 103 109
rect 91 100 93 108
rect 101 100 103 108
rect 91 99 103 100
rect 130 107 138 108
rect 130 99 138 104
rect 91 91 103 96
rect 91 83 103 88
rect 130 95 138 96
rect 130 86 138 87
rect 91 79 103 80
rect 91 71 93 79
rect 101 71 103 79
rect 130 78 138 83
rect 91 70 103 71
rect 130 74 138 75
rect 91 64 103 67
rect 93 60 103 64
rect 130 65 138 66
rect 130 57 138 62
rect 130 53 138 54
<< pdiffusion >>
rect 154 128 162 129
rect 184 128 202 129
rect 154 120 162 125
rect 184 120 202 125
rect 154 116 162 117
rect 154 107 162 108
rect 154 99 162 104
rect 184 116 202 117
rect 200 108 202 116
rect 184 107 202 108
rect 184 99 202 104
rect 154 95 162 96
rect 154 86 162 87
rect 184 95 202 96
rect 200 87 202 95
rect 184 86 202 87
rect 154 78 162 83
rect 154 74 162 75
rect 154 65 162 66
rect 184 82 202 83
rect 184 77 194 82
rect 154 57 162 62
rect 184 58 189 63
rect 197 58 202 63
rect 184 57 202 58
rect 154 53 162 54
rect 184 53 202 54
<< ntransistor >>
rect 91 125 103 128
rect 130 125 138 128
rect 91 117 103 120
rect 130 117 138 120
rect 91 109 103 112
rect 130 104 138 107
rect 91 96 103 99
rect 130 96 138 99
rect 91 88 103 91
rect 130 83 138 86
rect 91 80 103 83
rect 130 75 138 78
rect 91 67 103 70
rect 130 62 138 65
rect 130 54 138 57
<< ptransistor >>
rect 154 125 162 128
rect 184 125 202 128
rect 154 117 162 120
rect 184 117 202 120
rect 154 104 162 107
rect 184 104 202 107
rect 154 96 162 99
rect 184 96 202 99
rect 154 83 162 86
rect 154 75 162 78
rect 184 83 202 86
rect 154 62 162 65
rect 154 54 162 57
rect 184 54 202 57
<< polysilicon >>
rect 87 125 91 128
rect 103 125 107 128
rect 118 125 130 128
rect 138 125 154 128
rect 162 125 184 128
rect 202 125 206 128
rect 118 120 121 125
rect 87 117 91 120
rect 103 117 121 120
rect 126 117 130 120
rect 138 117 154 120
rect 162 117 174 120
rect 180 117 184 120
rect 202 117 204 120
rect 118 112 121 117
rect 87 109 91 112
rect 103 109 105 112
rect 126 104 130 107
rect 138 104 154 107
rect 162 104 166 107
rect 105 99 108 104
rect 171 99 174 117
rect 204 107 207 112
rect 180 104 184 107
rect 202 104 207 107
rect 87 96 91 99
rect 103 96 108 99
rect 125 96 130 99
rect 138 96 154 99
rect 162 96 184 99
rect 202 96 206 99
rect 125 91 128 96
rect 87 88 91 91
rect 103 88 128 91
rect 125 86 128 88
rect 166 91 174 96
rect 125 83 130 86
rect 138 83 154 86
rect 162 83 166 86
rect 87 80 91 83
rect 103 80 107 83
rect 126 75 130 78
rect 138 75 154 78
rect 162 75 166 78
rect 87 67 91 70
rect 103 67 105 70
rect 118 57 121 70
rect 171 65 174 83
rect 179 83 184 86
rect 202 83 206 86
rect 179 74 182 83
rect 126 62 130 65
rect 138 62 154 65
rect 162 62 174 65
rect 118 54 130 57
rect 138 54 154 57
rect 162 54 166 57
rect 180 54 184 57
rect 202 54 206 57
<< ndcontact >>
rect 91 129 103 137
rect 130 129 138 137
rect 93 100 101 108
rect 130 108 138 116
rect 130 87 138 95
rect 93 71 101 79
rect 85 56 93 64
rect 130 66 138 74
rect 130 45 138 53
<< pdcontact >>
rect 154 129 162 137
rect 184 129 202 137
rect 154 108 162 116
rect 184 108 200 116
rect 154 87 162 95
rect 184 87 200 95
rect 154 66 162 74
rect 194 74 202 82
rect 189 58 197 66
rect 154 45 162 53
rect 184 45 202 53
<< polycontact >>
rect 105 104 113 112
rect 118 104 126 112
rect 204 112 212 120
rect 166 83 174 91
rect 118 70 126 78
rect 105 62 113 70
rect 179 66 187 74
<< metal1 >>
rect 91 129 138 137
rect 154 129 202 137
rect 109 120 208 124
rect 109 116 113 120
rect 85 112 113 116
rect 85 64 89 112
rect 93 100 101 108
rect 105 104 113 112
rect 97 96 109 100
rect 93 71 101 79
rect 85 56 93 64
rect 97 53 101 71
rect 105 70 109 96
rect 118 70 126 112
rect 130 108 200 116
rect 204 112 212 120
rect 130 87 138 95
rect 142 74 150 108
rect 158 95 189 99
rect 154 87 162 95
rect 166 83 174 91
rect 184 87 200 95
rect 204 82 208 112
rect 194 78 208 82
rect 194 74 202 78
rect 105 66 113 70
rect 130 66 187 74
rect 105 62 134 66
rect 179 58 197 66
rect 97 45 138 53
rect 154 45 202 53
<< labels >>
rlabel metal1 134 112 134 112 1 x
rlabel metal1 158 112 158 112 1 x
rlabel metal1 158 133 158 133 5 Vdd!
rlabel metal1 134 133 134 133 5 GND!
rlabel metal1 158 91 158 91 1 Vdd!
rlabel metal1 134 49 134 49 1 GND!
rlabel metal1 158 49 158 49 1 Vdd!
rlabel metal1 158 70 158 70 1 x
rlabel metal1 134 70 134 70 1 x
rlabel polysilicon 90 126 90 126 1 _SReset!
rlabel polysilicon 90 81 90 81 1 _SReset!
rlabel metal1 97 104 97 104 1 x
rlabel metal1 134 91 134 91 1 GND!
rlabel metal1 192 91 192 91 1 Vdd!
rlabel metal1 192 112 192 112 5 x
rlabel polysilicon 203 55 203 55 1 _PReset!
rlabel metal1 193 62 193 62 1 x
rlabel metal1 193 49 193 49 1 Vdd!
rlabel metal1 193 133 193 133 5 Vdd!
rlabel metal1 170 87 170 87 1 b
rlabel metal1 122 108 122 108 1 a
rlabel metal1 122 74 122 74 1 a
rlabel metal1 97 75 97 75 1 GND!
rlabel metal1 97 133 97 133 5 GND!
rlabel space 84 44 137 138 7 ^n
rlabel space 155 44 213 138 3 ^p
<< end >>
