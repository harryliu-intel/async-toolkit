//                                                                             
// File:       toplevel_fuse_env.svh                                           
// Creator:    kmoses1                                                         
// Time:       Thursday Jan 16, 2014 [3:40:08 pm]                              
//                                                                             
// Path:       /tmp/kmoses1/nebulon_run/1248                                   
// Arguments:  /p/com/eda/denali/blueprint/3.7.4/Linux/blueprint -cspec -fuse  
//             -html -I /p/com/eda/intel/nebulon/2.07p1/include/               
//             fusegen-Nebulon.rdl                                             
//                                                                             
// Sources:    /nfs/iil/proj/mpg/kmoses1_wa/SOCFuseGen/MBY/fusegen-Nebulon.rdl:5b3e806ef7d09a39437507f3cfbd0ecb
//             /p/com/eda/intel/nebulon/2.07p1/generators/fuse.pm              
//             /p/com/eda/intel/nebulon/2.07p1/generators/generator_common.pm  
//             /p/com/eda/intel/nebulon/2.07p1/generators/html.pm              
//             /p/com/eda/intel/nebulon/2.07p1/include/fuse_udp.rdl:c11891ce81c95bc748bf1f2bdbde2f6f
//             /usr/intel/pkgs/perl/5.8.7/lib64/5.8.7/Digest/base.pm           
//             /usr/intel/pkgs/perl/5.8.7/lib64/site_perl/Devel/StackTrace.pm  
//                                                                             
// Blueprint:   3.7.4 (Tue Jun 23 00:17:01 PDT 2009)                           
// Machine:    ivnc0059                                                        
// OS:         Linux 2.6.16.60-0.58.1.3835.0.PTF.638363-smp                    
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2014 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY DENALI BLUEPRINT, DO NOT EDIT       
//                                                                             


//Fuse code compatible with Saola versions: v20131113 and newer 

`ifndef SLA_PATH_TO_STRING
`define SLA_PATH_TO_STRING(SIG_PATH) `"SIG_PATH`"
`endif

package sla_fusegen_pkg;
import ovm_pkg::*;
import sla_pkg::*;
`include "ovm_macros.svh"
`include "sla_macros.svh"

`include "mby_classes.svh"

class toplevel_fuse_env extends sla_fuse_env;
   `ovm_component_utils(toplevel_fuse_env)

 rand mby_fuse_fusegroup mby_fuse;

function new (string name="fuse_env", ovm_component parent = null);
   super.new(name, parent);
endfunction // new

function void build();
   super.build();
   mby_fuse = mby_fuse_fusegroup::type_id::create("mby_fuse", this);
   mby_fuse.set_env(this);
   mby_fuse.set_fuse_id(8'haa);
   mby_fuse.add_fuses();

   add_group(mby_fuse);
endfunction

function void connect();
   super.connect();
endfunction

 function void set_desired_val(string fuse_name, logic val[]);
    sla_fuse f = get_fuse(fuse_name);
    f.set_desired_val(val);
 endfunction


 function string sprint_sv_fuse_env();  
   return({"Generated SV FUSE Env ---> ", `__FILE__}); 
 endfunction 

endclass

endpackage
