magic
tech scmos
timestamp 988943070
<< nselect >>
rect -50 49 0 91
<< pselect >>
rect 0 49 58 92
<< ndiffusion >>
rect -46 75 -42 78
rect -16 63 -8 64
rect -46 59 -42 62
rect -16 59 -8 60
<< pdiffusion >>
rect 45 80 53 81
rect 22 76 26 80
rect 8 63 16 64
rect 8 59 16 60
rect 22 59 26 72
rect 45 72 53 77
rect 45 68 53 69
<< ntransistor >>
rect -46 62 -42 75
rect -16 60 -8 63
<< ptransistor >>
rect 45 77 53 80
rect 22 72 26 76
rect 8 60 16 63
rect 45 69 53 72
<< polysilicon >>
rect -50 62 -46 75
rect -42 74 -38 75
rect -42 66 -40 74
rect 41 77 45 80
rect 53 77 57 80
rect 18 72 22 76
rect 26 72 28 76
rect -42 62 -38 66
rect -2 63 2 72
rect -20 60 -16 63
rect -8 60 8 63
rect 16 60 20 63
rect 41 69 45 72
rect 53 69 57 72
<< ndcontact >>
rect -49 78 -41 86
rect -16 64 -8 72
rect -49 51 -41 59
rect -16 51 -8 59
<< pdcontact >>
rect 22 80 30 88
rect 45 81 53 89
rect 8 64 16 72
rect 8 51 16 59
rect 45 60 53 68
rect 22 51 30 59
<< polycontact >>
rect -40 66 -32 74
rect -4 72 4 80
rect 28 68 36 76
<< metal1 >>
rect -49 83 53 89
rect -49 78 -41 83
rect -40 70 -32 74
rect -4 72 4 83
rect 22 80 30 83
rect 45 81 53 83
rect 28 72 36 76
rect -16 70 -8 72
rect -40 68 -8 70
rect 8 68 36 72
rect -40 66 16 68
rect -16 64 16 66
rect 45 59 53 68
rect -49 51 -8 59
rect 8 51 53 59
<< labels >>
rlabel metal1 -49 83 53 89 1 x
rlabel space 53 49 59 92 3 ^p
rlabel polysilicon 41 69 45 72 1 a|pin|w|3|poly
rlabel polysilicon 53 69 57 72 1 a|pin|w|3|poly
rlabel polysilicon 41 77 45 80 1 b|pin|w|4|poly
rlabel polysilicon 53 77 57 80 1 b|pin|w|4|poly
rlabel metal1 8 51 53 59 1 Vdd!
rlabel metal1 45 51 53 68 1 Vdd!
rlabel metal1 -49 51 -8 59 1 GND!
rlabel metal1 -4 72 4 89 1 x
rlabel metal1 -49 78 -41 89 3 x
rlabel metal1 45 81 53 89 1 x
rlabel metal1 22 80 30 88 1 x
<< end >>
