magic
tech scmos
timestamp 982687203
<< nselect >>
rect -74 40 0 140
<< pselect >>
rect 0 40 78 140
<< ndiffusion >>
rect -67 128 -55 129
rect -28 128 -8 129
rect -67 120 -55 125
rect -28 120 -8 125
rect -67 112 -55 117
rect -28 116 -8 117
rect -67 108 -55 109
rect -67 100 -65 108
rect -57 100 -55 108
rect -67 99 -55 100
rect -28 107 -8 108
rect -28 99 -8 104
rect -67 91 -55 96
rect -67 83 -55 88
rect -28 95 -8 96
rect -28 86 -8 87
rect -67 79 -55 80
rect -67 71 -65 79
rect -57 71 -55 79
rect -28 78 -8 83
rect -67 70 -55 71
rect -28 74 -8 75
rect -67 64 -55 67
rect -65 60 -55 64
rect -28 65 -8 66
rect -28 57 -8 62
rect -28 53 -8 54
<< pdiffusion >>
rect 8 128 28 129
rect 50 128 68 129
rect 8 120 28 125
rect 50 120 68 125
rect 8 116 28 117
rect 8 107 28 108
rect 8 99 28 104
rect 50 116 68 117
rect 66 108 68 116
rect 50 107 68 108
rect 50 99 68 104
rect 8 95 28 96
rect 8 86 28 87
rect 50 95 68 96
rect 66 87 68 95
rect 50 86 68 87
rect 8 78 28 83
rect 8 74 28 75
rect 8 65 28 66
rect 50 82 68 83
rect 50 77 60 82
rect 8 57 28 62
rect 54 58 59 63
rect 67 58 72 63
rect 54 57 72 58
rect 8 53 28 54
rect 54 53 72 54
rect 69 45 72 53
<< ntransistor >>
rect -67 125 -55 128
rect -28 125 -8 128
rect -67 117 -55 120
rect -28 117 -8 120
rect -67 109 -55 112
rect -28 104 -8 107
rect -67 96 -55 99
rect -28 96 -8 99
rect -67 88 -55 91
rect -28 83 -8 86
rect -67 80 -55 83
rect -28 75 -8 78
rect -67 67 -55 70
rect -28 62 -8 65
rect -28 54 -8 57
<< ptransistor >>
rect 8 125 28 128
rect 50 125 68 128
rect 8 117 28 120
rect 50 117 68 120
rect 8 104 28 107
rect 50 104 68 107
rect 8 96 28 99
rect 50 96 68 99
rect 8 83 28 86
rect 8 75 28 78
rect 50 83 68 86
rect 8 62 28 65
rect 8 54 28 57
rect 54 54 72 57
<< polysilicon >>
rect -71 125 -67 128
rect -55 125 -51 128
rect -40 125 -28 128
rect -8 125 8 128
rect 28 125 50 128
rect 68 125 72 128
rect -40 120 -37 125
rect -71 117 -67 120
rect -55 117 -37 120
rect -32 117 -28 120
rect -8 117 8 120
rect 28 117 40 120
rect 46 117 50 120
rect 68 117 70 120
rect -40 112 -37 117
rect -71 109 -67 112
rect -55 109 -53 112
rect -32 104 -28 107
rect -8 104 8 107
rect 28 104 32 107
rect -53 99 -50 104
rect 37 99 40 117
rect 70 107 73 112
rect 46 104 50 107
rect 68 104 73 107
rect -71 96 -67 99
rect -55 96 -50 99
rect -33 96 -28 99
rect -8 96 8 99
rect 28 96 50 99
rect 68 96 72 99
rect -33 91 -30 96
rect -71 88 -67 91
rect -55 88 -30 91
rect -33 86 -30 88
rect 32 91 40 96
rect -33 83 -28 86
rect -8 83 8 86
rect 28 83 32 86
rect -71 80 -67 83
rect -55 80 -51 83
rect -32 75 -28 78
rect -8 75 8 78
rect 28 75 32 78
rect -71 67 -67 70
rect -55 67 -53 70
rect -40 57 -37 70
rect 37 65 40 83
rect 45 83 50 86
rect 68 83 72 86
rect 45 74 48 83
rect -32 62 -28 65
rect -8 62 8 65
rect 28 62 40 65
rect -40 54 -28 57
rect -8 54 8 57
rect 28 54 32 57
rect 50 54 54 57
rect 72 54 76 57
<< ndcontact >>
rect -67 129 -55 137
rect -28 129 -8 137
rect -65 100 -57 108
rect -28 108 -8 116
rect -28 87 -8 95
rect -65 71 -57 79
rect -73 56 -65 64
rect -28 66 -8 74
rect -28 45 -8 53
<< pdcontact >>
rect 8 129 28 137
rect 50 129 68 137
rect 8 108 28 116
rect 50 108 66 116
rect 8 87 28 95
rect 50 87 66 95
rect 8 66 28 74
rect 60 74 68 82
rect 59 58 67 66
rect 8 45 28 53
rect 54 45 69 53
<< polycontact >>
rect -53 104 -45 112
rect -40 104 -32 112
rect 70 112 78 120
rect 32 83 40 91
rect -40 70 -32 78
rect -53 62 -45 70
rect 45 66 53 74
<< metal1 >>
rect -67 135 -8 137
rect -67 129 -27 135
rect -9 129 -8 135
rect 8 135 68 137
rect 8 129 9 135
rect 27 129 68 135
rect -49 120 74 124
rect -49 116 -45 120
rect -73 112 -45 116
rect -73 64 -69 112
rect -65 100 -57 108
rect -53 104 -45 112
rect -61 96 -49 100
rect -65 71 -57 79
rect -73 56 -65 64
rect -61 53 -57 71
rect -53 70 -49 96
rect -40 70 -32 112
rect -28 108 66 116
rect 70 112 78 120
rect -28 90 -27 95
rect -9 90 -8 95
rect -28 87 -8 90
rect -4 74 4 108
rect 21 96 58 101
rect 8 90 9 95
rect 27 95 58 96
rect 27 90 28 95
rect 8 87 28 90
rect 32 83 40 91
rect 50 87 66 95
rect 70 82 74 112
rect 60 78 74 82
rect 60 74 68 78
rect -28 70 28 74
rect 45 70 53 74
rect -53 66 -45 70
rect -28 66 53 70
rect -53 62 -21 66
rect 49 62 67 66
rect 59 58 67 62
rect -61 48 -8 53
rect -61 45 -27 48
rect -9 45 -8 48
rect 8 48 69 53
rect 8 45 9 48
rect 27 45 69 48
<< m2contact >>
rect -27 129 -9 135
rect 9 129 27 135
rect -27 90 -9 96
rect 9 90 27 96
rect -27 42 -9 48
rect 9 42 27 48
<< m3contact >>
rect -27 129 -9 135
rect 9 129 27 135
rect -27 90 -9 96
rect 9 90 27 96
rect -27 42 -9 48
rect 9 42 27 48
<< metal3 >>
rect -27 40 -9 140
rect 9 40 27 140
<< labels >>
rlabel metal1 -61 104 -61 104 1 x
rlabel metal1 -40 70 -32 112 1 a
rlabel metal1 63 62 63 62 1 x
rlabel metal1 32 83 40 91 1 b
rlabel space -75 40 -28 140 7 ^n
rlabel space 28 40 79 140 3 ^p
rlabel metal3 -27 40 -9 140 1 GND!|pin|s|0
rlabel metal3 9 40 27 140 1 Vdd!|pin|s|1
rlabel metal1 -67 129 -8 137 1 GND!|pin|s|0
rlabel metal1 -61 45 -8 53 1 GND!|pin|s|0
rlabel metal1 -61 45 -57 79 1 GND!|pin|s|0
rlabel metal1 8 129 68 137 1 Vdd!|pin|s|1
rlabel metal1 50 87 66 95 1 Vdd!|pin|s|1
rlabel metal1 8 45 69 53 1 Vdd!|pin|s|1
rlabel metal1 -4 66 4 116 1 x|pin|s|2
rlabel metal1 -28 66 28 74 1 x|pin|s|2
rlabel metal1 -28 108 66 116 1 x|pin|s|2
rlabel polysilicon -71 80 -67 83 1 _SReset!|pin|w|3|poly
rlabel polysilicon -71 125 -67 128 1 _SReset!|pin|w|4|poly
rlabel polysilicon -55 125 -51 128 1 _SReset!|pin|w|4|poly
rlabel polysilicon 50 54 54 57 1 _PReset!|pin|w|5|poly
rlabel polysilicon 72 54 76 57 1 _PReset!|pin|w|5|poly
<< end >>
