magic
tech scmos
timestamp 969760391
<< ndiffusion >>
rect -65 -5 -57 -4
rect -87 -10 -79 -9
rect -87 -18 -79 -13
rect -65 -9 -57 -8
rect -65 -18 -57 -17
rect -87 -22 -79 -21
rect -65 -22 -57 -21
<< pdiffusion >>
rect -134 -5 -126 -4
rect -134 -9 -126 -8
rect -113 -15 -109 -12
rect -41 -5 -33 -4
rect -134 -18 -126 -17
rect -134 -22 -126 -21
rect -113 -22 -109 -19
rect -41 -9 -33 -8
rect -41 -18 -33 -17
rect -41 -22 -33 -21
<< ntransistor >>
rect -65 -8 -57 -5
rect -87 -13 -79 -10
rect -87 -21 -79 -18
rect -65 -21 -57 -18
<< ptransistor >>
rect -134 -8 -126 -5
rect -41 -8 -33 -5
rect -134 -21 -126 -18
rect -113 -19 -109 -15
rect -41 -21 -33 -18
<< polysilicon >>
rect -124 -2 -89 1
rect -124 -5 -121 -2
rect -139 -8 -134 -5
rect -126 -8 -121 -5
rect -139 -18 -136 -8
rect -92 -10 -89 -2
rect -69 -5 -67 -2
rect -70 -8 -65 -5
rect -57 -8 -41 -5
rect -33 -8 -29 -5
rect -92 -13 -87 -10
rect -79 -13 -75 -10
rect -139 -21 -134 -18
rect -126 -21 -122 -18
rect -117 -19 -113 -15
rect -109 -19 -105 -15
rect -70 -18 -67 -8
rect -97 -21 -87 -18
rect -79 -21 -75 -18
rect -70 -21 -65 -18
rect -57 -21 -41 -18
rect -33 -21 -29 -18
<< ndcontact >>
rect -87 -9 -79 -1
rect -65 -4 -57 4
rect -65 -17 -57 -9
rect -87 -30 -79 -22
rect -65 -30 -57 -22
<< pdcontact >>
rect -134 -4 -126 4
rect -134 -17 -126 -9
rect -117 -12 -109 -4
rect -41 -4 -33 4
rect -41 -17 -33 -9
rect -134 -30 -126 -22
rect -117 -30 -109 -22
rect -41 -30 -33 -22
<< polycontact >>
rect -77 -5 -69 3
rect -105 -21 -97 -13
<< metal1 >>
rect -134 -4 -126 4
rect -77 -1 -69 3
rect -87 -4 -69 -1
rect -65 -4 -57 4
rect -41 -4 -33 4
rect -117 -6 -69 -4
rect -117 -9 -79 -6
rect -134 -12 -109 -9
rect -134 -14 -113 -12
rect -65 -13 -33 -9
rect -134 -17 -126 -14
rect -105 -17 -33 -13
rect -105 -21 -97 -17
rect -134 -30 -109 -22
rect -87 -30 -57 -22
rect -41 -30 -33 -22
<< labels >>
rlabel polysilicon -88 -12 -88 -12 1 a
rlabel polysilicon -88 -20 -88 -20 1 x
rlabel metal1 -83 -5 -83 -5 1 _x
rlabel metal1 -83 -26 -83 -26 1 GND!
rlabel polysilicon -114 -18 -114 -18 1 x
rlabel metal1 -113 -8 -113 -8 1 _x
rlabel metal1 -113 -26 -113 -26 1 Vdd!
rlabel ndcontact -61 -13 -61 -13 1 x
rlabel ndcontact -61 -26 -61 -26 1 GND!
rlabel ndcontact -61 0 -61 0 5 GND!
rlabel polysilicon -66 -20 -66 -20 3 _x
rlabel polysilicon -66 -7 -66 -7 3 _x
rlabel polysilicon -32 -20 -32 -20 1 _x
rlabel polysilicon -32 -7 -32 -7 1 _x
rlabel pdcontact -37 0 -37 0 5 Vdd!
rlabel pdcontact -37 -13 -37 -13 1 x
rlabel pdcontact -37 -26 -37 -26 1 Vdd!
rlabel metal1 -130 -13 -130 -13 1 _x
rlabel metal1 -130 -26 -130 -26 1 Vdd!
rlabel metal1 -130 0 -130 0 5 Vdd!
rlabel polysilicon -135 -20 -135 -20 1 a
rlabel polysilicon -135 -7 -135 -7 1 a
rlabel space -140 -30 -134 4 7 ^p1
rlabel space -33 -30 -28 4 3 ^p2
rlabel space -57 -31 -27 5 3 ^n2
<< end >>
