// -----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Raghu P Gudla
// Created On   :  09/22/2018
// Description  :  This directed sequence demonstrates the way user can control AXI BFM to generate AXI master transactions.
//                 this class defines a sequence in which a AXI WRITE followed by a AXI READ sequence is generated by assigning 
//                 values to the transactions rather than randomization, and then transmitted using `uvm_send.
//
// ----------------------------------------------------------------------------------------------------

//class fc_axi_basic_txn_seq extends svt_axi_master_base_sequence;
class fc_axi_basic_txn_seq extends fc_axi_master_base_seq;

    // parameter that controls the number of transactions that will be generated 
    rand int unsigned sequence_length = 10;

    //constrain the sequence length to a reasonable value 
    constraint reasonable_sequence_length {
        sequence_length <= 100;
    }
    
    `uvm_object_utils(fc_axi_basic_txn_seq)

    // class constructor 
    function new(string name="fc_axi_basic_txn_seq");
        super.new(name);
    endfunction

    virtual task body();
        svt_axi_master_transaction write_tran, read_tran;
        svt_configuration get_cfg;
        bit status;
        `uvm_info("body", "started running fc_axi_basic_txn_seq..", UVM_LOW)

        super.body();

        status = uvm_config_db #(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
        `uvm_info("body", $sformatf("sequence_length is %0d as a result of %0s.", sequence_length, status ? "config DB" : "randomization"), UVM_LOW);

        // obtain a handle to the port configuration 
        p_sequencer.get_cfg(get_cfg);
        if (!$cast(cfg, get_cfg)) begin
            `uvm_fatal("body", "unable to $cast the configuration to a svt_axi_port_configuration class");
        end

        for(int i = 0; i < sequence_length; i++) begin
        //for(int i = 0; i < 1; i++) begin

            // set up the write transaction 
            `uvm_create(write_tran)
            write_tran.port_cfg     = cfg;
            write_tran.xact_type    = svt_axi_transaction::WRITE;
            write_tran.addr         = 32'h0000_0100 | ('h100 << i);
            write_tran.burst_type   = svt_axi_transaction::INCR;
            write_tran.burst_size   = svt_axi_transaction::BURST_SIZE_32BIT;
            write_tran.atomic_type  = svt_axi_transaction::NORMAL;
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
            write_tran.burst_length = 1;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
            write_tran.burst_length = 2;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
            write_tran.burst_length = 4;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_4
            write_tran.burst_length = 8;
`else
            write_tran.burst_length = 16;
`endif
            write_tran.data         = new[write_tran.burst_length];
            write_tran.wstrb        = new[write_tran.burst_length];
            write_tran.data_user    = new[write_tran.burst_length];
            foreach (write_tran.data[i]) begin
                write_tran.data[i] = i;
            end
            foreach(write_tran.wstrb[i]) begin
                write_tran.wstrb[i] = 4'hf;
            end
            write_tran.wvalid_delay = new[write_tran.burst_length];
            foreach (write_tran.wvalid_delay[i]) begin
                write_tran.wvalid_delay[i]=i;
            end

            // send the write transaction 
            `uvm_send(write_tran)

            // wait for the write transaction to complete 
            get_response(rsp);

            `uvm_info("body", "AXI WRITE transaction completed", UVM_LOW);

            // set up the read transaction 
            `uvm_create(read_tran)
            read_tran.port_cfg     = cfg;
            read_tran.xact_type    = svt_axi_transaction::READ;
            read_tran.addr         = 32'h0000_0100 | ('h100 << i);
            read_tran.burst_type   = svt_axi_transaction::INCR;
            read_tran.burst_size   = svt_axi_transaction::BURST_SIZE_32BIT;
            read_tran.atomic_type  = svt_axi_transaction::NORMAL;
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
            read_tran.burst_length = 1;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
            read_tran.burst_length = 2;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
            read_tran.burst_length = 4;
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_4
            read_tran.burst_length = 8;
`else
            read_tran.burst_length = 16;
`endif
            read_tran.rresp        = new[read_tran.burst_length];
            read_tran.data         = new[read_tran.burst_length];
            read_tran.rready_delay = new[read_tran.burst_length];
            read_tran.data_user    = new[read_tran.burst_length];
            foreach (read_tran.rready_delay[i]) begin
                read_tran.rready_delay[i]=i;
            end

            // send the read transaction 
            `uvm_send(read_tran)

            // wait for the read transaction to complete 
            get_response(rsp);

            `uvm_info("body", "AXI READ transaction completed", UVM_LOW);
        end

        `uvm_info("body", "exiting...", UVM_LOW)
    endtask: body

endclass: fc_axi_basic_txn_seq



