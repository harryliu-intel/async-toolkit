magic
tech scmos
timestamp 988943070
<< nselect >>
rect -46 99 0 125
rect -69 60 0 99
<< pselect >>
rect 0 99 46 125
rect 0 60 69 99
<< ndiffusion >>
rect -40 113 -8 114
rect -40 109 -8 110
rect -40 101 -28 109
rect -40 100 -8 101
rect -40 96 -8 97
rect -20 88 -8 96
rect -40 87 -8 88
rect -64 82 -60 86
rect -40 83 -8 84
rect -40 74 -8 75
rect -64 70 -60 74
rect -40 70 -8 71
<< pdiffusion >>
rect 8 113 40 114
rect 8 109 40 110
rect 28 101 40 109
rect 8 100 40 101
rect 8 96 40 97
rect 8 88 26 96
rect 8 87 40 88
rect 8 83 40 84
rect 8 74 40 75
rect 60 82 64 86
rect 8 70 40 71
rect 60 70 64 78
<< ntransistor >>
rect -40 110 -8 113
rect -40 97 -8 100
rect -40 84 -8 87
rect -64 74 -60 82
rect -40 71 -8 74
<< ptransistor >>
rect 8 110 40 113
rect 8 97 40 100
rect 8 84 40 87
rect 60 78 64 82
rect 8 71 40 74
<< polysilicon >>
rect -45 110 -40 113
rect -8 110 8 113
rect 40 110 45 113
rect -45 100 -42 110
rect -4 100 4 110
rect 42 100 45 110
rect -45 97 -40 100
rect -8 97 8 100
rect 40 97 45 100
rect -45 95 -42 97
rect -44 87 -42 95
rect -4 96 4 97
rect -45 84 -40 87
rect -8 84 -4 87
rect -68 74 -64 82
rect -60 74 -58 82
rect -45 74 -42 84
rect 42 95 45 97
rect 42 87 44 95
rect 4 84 8 87
rect 40 84 45 87
rect 42 74 45 84
rect 58 78 60 82
rect 64 78 68 82
rect -45 71 -40 74
rect -8 71 8 74
rect 40 71 45 74
<< ndcontact >>
rect -40 114 -8 122
rect -28 101 -8 109
rect -64 86 -56 94
rect -40 88 -20 96
rect -40 75 -8 83
rect -64 62 -56 70
rect -40 62 -8 70
<< pdcontact >>
rect 8 114 40 122
rect 8 101 28 109
rect 26 88 40 96
rect 56 86 64 94
rect 8 75 40 83
rect 8 62 40 70
rect 56 62 64 70
<< polycontact >>
rect -52 87 -44 95
rect -58 74 -50 82
rect -4 74 4 96
rect 44 87 52 95
rect 50 74 58 82
<< metal1 >>
rect -40 114 -8 122
rect 8 114 40 122
rect -40 96 -32 114
rect -28 101 28 109
rect -52 94 -44 95
rect -64 87 -44 94
rect -40 88 -20 96
rect -64 86 -56 87
rect -16 83 -8 101
rect -40 82 -8 83
rect -58 75 -8 82
rect -58 74 -50 75
rect -4 74 4 96
rect 8 83 16 101
rect 32 96 40 114
rect 26 88 40 96
rect 44 94 52 95
rect 44 87 64 94
rect 56 86 64 87
rect 8 82 40 83
rect 8 75 58 82
rect 50 74 58 75
rect -64 62 -8 70
rect 8 62 64 70
<< labels >>
rlabel metal1 -4 74 4 96 1 _x
rlabel metal1 -48 91 -48 91 1 _x
rlabel metal1 48 91 48 91 1 _x
rlabel space -69 60 -28 125 7 ^n
rlabel space 28 60 69 125 3 ^p
rlabel metal1 -40 88 -32 122 1 GND!|pin|s|0
rlabel metal1 -40 88 -20 96 1 GND!|pin|s|0
rlabel metal1 26 88 40 96 1 Vdd!|pin|s|1
rlabel metal1 32 88 40 122 1 Vdd!|pin|s|1
rlabel metal1 -58 75 -8 82 1 x|pin|s|2
rlabel metal1 -28 101 28 109 1 x|pin|s|2
rlabel metal1 8 75 58 82 1 x|pin|s|2
rlabel metal1 8 75 16 109 1 x|pin|s|2
rlabel metal1 -16 75 -8 109 1 x|pin|s|2
rlabel metal1 -40 114 -8 122 1 GND!|pin|s|0
rlabel metal1 8 114 40 122 1 Vdd!|pin|s|1
rlabel metal1 -64 62 -8 70 1 GND!|pin|s|1
rlabel metal1 8 62 64 70 1 Vdd!|pin|s|0
<< end >>
