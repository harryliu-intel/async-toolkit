///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Jon Bagge <jon.bagge.com> 
// -- Project Name : MBY 
// -- Description  : parser netlist. 
// ------------------------------------------------------------------- 

module parser_top (
input reset, 
ahb_rx_ppe_if.ppe ahb_rx_ppe_if, 
glb_rx_ppe_if.ppe glb_rx_ppe_if, 
igr_rx_ppe_if.ppe igr_rx_ppe_if, 
//Input List
input                   cclk                                      
);

logic [104:0] parser_parser_ana_cam_0_from_mem;
logic [119:0] parser_parser_ana_cam_0_to_mem; 
logic [104:0] parser_parser_ana_cam_10_from_mem;
logic [119:0] parser_parser_ana_cam_10_to_mem;
logic [104:0] parser_parser_ana_cam_11_from_mem;
logic [119:0] parser_parser_ana_cam_11_to_mem;
logic [104:0] parser_parser_ana_cam_12_from_mem;
logic [119:0] parser_parser_ana_cam_12_to_mem;
logic [104:0] parser_parser_ana_cam_13_from_mem;
logic [119:0] parser_parser_ana_cam_13_to_mem;
logic [104:0] parser_parser_ana_cam_14_from_mem;
logic [119:0] parser_parser_ana_cam_14_to_mem;
logic [104:0] parser_parser_ana_cam_15_from_mem;
logic [119:0] parser_parser_ana_cam_15_to_mem;
logic [104:0] parser_parser_ana_cam_16_from_mem;
logic [119:0] parser_parser_ana_cam_16_to_mem;
logic [104:0] parser_parser_ana_cam_17_from_mem;
logic [119:0] parser_parser_ana_cam_17_to_mem;
logic [104:0] parser_parser_ana_cam_18_from_mem;
logic [119:0] parser_parser_ana_cam_18_to_mem;
logic [104:0] parser_parser_ana_cam_19_from_mem;
logic [119:0] parser_parser_ana_cam_19_to_mem;
logic [104:0] parser_parser_ana_cam_1_from_mem;
logic [119:0] parser_parser_ana_cam_1_to_mem; 
logic [104:0] parser_parser_ana_cam_20_from_mem;
logic [119:0] parser_parser_ana_cam_20_to_mem;
logic [104:0] parser_parser_ana_cam_21_from_mem;
logic [119:0] parser_parser_ana_cam_21_to_mem;
logic [104:0] parser_parser_ana_cam_22_from_mem;
logic [119:0] parser_parser_ana_cam_22_to_mem;
logic [104:0] parser_parser_ana_cam_23_from_mem;
logic [119:0] parser_parser_ana_cam_23_to_mem;
logic [104:0] parser_parser_ana_cam_24_from_mem;
logic [119:0] parser_parser_ana_cam_24_to_mem;
logic [104:0] parser_parser_ana_cam_25_from_mem;
logic [119:0] parser_parser_ana_cam_25_to_mem;
logic [104:0] parser_parser_ana_cam_26_from_mem;
logic [119:0] parser_parser_ana_cam_26_to_mem;
logic [104:0] parser_parser_ana_cam_27_from_mem;
logic [119:0] parser_parser_ana_cam_27_to_mem;
logic [104:0] parser_parser_ana_cam_28_from_mem;
logic [119:0] parser_parser_ana_cam_28_to_mem;
logic [104:0] parser_parser_ana_cam_29_from_mem;
logic [119:0] parser_parser_ana_cam_29_to_mem;
logic [104:0] parser_parser_ana_cam_2_from_mem;
logic [119:0] parser_parser_ana_cam_2_to_mem; 
logic [104:0] parser_parser_ana_cam_30_from_mem;
logic [119:0] parser_parser_ana_cam_30_to_mem;
logic [104:0] parser_parser_ana_cam_31_from_mem;
logic [119:0] parser_parser_ana_cam_31_to_mem;
logic [104:0] parser_parser_ana_cam_3_from_mem;
logic [119:0] parser_parser_ana_cam_3_to_mem; 
logic [104:0] parser_parser_ana_cam_4_from_mem;
logic [119:0] parser_parser_ana_cam_4_to_mem; 
logic [104:0] parser_parser_ana_cam_5_from_mem;
logic [119:0] parser_parser_ana_cam_5_to_mem; 
logic [104:0] parser_parser_ana_cam_6_from_mem;
logic [119:0] parser_parser_ana_cam_6_to_mem; 
logic [104:0] parser_parser_ana_cam_7_from_mem;
logic [119:0] parser_parser_ana_cam_7_to_mem; 
logic [104:0] parser_parser_ana_cam_8_from_mem;
logic [119:0] parser_parser_ana_cam_8_to_mem; 
logic [104:0] parser_parser_ana_cam_9_from_mem;
logic [119:0] parser_parser_ana_cam_9_to_mem; 
logic  [14:0] parser_parser_ana_exc_0_from_mem;
logic  [29:0] parser_parser_ana_exc_0_to_mem; 
logic  [14:0] parser_parser_ana_exc_10_from_mem;
logic  [29:0] parser_parser_ana_exc_10_to_mem;
logic  [14:0] parser_parser_ana_exc_11_from_mem;
logic  [29:0] parser_parser_ana_exc_11_to_mem;
logic  [14:0] parser_parser_ana_exc_12_from_mem;
logic  [29:0] parser_parser_ana_exc_12_to_mem;
logic  [14:0] parser_parser_ana_exc_13_from_mem;
logic  [29:0] parser_parser_ana_exc_13_to_mem;
logic  [14:0] parser_parser_ana_exc_14_from_mem;
logic  [29:0] parser_parser_ana_exc_14_to_mem;
logic  [14:0] parser_parser_ana_exc_15_from_mem;
logic  [29:0] parser_parser_ana_exc_15_to_mem;
logic  [14:0] parser_parser_ana_exc_16_from_mem;
logic  [29:0] parser_parser_ana_exc_16_to_mem;
logic  [14:0] parser_parser_ana_exc_17_from_mem;
logic  [29:0] parser_parser_ana_exc_17_to_mem;
logic  [14:0] parser_parser_ana_exc_18_from_mem;
logic  [29:0] parser_parser_ana_exc_18_to_mem;
logic  [14:0] parser_parser_ana_exc_19_from_mem;
logic  [29:0] parser_parser_ana_exc_19_to_mem;
logic  [14:0] parser_parser_ana_exc_1_from_mem;
logic  [29:0] parser_parser_ana_exc_1_to_mem; 
logic  [14:0] parser_parser_ana_exc_20_from_mem;
logic  [29:0] parser_parser_ana_exc_20_to_mem;
logic  [14:0] parser_parser_ana_exc_21_from_mem;
logic  [29:0] parser_parser_ana_exc_21_to_mem;
logic  [14:0] parser_parser_ana_exc_22_from_mem;
logic  [29:0] parser_parser_ana_exc_22_to_mem;
logic  [14:0] parser_parser_ana_exc_23_from_mem;
logic  [29:0] parser_parser_ana_exc_23_to_mem;
logic  [14:0] parser_parser_ana_exc_24_from_mem;
logic  [29:0] parser_parser_ana_exc_24_to_mem;
logic  [14:0] parser_parser_ana_exc_25_from_mem;
logic  [29:0] parser_parser_ana_exc_25_to_mem;
logic  [14:0] parser_parser_ana_exc_26_from_mem;
logic  [29:0] parser_parser_ana_exc_26_to_mem;
logic  [14:0] parser_parser_ana_exc_27_from_mem;
logic  [29:0] parser_parser_ana_exc_27_to_mem;
logic  [14:0] parser_parser_ana_exc_28_from_mem;
logic  [29:0] parser_parser_ana_exc_28_to_mem;
logic  [14:0] parser_parser_ana_exc_29_from_mem;
logic  [29:0] parser_parser_ana_exc_29_to_mem;
logic  [14:0] parser_parser_ana_exc_2_from_mem;
logic  [29:0] parser_parser_ana_exc_2_to_mem; 
logic  [14:0] parser_parser_ana_exc_30_from_mem;
logic  [29:0] parser_parser_ana_exc_30_to_mem;
logic  [14:0] parser_parser_ana_exc_31_from_mem;
logic  [29:0] parser_parser_ana_exc_31_to_mem;
logic  [14:0] parser_parser_ana_exc_3_from_mem;
logic  [29:0] parser_parser_ana_exc_3_to_mem; 
logic  [14:0] parser_parser_ana_exc_4_from_mem;
logic  [29:0] parser_parser_ana_exc_4_to_mem; 
logic  [14:0] parser_parser_ana_exc_5_from_mem;
logic  [29:0] parser_parser_ana_exc_5_to_mem; 
logic  [14:0] parser_parser_ana_exc_6_from_mem;
logic  [29:0] parser_parser_ana_exc_6_to_mem; 
logic  [14:0] parser_parser_ana_exc_7_from_mem;
logic  [29:0] parser_parser_ana_exc_7_to_mem; 
logic  [14:0] parser_parser_ana_exc_8_from_mem;
logic  [29:0] parser_parser_ana_exc_8_to_mem; 
logic  [14:0] parser_parser_ana_exc_9_from_mem;
logic  [29:0] parser_parser_ana_exc_9_to_mem; 
logic  [32:0] parser_parser_ana_ext_0_from_mem;
logic  [49:0] parser_parser_ana_ext_0_to_mem; 
logic  [32:0] parser_parser_ana_ext_10_from_mem;
logic  [49:0] parser_parser_ana_ext_10_to_mem;
logic  [32:0] parser_parser_ana_ext_11_from_mem;
logic  [49:0] parser_parser_ana_ext_11_to_mem;
logic  [32:0] parser_parser_ana_ext_12_from_mem;
logic  [49:0] parser_parser_ana_ext_12_to_mem;
logic  [32:0] parser_parser_ana_ext_13_from_mem;
logic  [49:0] parser_parser_ana_ext_13_to_mem;
logic  [32:0] parser_parser_ana_ext_14_from_mem;
logic  [49:0] parser_parser_ana_ext_14_to_mem;
logic  [32:0] parser_parser_ana_ext_15_from_mem;
logic  [49:0] parser_parser_ana_ext_15_to_mem;
logic  [32:0] parser_parser_ana_ext_16_from_mem;
logic  [49:0] parser_parser_ana_ext_16_to_mem;
logic  [32:0] parser_parser_ana_ext_17_from_mem;
logic  [49:0] parser_parser_ana_ext_17_to_mem;
logic  [32:0] parser_parser_ana_ext_18_from_mem;
logic  [49:0] parser_parser_ana_ext_18_to_mem;
logic  [32:0] parser_parser_ana_ext_19_from_mem;
logic  [49:0] parser_parser_ana_ext_19_to_mem;
logic  [32:0] parser_parser_ana_ext_1_from_mem;
logic  [49:0] parser_parser_ana_ext_1_to_mem; 
logic  [32:0] parser_parser_ana_ext_20_from_mem;
logic  [49:0] parser_parser_ana_ext_20_to_mem;
logic  [32:0] parser_parser_ana_ext_21_from_mem;
logic  [49:0] parser_parser_ana_ext_21_to_mem;
logic  [32:0] parser_parser_ana_ext_22_from_mem;
logic  [49:0] parser_parser_ana_ext_22_to_mem;
logic  [32:0] parser_parser_ana_ext_23_from_mem;
logic  [49:0] parser_parser_ana_ext_23_to_mem;
logic  [32:0] parser_parser_ana_ext_24_from_mem;
logic  [49:0] parser_parser_ana_ext_24_to_mem;
logic  [32:0] parser_parser_ana_ext_25_from_mem;
logic  [49:0] parser_parser_ana_ext_25_to_mem;
logic  [32:0] parser_parser_ana_ext_26_from_mem;
logic  [49:0] parser_parser_ana_ext_26_to_mem;
logic  [32:0] parser_parser_ana_ext_27_from_mem;
logic  [49:0] parser_parser_ana_ext_27_to_mem;
logic  [32:0] parser_parser_ana_ext_28_from_mem;
logic  [49:0] parser_parser_ana_ext_28_to_mem;
logic  [32:0] parser_parser_ana_ext_29_from_mem;
logic  [49:0] parser_parser_ana_ext_29_to_mem;
logic  [32:0] parser_parser_ana_ext_2_from_mem;
logic  [49:0] parser_parser_ana_ext_2_to_mem; 
logic  [32:0] parser_parser_ana_ext_30_from_mem;
logic  [49:0] parser_parser_ana_ext_30_to_mem;
logic  [32:0] parser_parser_ana_ext_31_from_mem;
logic  [49:0] parser_parser_ana_ext_31_to_mem;
logic  [32:0] parser_parser_ana_ext_3_from_mem;
logic  [49:0] parser_parser_ana_ext_3_to_mem; 
logic  [32:0] parser_parser_ana_ext_4_from_mem;
logic  [49:0] parser_parser_ana_ext_4_to_mem; 
logic  [32:0] parser_parser_ana_ext_5_from_mem;
logic  [49:0] parser_parser_ana_ext_5_to_mem; 
logic  [32:0] parser_parser_ana_ext_6_from_mem;
logic  [49:0] parser_parser_ana_ext_6_to_mem; 
logic  [32:0] parser_parser_ana_ext_7_from_mem;
logic  [49:0] parser_parser_ana_ext_7_to_mem; 
logic  [32:0] parser_parser_ana_ext_8_from_mem;
logic  [49:0] parser_parser_ana_ext_8_to_mem; 
logic  [32:0] parser_parser_ana_ext_9_from_mem;
logic  [49:0] parser_parser_ana_ext_9_to_mem; 
logic  [55:0] parser_parser_ana_s_0_from_mem; 
logic  [70:0] parser_parser_ana_s_0_to_mem;   
logic  [55:0] parser_parser_ana_s_10_from_mem;
logic  [70:0] parser_parser_ana_s_10_to_mem;  
logic  [55:0] parser_parser_ana_s_11_from_mem;
logic  [70:0] parser_parser_ana_s_11_to_mem;  
logic  [55:0] parser_parser_ana_s_12_from_mem;
logic  [70:0] parser_parser_ana_s_12_to_mem;  
logic  [55:0] parser_parser_ana_s_13_from_mem;
logic  [70:0] parser_parser_ana_s_13_to_mem;  
logic  [55:0] parser_parser_ana_s_14_from_mem;
logic  [70:0] parser_parser_ana_s_14_to_mem;  
logic  [55:0] parser_parser_ana_s_15_from_mem;
logic  [70:0] parser_parser_ana_s_15_to_mem;  
logic  [55:0] parser_parser_ana_s_16_from_mem;
logic  [70:0] parser_parser_ana_s_16_to_mem;  
logic  [55:0] parser_parser_ana_s_17_from_mem;
logic  [70:0] parser_parser_ana_s_17_to_mem;  
logic  [55:0] parser_parser_ana_s_18_from_mem;
logic  [70:0] parser_parser_ana_s_18_to_mem;  
logic  [55:0] parser_parser_ana_s_19_from_mem;
logic  [70:0] parser_parser_ana_s_19_to_mem;  
logic  [55:0] parser_parser_ana_s_1_from_mem; 
logic  [70:0] parser_parser_ana_s_1_to_mem;   
logic  [55:0] parser_parser_ana_s_20_from_mem;
logic  [70:0] parser_parser_ana_s_20_to_mem;  
logic  [55:0] parser_parser_ana_s_21_from_mem;
logic  [70:0] parser_parser_ana_s_21_to_mem;  
logic  [55:0] parser_parser_ana_s_22_from_mem;
logic  [70:0] parser_parser_ana_s_22_to_mem;  
logic  [55:0] parser_parser_ana_s_23_from_mem;
logic  [70:0] parser_parser_ana_s_23_to_mem;  
logic  [55:0] parser_parser_ana_s_24_from_mem;
logic  [70:0] parser_parser_ana_s_24_to_mem;  
logic  [55:0] parser_parser_ana_s_25_from_mem;
logic  [70:0] parser_parser_ana_s_25_to_mem;  
logic  [55:0] parser_parser_ana_s_26_from_mem;
logic  [70:0] parser_parser_ana_s_26_to_mem;  
logic  [55:0] parser_parser_ana_s_27_from_mem;
logic  [70:0] parser_parser_ana_s_27_to_mem;  
logic  [55:0] parser_parser_ana_s_28_from_mem;
logic  [70:0] parser_parser_ana_s_28_to_mem;  
logic  [55:0] parser_parser_ana_s_29_from_mem;
logic  [70:0] parser_parser_ana_s_29_to_mem;  
logic  [55:0] parser_parser_ana_s_2_from_mem; 
logic  [70:0] parser_parser_ana_s_2_to_mem;   
logic  [55:0] parser_parser_ana_s_30_from_mem;
logic  [70:0] parser_parser_ana_s_30_to_mem;  
logic  [55:0] parser_parser_ana_s_31_from_mem;
logic  [70:0] parser_parser_ana_s_31_to_mem;  
logic  [55:0] parser_parser_ana_s_3_from_mem; 
logic  [70:0] parser_parser_ana_s_3_to_mem;   
logic  [55:0] parser_parser_ana_s_4_from_mem; 
logic  [70:0] parser_parser_ana_s_4_to_mem;   
logic  [55:0] parser_parser_ana_s_5_from_mem; 
logic  [70:0] parser_parser_ana_s_5_to_mem;   
logic  [55:0] parser_parser_ana_s_6_from_mem; 
logic  [70:0] parser_parser_ana_s_6_to_mem;   
logic  [55:0] parser_parser_ana_s_7_from_mem; 
logic  [70:0] parser_parser_ana_s_7_to_mem;   
logic  [55:0] parser_parser_ana_s_8_from_mem; 
logic  [70:0] parser_parser_ana_s_8_to_mem;   
logic  [55:0] parser_parser_ana_s_9_from_mem; 
logic  [70:0] parser_parser_ana_s_9_to_mem;   
logic  [39:0] parser_parser_ana_w_0_from_mem; 
logic  [54:0] parser_parser_ana_w_0_to_mem;   
logic  [39:0] parser_parser_ana_w_10_from_mem;
logic  [54:0] parser_parser_ana_w_10_to_mem;  
logic  [39:0] parser_parser_ana_w_11_from_mem;
logic  [54:0] parser_parser_ana_w_11_to_mem;  
logic  [39:0] parser_parser_ana_w_12_from_mem;
logic  [54:0] parser_parser_ana_w_12_to_mem;  
logic  [39:0] parser_parser_ana_w_13_from_mem;
logic  [54:0] parser_parser_ana_w_13_to_mem;  
logic  [39:0] parser_parser_ana_w_14_from_mem;
logic  [54:0] parser_parser_ana_w_14_to_mem;  
logic  [39:0] parser_parser_ana_w_15_from_mem;
logic  [54:0] parser_parser_ana_w_15_to_mem;  
logic  [39:0] parser_parser_ana_w_16_from_mem;
logic  [54:0] parser_parser_ana_w_16_to_mem;  
logic  [39:0] parser_parser_ana_w_17_from_mem;
logic  [54:0] parser_parser_ana_w_17_to_mem;  
logic  [39:0] parser_parser_ana_w_18_from_mem;
logic  [54:0] parser_parser_ana_w_18_to_mem;  
logic  [39:0] parser_parser_ana_w_19_from_mem;
logic  [54:0] parser_parser_ana_w_19_to_mem;  
logic  [39:0] parser_parser_ana_w_1_from_mem; 
logic  [54:0] parser_parser_ana_w_1_to_mem;   
logic  [39:0] parser_parser_ana_w_20_from_mem;
logic  [54:0] parser_parser_ana_w_20_to_mem;  
logic  [39:0] parser_parser_ana_w_21_from_mem;
logic  [54:0] parser_parser_ana_w_21_to_mem;  
logic  [39:0] parser_parser_ana_w_22_from_mem;
logic  [54:0] parser_parser_ana_w_22_to_mem;  
logic  [39:0] parser_parser_ana_w_23_from_mem;
logic  [54:0] parser_parser_ana_w_23_to_mem;  
logic  [39:0] parser_parser_ana_w_24_from_mem;
logic  [54:0] parser_parser_ana_w_24_to_mem;  
logic  [39:0] parser_parser_ana_w_25_from_mem;
logic  [54:0] parser_parser_ana_w_25_to_mem;  
logic  [39:0] parser_parser_ana_w_26_from_mem;
logic  [54:0] parser_parser_ana_w_26_to_mem;  
logic  [39:0] parser_parser_ana_w_27_from_mem;
logic  [54:0] parser_parser_ana_w_27_to_mem;  
logic  [39:0] parser_parser_ana_w_28_from_mem;
logic  [54:0] parser_parser_ana_w_28_to_mem;  
logic  [39:0] parser_parser_ana_w_29_from_mem;
logic  [54:0] parser_parser_ana_w_29_to_mem;  
logic  [39:0] parser_parser_ana_w_2_from_mem; 
logic  [54:0] parser_parser_ana_w_2_to_mem;   
logic  [39:0] parser_parser_ana_w_30_from_mem;
logic  [54:0] parser_parser_ana_w_30_to_mem;  
logic  [39:0] parser_parser_ana_w_31_from_mem;
logic  [54:0] parser_parser_ana_w_31_to_mem;  
logic  [39:0] parser_parser_ana_w_3_from_mem; 
logic  [54:0] parser_parser_ana_w_3_to_mem;   
logic  [39:0] parser_parser_ana_w_4_from_mem; 
logic  [54:0] parser_parser_ana_w_4_to_mem;   
logic  [39:0] parser_parser_ana_w_5_from_mem; 
logic  [54:0] parser_parser_ana_w_5_to_mem;   
logic  [39:0] parser_parser_ana_w_6_from_mem; 
logic  [54:0] parser_parser_ana_w_6_to_mem;   
logic  [39:0] parser_parser_ana_w_7_from_mem; 
logic  [54:0] parser_parser_ana_w_7_to_mem;   
logic  [39:0] parser_parser_ana_w_8_from_mem; 
logic  [54:0] parser_parser_ana_w_8_to_mem;   
logic  [39:0] parser_parser_ana_w_9_from_mem; 
logic  [54:0] parser_parser_ana_w_9_to_mem;   
logic  [11:0] parser_parser_csum_cfg_0_from_mem;
logic  [28:0] parser_parser_csum_cfg_0_to_mem;
logic  [11:0] parser_parser_csum_cfg_1_from_mem;
logic  [28:0] parser_parser_csum_cfg_1_to_mem;
logic  [88:0] parser_parser_extract_cfg_0_from_mem;
logic [103:0] parser_parser_extract_cfg_0_to_mem;
logic  [88:0] parser_parser_extract_cfg_10_from_mem;
logic [103:0] parser_parser_extract_cfg_10_to_mem;
logic  [88:0] parser_parser_extract_cfg_11_from_mem;
logic [103:0] parser_parser_extract_cfg_11_to_mem;
logic  [88:0] parser_parser_extract_cfg_12_from_mem;
logic [103:0] parser_parser_extract_cfg_12_to_mem;
logic  [88:0] parser_parser_extract_cfg_13_from_mem;
logic [103:0] parser_parser_extract_cfg_13_to_mem;
logic  [88:0] parser_parser_extract_cfg_14_from_mem;
logic [103:0] parser_parser_extract_cfg_14_to_mem;
logic  [88:0] parser_parser_extract_cfg_15_from_mem;
logic [103:0] parser_parser_extract_cfg_15_to_mem;
logic  [88:0] parser_parser_extract_cfg_1_from_mem;
logic [103:0] parser_parser_extract_cfg_1_to_mem;
logic  [88:0] parser_parser_extract_cfg_2_from_mem;
logic [103:0] parser_parser_extract_cfg_2_to_mem;
logic  [88:0] parser_parser_extract_cfg_3_from_mem;
logic [103:0] parser_parser_extract_cfg_3_to_mem;
logic  [88:0] parser_parser_extract_cfg_4_from_mem;
logic [103:0] parser_parser_extract_cfg_4_to_mem;
logic  [88:0] parser_parser_extract_cfg_5_from_mem;
logic [103:0] parser_parser_extract_cfg_5_to_mem;
logic  [88:0] parser_parser_extract_cfg_6_from_mem;
logic [103:0] parser_parser_extract_cfg_6_to_mem;
logic  [88:0] parser_parser_extract_cfg_7_from_mem;
logic [103:0] parser_parser_extract_cfg_7_to_mem;
logic  [88:0] parser_parser_extract_cfg_8_from_mem;
logic [103:0] parser_parser_extract_cfg_8_to_mem;
logic  [88:0] parser_parser_extract_cfg_9_from_mem;
logic [103:0] parser_parser_extract_cfg_9_to_mem;
logic  [39:0] parser_parser_key_s_0_from_mem; 
logic  [54:0] parser_parser_key_s_0_to_mem;   
logic  [39:0] parser_parser_key_s_10_from_mem;
logic  [54:0] parser_parser_key_s_10_to_mem;  
logic  [39:0] parser_parser_key_s_11_from_mem;
logic  [54:0] parser_parser_key_s_11_to_mem;  
logic  [39:0] parser_parser_key_s_12_from_mem;
logic  [54:0] parser_parser_key_s_12_to_mem;  
logic  [39:0] parser_parser_key_s_13_from_mem;
logic  [54:0] parser_parser_key_s_13_to_mem;  
logic  [39:0] parser_parser_key_s_14_from_mem;
logic  [54:0] parser_parser_key_s_14_to_mem;  
logic  [39:0] parser_parser_key_s_15_from_mem;
logic  [54:0] parser_parser_key_s_15_to_mem;  
logic  [39:0] parser_parser_key_s_16_from_mem;
logic  [54:0] parser_parser_key_s_16_to_mem;  
logic  [39:0] parser_parser_key_s_17_from_mem;
logic  [54:0] parser_parser_key_s_17_to_mem;  
logic  [39:0] parser_parser_key_s_18_from_mem;
logic  [54:0] parser_parser_key_s_18_to_mem;  
logic  [39:0] parser_parser_key_s_19_from_mem;
logic  [54:0] parser_parser_key_s_19_to_mem;  
logic  [39:0] parser_parser_key_s_1_from_mem; 
logic  [54:0] parser_parser_key_s_1_to_mem;   
logic  [39:0] parser_parser_key_s_20_from_mem;
logic  [54:0] parser_parser_key_s_20_to_mem;  
logic  [39:0] parser_parser_key_s_21_from_mem;
logic  [54:0] parser_parser_key_s_21_to_mem;  
logic  [39:0] parser_parser_key_s_22_from_mem;
logic  [54:0] parser_parser_key_s_22_to_mem;  
logic  [39:0] parser_parser_key_s_23_from_mem;
logic  [54:0] parser_parser_key_s_23_to_mem;  
logic  [39:0] parser_parser_key_s_24_from_mem;
logic  [54:0] parser_parser_key_s_24_to_mem;  
logic  [39:0] parser_parser_key_s_25_from_mem;
logic  [54:0] parser_parser_key_s_25_to_mem;  
logic  [39:0] parser_parser_key_s_26_from_mem;
logic  [54:0] parser_parser_key_s_26_to_mem;  
logic  [39:0] parser_parser_key_s_27_from_mem;
logic  [54:0] parser_parser_key_s_27_to_mem;  
logic  [39:0] parser_parser_key_s_28_from_mem;
logic  [54:0] parser_parser_key_s_28_to_mem;  
logic  [39:0] parser_parser_key_s_29_from_mem;
logic  [54:0] parser_parser_key_s_29_to_mem;  
logic  [39:0] parser_parser_key_s_2_from_mem; 
logic  [54:0] parser_parser_key_s_2_to_mem;   
logic  [39:0] parser_parser_key_s_30_from_mem;
logic  [54:0] parser_parser_key_s_30_to_mem;  
logic  [39:0] parser_parser_key_s_31_from_mem;
logic  [54:0] parser_parser_key_s_31_to_mem;  
logic  [39:0] parser_parser_key_s_3_from_mem; 
logic  [54:0] parser_parser_key_s_3_to_mem;   
logic  [39:0] parser_parser_key_s_4_from_mem; 
logic  [54:0] parser_parser_key_s_4_to_mem;   
logic  [39:0] parser_parser_key_s_5_from_mem; 
logic  [54:0] parser_parser_key_s_5_to_mem;   
logic  [39:0] parser_parser_key_s_6_from_mem; 
logic  [54:0] parser_parser_key_s_6_to_mem;   
logic  [39:0] parser_parser_key_s_7_from_mem; 
logic  [54:0] parser_parser_key_s_7_to_mem;   
logic  [39:0] parser_parser_key_s_8_from_mem; 
logic  [54:0] parser_parser_key_s_8_to_mem;   
logic  [39:0] parser_parser_key_s_9_from_mem; 
logic  [54:0] parser_parser_key_s_9_to_mem;   
logic  [72:0] parser_parser_key_w_0_from_mem; 
logic  [87:0] parser_parser_key_w_0_to_mem;   
logic  [72:0] parser_parser_key_w_10_from_mem;
logic  [87:0] parser_parser_key_w_10_to_mem;  
logic  [72:0] parser_parser_key_w_11_from_mem;
logic  [87:0] parser_parser_key_w_11_to_mem;  
logic  [72:0] parser_parser_key_w_12_from_mem;
logic  [87:0] parser_parser_key_w_12_to_mem;  
logic  [72:0] parser_parser_key_w_13_from_mem;
logic  [87:0] parser_parser_key_w_13_to_mem;  
logic  [72:0] parser_parser_key_w_14_from_mem;
logic  [87:0] parser_parser_key_w_14_to_mem;  
logic  [72:0] parser_parser_key_w_15_from_mem;
logic  [87:0] parser_parser_key_w_15_to_mem;  
logic  [72:0] parser_parser_key_w_16_from_mem;
logic  [87:0] parser_parser_key_w_16_to_mem;  
logic  [72:0] parser_parser_key_w_17_from_mem;
logic  [87:0] parser_parser_key_w_17_to_mem;  
logic  [72:0] parser_parser_key_w_18_from_mem;
logic  [87:0] parser_parser_key_w_18_to_mem;  
logic  [72:0] parser_parser_key_w_19_from_mem;
logic  [87:0] parser_parser_key_w_19_to_mem;  
logic  [72:0] parser_parser_key_w_1_from_mem; 
logic  [87:0] parser_parser_key_w_1_to_mem;   
logic  [72:0] parser_parser_key_w_20_from_mem;
logic  [87:0] parser_parser_key_w_20_to_mem;  
logic  [72:0] parser_parser_key_w_21_from_mem;
logic  [87:0] parser_parser_key_w_21_to_mem;  
logic  [72:0] parser_parser_key_w_22_from_mem;
logic  [87:0] parser_parser_key_w_22_to_mem;  
logic  [72:0] parser_parser_key_w_23_from_mem;
logic  [87:0] parser_parser_key_w_23_to_mem;  
logic  [72:0] parser_parser_key_w_24_from_mem;
logic  [87:0] parser_parser_key_w_24_to_mem;  
logic  [72:0] parser_parser_key_w_25_from_mem;
logic  [87:0] parser_parser_key_w_25_to_mem;  
logic  [72:0] parser_parser_key_w_26_from_mem;
logic  [87:0] parser_parser_key_w_26_to_mem;  
logic  [72:0] parser_parser_key_w_27_from_mem;
logic  [87:0] parser_parser_key_w_27_to_mem;  
logic  [72:0] parser_parser_key_w_28_from_mem;
logic  [87:0] parser_parser_key_w_28_to_mem;  
logic  [72:0] parser_parser_key_w_29_from_mem;
logic  [87:0] parser_parser_key_w_29_to_mem;  
logic  [72:0] parser_parser_key_w_2_from_mem; 
logic  [87:0] parser_parser_key_w_2_to_mem;   
logic  [72:0] parser_parser_key_w_30_from_mem;
logic  [87:0] parser_parser_key_w_30_to_mem;  
logic  [72:0] parser_parser_key_w_31_from_mem;
logic  [87:0] parser_parser_key_w_31_to_mem;  
logic  [72:0] parser_parser_key_w_3_from_mem; 
logic  [87:0] parser_parser_key_w_3_to_mem;   
logic  [72:0] parser_parser_key_w_4_from_mem; 
logic  [87:0] parser_parser_key_w_4_to_mem;   
logic  [72:0] parser_parser_key_w_5_from_mem; 
logic  [87:0] parser_parser_key_w_5_to_mem;   
logic  [72:0] parser_parser_key_w_6_from_mem; 
logic  [87:0] parser_parser_key_w_6_to_mem;   
logic  [72:0] parser_parser_key_w_7_from_mem; 
logic  [87:0] parser_parser_key_w_7_to_mem;   
logic  [72:0] parser_parser_key_w_8_from_mem; 
logic  [87:0] parser_parser_key_w_8_to_mem;   
logic  [72:0] parser_parser_key_w_9_from_mem; 
logic  [87:0] parser_parser_key_w_9_to_mem;   
logic  [69:0] parser_parser_metadata_fifo_from_mem;
logic  [88:0] parser_parser_metadata_fifo_to_mem;
logic  [72:0] parser_parser_port_cfg_0_from_mem;
logic  [89:0] parser_parser_port_cfg_0_to_mem;
logic  [72:0] parser_parser_port_cfg_1_from_mem;
logic  [89:0] parser_parser_port_cfg_1_to_mem;
logic  [20:0] parser_parser_ptype_ram_from_mem;
logic  [34:0] parser_parser_ptype_ram_to_mem; 
logic reset_n; 
assign reset_n = !reset;


// module parser_shells_wrapper    from parser_shells_wrapper using parser_shells_wrapper.map 
parser_shells_wrapper    parser_shells_wrapper(
/* input  logic          */ .PARSER_ANA_EXT_4_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_4_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_5_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_5_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_6_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_6_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_7_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_7_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_8_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_8_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_9_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_9_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_S_0_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_0_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_10_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_10_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_11_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_11_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_12_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_12_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_13_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_13_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_14_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_14_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_15_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_15_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_16_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_16_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_17_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_17_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_18_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_18_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_19_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_19_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_1_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_1_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_20_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_20_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_21_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_21_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_22_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_22_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_23_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_23_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_24_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_24_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_25_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_25_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_26_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_26_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_27_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_27_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_28_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_28_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_29_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_29_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_2_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_2_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_30_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_30_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_31_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_S_31_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_S_3_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_5_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_5_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_6_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_6_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_7_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_7_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_8_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_8_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_9_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_9_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_0_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_0_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_10_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_10_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_11_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_11_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_12_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_12_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_13_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_13_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_14_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_14_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_15_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_15_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_16_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_16_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_17_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_17_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_18_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_18_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_19_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_19_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_1_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_1_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_20_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_20_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_21_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_21_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_22_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_22_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_23_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_23_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_24_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_24_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_25_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_25_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_26_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_26_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_27_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_27_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_28_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_28_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_29_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_29_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_2_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_2_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_30_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_30_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_31_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_ANA_W_31_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_ANA_W_3_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_3_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_4_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_4_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_5_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_5_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_6_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_6_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_7_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_7_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_8_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_8_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_W_9_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_W_9_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_CSUM_CFG_0_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_CSUM_CFG_0_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_CSUM_CFG_1_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_CSUM_CFG_1_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ECC_COR_ERR_reg_sel            (),                                                
/* input  logic          */ .PARSER_ECC_UNCOR_ERR_reg_sel          (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_0_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_0_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_10_CFG_reg_sel     (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_10_STATUS_reg_sel  (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_11_CFG_reg_sel     (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_11_STATUS_reg_sel  (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_12_CFG_reg_sel     (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_12_STATUS_reg_sel  (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_13_CFG_reg_sel     (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_13_STATUS_reg_sel  (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_14_CFG_reg_sel     (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_14_STATUS_reg_sel  (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_15_CFG_reg_sel     (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_15_STATUS_reg_sel  (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_1_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_1_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_2_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_2_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_3_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_3_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_4_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_4_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_5_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_5_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_6_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_6_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_7_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_7_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_8_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_8_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_9_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_EXTRACT_CFG_9_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_KEY_S_0_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_0_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_10_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_10_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_11_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_11_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_12_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_12_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_13_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_13_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_14_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_14_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_15_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_15_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_16_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_16_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_17_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_17_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_18_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_18_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_19_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_19_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_1_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_1_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_20_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_20_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_21_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_21_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_22_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_22_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_23_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_23_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_24_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_24_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_25_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_25_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_26_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_26_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_27_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_27_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_28_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_28_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_29_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_29_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_2_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_2_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_30_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_30_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_31_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_S_31_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_S_3_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_3_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_4_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_4_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_5_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_5_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_6_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_8_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_9_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_9_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_0_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_0_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_10_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_10_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_11_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_11_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_12_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_12_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_13_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_13_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_14_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_14_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_15_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_15_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_16_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_16_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_17_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_17_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_18_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_18_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_19_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_19_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_1_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_1_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_20_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_20_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_21_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_21_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_22_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_22_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_23_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_23_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_24_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_24_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_25_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_25_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_26_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_26_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_27_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_27_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_28_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_28_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_29_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_29_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_2_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_2_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_30_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_30_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_31_CFG_reg_sel           (),                                                
/* input  logic          */ .PARSER_KEY_W_31_STATUS_reg_sel        (),                                                
/* input  logic          */ .PARSER_KEY_W_3_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_3_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_4_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_4_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_5_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_5_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_6_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_6_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_7_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_7_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_8_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_8_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_W_9_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_W_9_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_METADATA_FIFO_CFG_reg_sel      (),                                                
/* input  logic          */ .PARSER_METADATA_FIFO_STATUS_reg_sel   (),                                                
/* input  logic          */ .PARSER_PORT_CFG_0_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_PORT_CFG_0_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_PORT_CFG_1_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_PORT_CFG_1_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_PTYPE_RAM_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_PTYPE_RAM_STATUS_reg_sel       (),                                                
/* input  logic          */ .clk                                   (cclk),                                            
/* input  logic          */ .parser_ana_cam_0_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_0_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_0_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_0_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_0_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_0_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_10_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_10_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_10_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_30_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_30_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_30_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_30_wr_data             (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_11_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_11_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_11_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_11_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_11_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_12_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_12_rd_adr              (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_31_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_31_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_31_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_3_mem_ls_enter         (),                                                
/* input  logic          */ .parser_ana_cam_12_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_12_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_12_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_12_wr_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_3_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_3_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_3_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_3_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_13_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_13_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_13_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_13_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_13_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_13_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_14_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_14_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_14_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_14_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_14_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_14_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_15_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_15_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_15_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_15_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_15_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_15_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_16_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_16_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_16_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_16_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_16_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_16_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_17_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_17_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_17_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_17_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_17_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_17_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_18_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_18_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_18_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_18_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_18_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_18_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_19_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_19_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_19_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_19_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_19_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_19_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_1_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_1_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_1_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_1_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_1_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_1_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_20_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_20_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_20_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_20_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_20_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_20_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_21_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_21_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_21_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_21_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_21_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_21_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_22_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_22_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_22_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_22_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_22_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_22_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_23_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_23_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_23_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_24_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_24_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_24_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_24_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_24_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_25_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_25_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_25_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_25_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_25_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_25_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_26_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_26_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_26_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_26_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_26_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_26_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_27_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_27_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_27_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_27_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_27_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_27_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_28_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_28_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_28_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_28_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_28_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_28_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_29_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_29_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_29_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_29_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_29_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_29_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_2_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_2_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_2_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_2_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_2_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_2_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_30_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_30_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_30_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_30_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_30_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_30_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_31_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_31_rd_adr              (),                                                
/* input  logic          */ .parser_ana_cam_31_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_31_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_31_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_31_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_3_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_3_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_3_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_3_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_3_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_3_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_4_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_4_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_4_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_4_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_4_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_4_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_5_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_5_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_5_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_5_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_5_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_5_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_6_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_6_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_6_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_6_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_6_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_6_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_7_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_7_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_7_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_7_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_7_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_7_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_8_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_8_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_8_wr_en                (),                                                
/* input  logic          */ .parser_ana_cam_9_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_9_rd_adr               (),                                                
/* input  logic          */ .parser_ana_cam_9_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_9_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_9_wr_data              (),                                                
/* input  logic          */ .parser_ana_cam_9_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_0_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_0_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_0_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_0_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_0_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_0_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_10_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_10_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_10_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_10_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_10_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_10_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_11_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_11_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_11_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_11_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_11_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_11_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_12_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_12_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_12_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_12_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_12_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_12_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_13_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_13_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_13_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_13_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_13_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_13_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_14_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_14_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_14_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_14_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_14_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_14_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_15_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_15_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_15_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_15_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_15_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_15_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_16_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_16_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_16_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_16_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_16_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_16_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_17_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_17_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_17_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_17_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_17_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_17_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_18_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_18_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_18_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_18_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_18_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_18_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_19_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_19_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_19_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_19_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_19_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_19_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_1_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_1_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_1_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_1_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_1_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_1_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_20_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_20_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_21_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_21_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_21_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_21_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_21_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_21_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_22_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_22_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_22_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_22_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_22_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_22_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_23_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_23_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_23_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_23_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_23_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_23_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_24_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_24_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_24_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_24_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_24_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_24_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_25_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_25_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_25_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_25_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_25_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_25_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_26_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_26_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_26_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_26_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_26_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_26_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_27_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_27_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_27_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_27_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_27_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_27_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_28_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_28_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_28_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_28_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_28_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_28_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_29_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_29_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_29_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_29_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_29_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_29_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_2_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_2_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_2_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_2_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_2_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_2_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_30_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_30_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_30_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_30_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_30_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_30_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_31_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_31_rd_adr              (),                                                
/* input  logic          */ .parser_ana_exc_31_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_31_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_31_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_31_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_3_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_3_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_3_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_3_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_3_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_3_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_4_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_4_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_4_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_4_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_4_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_4_wr_en                (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_5_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_5_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_6_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_6_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_6_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_6_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_6_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_6_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_7_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_7_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_7_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_7_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_7_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_7_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_8_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_8_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_8_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_8_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_8_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_8_wr_en                (),                                                
/* input  logic          */ .parser_ana_exc_9_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_9_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_9_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_9_wr_adr               (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_9_wr_data              (),                                                
/* input  logic          */ .parser_ana_exc_9_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_0_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_0_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_0_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_0_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_0_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_0_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_10_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_10_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_10_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_10_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_10_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_10_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_11_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_11_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_11_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_11_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_11_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_11_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_12_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_12_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_12_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_12_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_12_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_12_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_13_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_13_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_13_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_13_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_13_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_13_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_14_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_14_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_14_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_14_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_14_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_14_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_15_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_15_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_15_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_15_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_15_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_15_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_16_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_16_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_16_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_16_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_16_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_16_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_17_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_17_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_17_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_17_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_17_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_17_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_18_mem_ls_enter        (),                                                
/* input  logic          */ .parser_ana_ext_18_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_19_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_19_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_19_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_19_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_19_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_19_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_1_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_1_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_1_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_1_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_1_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_1_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_20_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_20_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_20_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_20_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_20_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_20_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_21_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_21_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_21_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_21_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_21_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_21_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_22_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_22_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_22_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_22_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_22_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_22_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_23_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_23_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_23_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_23_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_23_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_23_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_24_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_24_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_24_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_24_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_24_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_24_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_25_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_25_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_25_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_25_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_25_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_25_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_26_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_26_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_26_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_26_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_26_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_26_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_27_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_27_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_27_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_27_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_27_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_27_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_28_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_28_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_28_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_28_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_28_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_28_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_29_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_29_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_29_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_29_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_29_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_29_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_2_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_2_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_2_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_2_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_2_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_2_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_30_mem_ls_enter        (),                                                
/* input  logic   [32:0] */ .parser_parser_ana_ext_5_from_mem      (parser_parser_ana_ext_5_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_6_from_mem      (parser_parser_ana_ext_6_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_7_from_mem      (parser_parser_ana_ext_7_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_8_from_mem      (parser_parser_ana_ext_8_from_mem),                
/* input  logic   [55:0] */ .parser_parser_ana_s_12_from_mem       (parser_parser_ana_s_12_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_13_from_mem       (parser_parser_ana_s_13_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_14_from_mem       (parser_parser_ana_s_14_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_15_from_mem       (parser_parser_ana_s_15_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_16_from_mem       (parser_parser_ana_s_16_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_17_from_mem       (parser_parser_ana_s_17_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_18_from_mem       (parser_parser_ana_s_18_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_19_from_mem       (parser_parser_ana_s_19_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_1_from_mem        (parser_parser_ana_s_1_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_20_from_mem       (parser_parser_ana_s_20_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_21_from_mem       (parser_parser_ana_s_21_from_mem),                 
/* input  logic          */ .parser_ana_ext_3_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_4_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_4_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_4_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_4_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_4_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_4_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_5_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_5_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_5_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_5_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_5_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_5_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_6_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_6_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_6_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_6_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_6_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_6_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_7_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_7_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_7_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_7_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_7_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_7_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_8_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_8_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_8_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_8_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_8_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_8_wr_en                (),                                                
/* input  logic          */ .parser_ana_ext_9_mem_ls_enter         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_9_rd_adr               (),                                                
/* input  logic          */ .parser_ana_ext_9_rd_en                (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_9_wr_adr               (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_9_wr_data              (),                                                
/* input  logic          */ .parser_ana_ext_9_wr_en                (),                                                
/* input  logic          */ .parser_ana_s_0_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_0_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_0_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_0_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_0_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_0_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_10_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_10_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_10_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_10_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_10_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_10_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_11_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_11_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_11_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_11_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_11_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_11_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_12_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_12_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_12_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_12_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_12_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_12_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_13_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_13_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_13_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_13_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_13_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_13_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_14_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_14_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_14_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_14_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_14_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_14_wr_en                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_15_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_15_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_16_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_16_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_16_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_16_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_16_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_16_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_17_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_17_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_17_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_17_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_17_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_17_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_18_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_18_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_18_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_18_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_18_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_18_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_19_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_19_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_19_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_19_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_19_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_19_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_1_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_1_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_1_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_1_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_1_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_1_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_20_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_20_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_20_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_20_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_20_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_20_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_21_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_21_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_21_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_21_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_21_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_21_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_22_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_22_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_22_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_22_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_22_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_22_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_23_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_23_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_23_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_23_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_23_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_23_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_24_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_24_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_24_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_24_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_24_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_24_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_25_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_25_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_25_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_25_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_25_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_25_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_26_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_26_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_26_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_26_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_26_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_26_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_27_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_27_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_27_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_27_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_27_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_27_wr_en                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_28_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_28_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_29_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_29_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_29_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_29_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_29_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_29_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_2_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_2_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_2_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_2_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_2_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_2_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_30_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_30_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_30_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_30_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_30_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_30_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_31_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_31_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_31_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_31_wr_adr                (),                                                
/* input  logic   [47:0] */ .parser_ana_s_31_wr_data               (),                                                
/* input  logic          */ .parser_ana_s_31_wr_en                 (),                                                
/* input  logic          */ .parser_ana_s_3_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_3_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_3_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_3_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_3_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_3_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_4_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_4_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_4_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_4_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_4_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_4_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_5_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_5_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_5_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_5_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_5_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_5_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_6_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_6_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_6_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_6_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_6_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_6_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_7_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_7_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_7_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_7_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_7_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_7_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_8_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_8_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_8_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_8_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_8_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_8_wr_en                  (),                                                
/* input  logic          */ .parser_ana_s_9_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_s_9_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_s_9_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_s_9_wr_adr                 (),                                                
/* input  logic   [47:0] */ .parser_ana_s_9_wr_data                (),                                                
/* input  logic          */ .parser_ana_s_9_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_0_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_0_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_0_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_0_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_0_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_0_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_10_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_10_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_10_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_10_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_10_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_10_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_11_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_11_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_11_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_11_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_11_wr_data               (),                                                
/* input  logic    [3:0] */ .parser_ana_w_12_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_12_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_12_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_13_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_13_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_13_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_13_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_13_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_13_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_14_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_14_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_14_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_14_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_14_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_14_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_15_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_15_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_15_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_15_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_15_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_15_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_16_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_16_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_16_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_16_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_16_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_16_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_17_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_17_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_17_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_17_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_17_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_17_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_18_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_18_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_18_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_18_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_18_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_18_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_19_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_19_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_19_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_19_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_19_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_19_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_1_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_1_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_1_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_1_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_1_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_1_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_20_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_20_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_20_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_20_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_20_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_20_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_21_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_21_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_21_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_21_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_21_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_21_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_22_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_22_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_22_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_22_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_22_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_22_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_23_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_23_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_23_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_23_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_23_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_23_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_24_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_24_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_24_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_24_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_24_wr_data               (),                                                
/* input  logic    [3:0] */ .parser_ana_w_25_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_25_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_25_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_26_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_26_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_26_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_26_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_26_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_26_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_27_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_27_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_27_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_27_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_27_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_27_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_28_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_28_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_28_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_28_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_28_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_28_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_29_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_29_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_29_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_29_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_29_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_29_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_2_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_2_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_2_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_2_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_2_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_2_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_30_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_30_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_30_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_30_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_30_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_30_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_31_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_31_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_31_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_w_31_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_ana_w_31_wr_data               (),                                                
/* input  logic          */ .parser_ana_w_31_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_3_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_3_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_3_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_3_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_3_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_3_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_4_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_4_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_4_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_4_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_4_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_4_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_5_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_5_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_5_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_5_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_5_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_5_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_6_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_6_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_6_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_6_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_6_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_6_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_7_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_7_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_7_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_7_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_7_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_7_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_8_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_8_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_8_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_8_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_8_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_8_wr_en                  (),                                                
/* input  logic          */ .parser_ana_w_9_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_ana_w_9_rd_adr                 (),                                                
/* input  logic          */ .parser_ana_w_9_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_ana_w_9_wr_adr                 (),                                                
/* input  logic    [4:0] */ .parser_csum_cfg_0_rd_adr              (),                                                
/* input  logic          */ .parser_csum_cfg_0_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_csum_cfg_0_wr_adr              (),                                                
/* input  logic    [5:0] */ .parser_csum_cfg_0_wr_data             (),                                                
/* input  logic          */ .parser_csum_cfg_0_wr_en               (),                                                
/* input  logic          */ .parser_csum_cfg_1_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_csum_cfg_1_rd_adr              (),                                                
/* input  logic          */ .parser_csum_cfg_1_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_csum_cfg_1_wr_adr              (),                                                
/* input  logic    [5:0] */ .parser_csum_cfg_1_wr_data             (),                                                
/* input  logic          */ .parser_csum_cfg_1_wr_en               (),                                                
/* input  logic          */ .parser_extract_cfg_0_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_0_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_0_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_0_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_0_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_0_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_10_mem_ls_enter    (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_10_rd_adr          (),                                                
/* input  logic          */ .parser_extract_cfg_10_rd_en           (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_10_wr_adr          (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_10_wr_data         (),                                                
/* input  logic          */ .parser_extract_cfg_10_wr_en           (),                                                
/* input  logic          */ .parser_extract_cfg_11_mem_ls_enter    (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_11_rd_adr          (),                                                
/* input  logic          */ .parser_extract_cfg_11_rd_en           (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_11_wr_adr          (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_11_wr_data         (),                                                
/* input  logic          */ .parser_extract_cfg_11_wr_en           (),                                                
/* input  logic          */ .parser_extract_cfg_12_mem_ls_enter    (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_12_rd_adr          (),                                                
/* input  logic          */ .parser_extract_cfg_12_rd_en           (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_12_wr_adr          (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_12_wr_data         (),                                                
/* input  logic          */ .parser_extract_cfg_12_wr_en           (),                                                
/* input  logic          */ .parser_extract_cfg_13_mem_ls_enter    (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_13_rd_adr          (),                                                
/* input  logic          */ .parser_extract_cfg_13_rd_en           (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_13_wr_adr          (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_13_wr_data         (),                                                
/* input  logic          */ .parser_extract_cfg_13_wr_en           (),                                                
/* input  logic          */ .parser_extract_cfg_14_mem_ls_enter    (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_14_rd_adr          (),                                                
/* input  logic          */ .parser_extract_cfg_14_rd_en           (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_14_wr_adr          (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_14_wr_data         (),                                                
/* input  logic          */ .parser_extract_cfg_14_wr_en           (),                                                
/* input  logic          */ .parser_extract_cfg_15_mem_ls_enter    (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_15_rd_adr          (),                                                
/* input  logic          */ .parser_extract_cfg_15_rd_en           (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_15_wr_adr          (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_15_wr_data         (),                                                
/* input  logic          */ .parser_extract_cfg_15_wr_en           (),                                                
/* input  logic          */ .parser_extract_cfg_1_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_1_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_1_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_1_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_1_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_1_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_2_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_2_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_2_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_2_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_2_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_2_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_3_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_3_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_3_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_3_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_3_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_3_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_4_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_4_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_4_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_4_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_4_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_4_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_5_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_5_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_5_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_5_wr_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_6_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_6_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_6_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_6_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_7_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_7_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_7_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_7_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_7_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_7_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_8_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_8_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_8_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_8_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_8_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_8_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_9_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_9_rd_adr           (),                                                
/* input  logic          */ .parser_extract_cfg_9_rd_en            (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_9_wr_adr           (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_9_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_9_wr_en            (),                                                
/* input  logic          */ .parser_key_s_0_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_0_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_0_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_0_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_0_wr_data                (),                                                
/* input  logic          */ .parser_key_s_0_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_10_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_10_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_10_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_10_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_10_wr_data               (),                                                
/* input  logic          */ .parser_key_s_10_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_11_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_11_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_11_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_11_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_11_wr_data               (),                                                
/* input  logic          */ .parser_key_s_11_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_12_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_12_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_12_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_12_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_12_wr_data               (),                                                
/* input  logic          */ .parser_key_s_12_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_13_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_13_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_13_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_13_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_13_wr_data               (),                                                
/* input  logic          */ .parser_key_s_13_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_14_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_14_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_14_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_14_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_14_wr_data               (),                                                
/* input  logic          */ .parser_key_s_14_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_15_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_15_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_15_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_15_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_15_wr_data               (),                                                
/* input  logic          */ .parser_key_s_15_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_16_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_16_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_16_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_16_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_16_wr_data               (),                                                
/* input  logic          */ .parser_key_s_16_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_17_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_17_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_17_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_17_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_17_wr_data               (),                                                
/* input  logic          */ .parser_key_s_17_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_18_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_18_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_18_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_18_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_18_wr_data               (),                                                
/* input  logic          */ .parser_key_s_18_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_19_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_19_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_1_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_1_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_1_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_1_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_1_wr_data                (),                                                
/* input  logic          */ .parser_key_s_1_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_20_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_20_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_20_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_20_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_20_wr_data               (),                                                
/* input  logic          */ .parser_key_s_20_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_21_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_21_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_21_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_21_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_21_wr_data               (),                                                
/* input  logic          */ .parser_key_s_21_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_22_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_22_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_22_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_22_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_22_wr_data               (),                                                
/* input  logic          */ .parser_key_s_22_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_23_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_23_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_23_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_23_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_23_wr_data               (),                                                
/* input  logic          */ .parser_key_s_23_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_24_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_24_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_24_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_24_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_24_wr_data               (),                                                
/* input  logic          */ .parser_key_s_24_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_25_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_25_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_25_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_25_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_25_wr_data               (),                                                
/* input  logic          */ .parser_key_s_25_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_26_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_26_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_26_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_26_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_26_wr_data               (),                                                
/* input  logic          */ .parser_key_s_26_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_27_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_27_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_27_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_27_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_27_wr_data               (),                                                
/* input  logic          */ .parser_key_s_27_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_28_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_28_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_28_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_28_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_28_wr_data               (),                                                
/* input  logic          */ .parser_key_s_28_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_29_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_29_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_29_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_29_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_29_wr_data               (),                                                
/* input  logic          */ .parser_key_s_29_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_2_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_2_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_2_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_2_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_2_wr_data                (),                                                
/* input  logic          */ .parser_key_s_2_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_30_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_30_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_30_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_30_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_30_wr_data               (),                                                
/* input  logic          */ .parser_key_s_30_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_31_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_s_31_rd_adr                (),                                                
/* input  logic          */ .parser_key_s_31_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_3_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_3_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_3_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_3_wr_data                (),                                                
/* input  logic          */ .parser_key_s_3_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_4_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_4_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_4_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_4_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_4_wr_data                (),                                                
/* input  logic          */ .parser_key_s_4_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_5_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_5_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_5_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_5_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_5_wr_data                (),                                                
/* input  logic          */ .parser_key_s_5_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_6_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_6_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_6_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_6_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_6_wr_data                (),                                                
/* input  logic          */ .parser_key_s_6_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_7_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_7_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_7_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_7_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_7_wr_data                (),                                                
/* input  logic          */ .parser_key_s_7_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_8_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_8_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_8_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_8_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_8_wr_data                (),                                                
/* input  logic          */ .parser_key_s_8_wr_en                  (),                                                
/* input  logic          */ .parser_key_s_9_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_s_9_rd_adr                 (),                                                
/* input  logic          */ .parser_key_s_9_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_s_9_wr_adr                 (),                                                
/* input  logic   [31:0] */ .parser_key_s_9_wr_data                (),                                                
/* input  logic          */ .parser_key_s_9_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_0_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_0_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_0_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_0_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_0_wr_data                (),                                                
/* input  logic          */ .parser_key_w_0_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_10_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_10_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_10_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_10_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_10_wr_data               (),                                                
/* input  logic          */ .parser_key_w_10_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_11_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_11_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_11_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_11_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_11_wr_data               (),                                                
/* input  logic          */ .parser_key_w_11_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_12_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_12_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_12_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_12_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_12_wr_data               (),                                                
/* input  logic          */ .parser_key_w_12_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_13_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_13_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_13_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_13_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_13_wr_data               (),                                                
/* input  logic          */ .parser_key_w_13_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_14_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_14_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_14_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_14_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_14_wr_data               (),                                                
/* input  logic          */ .parser_key_w_14_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_15_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_15_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_15_rd_en                 (),                                                
/* input  logic          */ .parser_key_w_16_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_17_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_17_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_17_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_17_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_17_wr_data               (),                                                
/* input  logic          */ .parser_key_w_17_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_18_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_18_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_18_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_18_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_18_wr_data               (),                                                
/* input  logic   [63:0] */ .parser_key_w_1_wr_data                (),                                                
/* input  logic          */ .parser_key_w_1_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_20_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_20_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_20_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_20_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_20_wr_data               (),                                                
/* input  logic          */ .parser_key_w_20_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_21_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_21_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_21_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_21_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_21_wr_data               (),                                                
/* input  logic          */ .parser_key_w_21_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_22_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_22_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_22_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_22_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_22_wr_data               (),                                                
/* input  logic          */ .parser_key_w_22_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_23_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_23_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_23_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_23_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_23_wr_data               (),                                                
/* input  logic          */ .parser_key_w_23_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_24_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_24_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_24_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_24_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_24_wr_data               (),                                                
/* input  logic          */ .parser_key_w_24_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_25_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_25_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_25_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_25_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_25_wr_data               (),                                                
/* input  logic          */ .parser_key_w_25_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_26_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_26_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_26_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_26_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_26_wr_data               (),                                                
/* input  logic          */ .parser_key_w_26_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_27_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_27_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_27_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_27_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_27_wr_data               (),                                                
/* input  logic          */ .parser_key_w_27_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_28_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_28_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_28_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_28_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_28_wr_data               (),                                                
/* input  logic          */ .parser_key_w_28_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_29_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_29_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_2_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_2_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_2_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_2_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_2_wr_data                (),                                                
/* input  logic          */ .parser_key_w_2_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_30_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_30_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_30_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_30_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_30_wr_data               (),                                                
/* input  logic          */ .parser_key_w_30_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_31_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_31_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_31_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_31_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_31_wr_data               (),                                                
/* input  logic          */ .parser_key_w_31_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_3_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_3_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_3_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_3_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_3_wr_data                (),                                                
/* input  logic          */ .parser_key_w_3_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_4_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_4_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_4_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_4_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_4_wr_data                (),                                                
/* input  logic          */ .parser_key_w_4_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_5_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_5_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_5_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_5_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_5_wr_data                (),                                                
/* input  logic          */ .parser_key_w_5_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_6_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_6_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_6_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_6_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_6_wr_data                (),                                                
/* input  logic          */ .parser_key_w_6_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_7_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_7_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_7_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_7_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_7_wr_data                (),                                                
/* input  logic          */ .parser_key_w_7_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_8_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_8_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_8_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_8_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_8_wr_data                (),                                                
/* input  logic          */ .parser_key_w_8_wr_en                  (),                                                
/* input  logic          */ .parser_key_w_9_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_9_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_9_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_9_wr_adr                 (),                                                
/* input  logic   [63:0] */ .parser_key_w_9_wr_data                (),                                                
/* input  logic          */ .parser_key_w_9_wr_en                  (),                                                
/* input  logic          */ .parser_metadata_fifo_mem_ls_enter     (),                                                
/* input  logic    [5:0] */ .parser_metadata_fifo_rd_adr           (),                                                
/* input  logic          */ .parser_metadata_fifo_rd_en            (),                                                
/* input  logic    [5:0] */ .parser_metadata_fifo_wr_adr           (),                                                
/* input  logic   [60:0] */ .parser_metadata_fifo_wr_data          (),                                                
/* input  logic          */ .parser_metadata_fifo_wr_en            (),                                                
/* input  logic  [104:0] */ .parser_parser_ana_cam_0_from_mem      (parser_parser_ana_cam_0_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_10_from_mem     (parser_parser_ana_cam_10_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_11_from_mem     (parser_parser_ana_cam_11_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_12_from_mem     (parser_parser_ana_cam_12_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_13_from_mem     (parser_parser_ana_cam_13_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_14_from_mem     (parser_parser_ana_cam_14_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_15_from_mem     (parser_parser_ana_cam_15_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_16_from_mem     (parser_parser_ana_cam_16_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_17_from_mem     (parser_parser_ana_cam_17_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_18_from_mem     (parser_parser_ana_cam_18_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_19_from_mem     (parser_parser_ana_cam_19_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_1_from_mem      (parser_parser_ana_cam_1_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_20_from_mem     (parser_parser_ana_cam_20_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_21_from_mem     (parser_parser_ana_cam_21_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_22_from_mem     (parser_parser_ana_cam_22_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_23_from_mem     (parser_parser_ana_cam_23_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_24_from_mem     (parser_parser_ana_cam_24_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_25_from_mem     (parser_parser_ana_cam_25_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_26_from_mem     (parser_parser_ana_cam_26_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_27_from_mem     (parser_parser_ana_cam_27_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_28_from_mem     (parser_parser_ana_cam_28_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_29_from_mem     (parser_parser_ana_cam_29_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_4_from_mem      (parser_parser_ana_cam_4_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_5_from_mem      (parser_parser_ana_cam_5_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_6_from_mem      (parser_parser_ana_cam_6_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_7_from_mem      (parser_parser_ana_cam_7_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_8_from_mem      (parser_parser_ana_cam_8_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_9_from_mem      (parser_parser_ana_cam_9_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_0_from_mem      (parser_parser_ana_exc_0_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_10_from_mem     (parser_parser_ana_exc_10_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_11_from_mem     (parser_parser_ana_exc_11_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_12_from_mem     (parser_parser_ana_exc_12_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_13_from_mem     (parser_parser_ana_exc_13_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_14_from_mem     (parser_parser_ana_exc_14_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_15_from_mem     (parser_parser_ana_exc_15_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_16_from_mem     (parser_parser_ana_exc_16_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_17_from_mem     (parser_parser_ana_exc_17_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_18_from_mem     (parser_parser_ana_exc_18_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_19_from_mem     (parser_parser_ana_exc_19_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_1_from_mem      (parser_parser_ana_exc_1_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_20_from_mem     (parser_parser_ana_exc_20_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_21_from_mem     (parser_parser_ana_exc_21_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_22_from_mem     (parser_parser_ana_exc_22_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_23_from_mem     (parser_parser_ana_exc_23_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_24_from_mem     (parser_parser_ana_exc_24_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_25_from_mem     (parser_parser_ana_exc_25_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_26_from_mem     (parser_parser_ana_exc_26_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_27_from_mem     (parser_parser_ana_exc_27_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_28_from_mem     (parser_parser_ana_exc_28_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_29_from_mem     (parser_parser_ana_exc_29_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_2_from_mem      (parser_parser_ana_exc_2_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_30_from_mem     (parser_parser_ana_exc_30_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_31_from_mem     (parser_parser_ana_exc_31_from_mem),               
/* input  logic   [14:0] */ .parser_parser_ana_exc_3_from_mem      (parser_parser_ana_exc_3_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_4_from_mem      (parser_parser_ana_exc_4_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_5_from_mem      (parser_parser_ana_exc_5_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_6_from_mem      (parser_parser_ana_exc_6_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_7_from_mem      (parser_parser_ana_exc_7_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_8_from_mem      (parser_parser_ana_exc_8_from_mem),                
/* input  logic   [14:0] */ .parser_parser_ana_exc_9_from_mem      (parser_parser_ana_exc_9_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_0_from_mem      (parser_parser_ana_ext_0_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_10_from_mem     (parser_parser_ana_ext_10_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_11_from_mem     (parser_parser_ana_ext_11_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_12_from_mem     (parser_parser_ana_ext_12_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_13_from_mem     (parser_parser_ana_ext_13_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_14_from_mem     (parser_parser_ana_ext_14_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_15_from_mem     (parser_parser_ana_ext_15_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_16_from_mem     (parser_parser_ana_ext_16_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_17_from_mem     (parser_parser_ana_ext_17_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_18_from_mem     (parser_parser_ana_ext_18_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_19_from_mem     (parser_parser_ana_ext_19_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_1_from_mem      (parser_parser_ana_ext_1_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_20_from_mem     (parser_parser_ana_ext_20_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_21_from_mem     (parser_parser_ana_ext_21_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_22_from_mem     (parser_parser_ana_ext_22_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_23_from_mem     (parser_parser_ana_ext_23_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_24_from_mem     (parser_parser_ana_ext_24_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_25_from_mem     (parser_parser_ana_ext_25_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_26_from_mem     (parser_parser_ana_ext_26_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_27_from_mem     (parser_parser_ana_ext_27_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_28_from_mem     (parser_parser_ana_ext_28_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_29_from_mem     (parser_parser_ana_ext_29_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_2_from_mem      (parser_parser_ana_ext_2_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_30_from_mem     (parser_parser_ana_ext_30_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_31_from_mem     (parser_parser_ana_ext_31_from_mem),               
/* input  logic   [32:0] */ .parser_parser_ana_ext_3_from_mem      (parser_parser_ana_ext_3_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_4_from_mem      (parser_parser_ana_ext_4_from_mem),                
/* input  logic   [32:0] */ .parser_parser_ana_ext_9_from_mem      (parser_parser_ana_ext_9_from_mem),                
/* input  logic   [55:0] */ .parser_parser_ana_s_0_from_mem        (parser_parser_ana_s_0_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_10_from_mem       (parser_parser_ana_s_10_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_11_from_mem       (parser_parser_ana_s_11_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_22_from_mem       (parser_parser_ana_s_22_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_23_from_mem       (parser_parser_ana_s_23_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_24_from_mem       (parser_parser_ana_s_24_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_25_from_mem       (parser_parser_ana_s_25_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_26_from_mem       (parser_parser_ana_s_26_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_27_from_mem       (parser_parser_ana_s_27_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_28_from_mem       (parser_parser_ana_s_28_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_29_from_mem       (parser_parser_ana_s_29_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_2_from_mem        (parser_parser_ana_s_2_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_30_from_mem       (parser_parser_ana_s_30_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_31_from_mem       (parser_parser_ana_s_31_from_mem),                 
/* input  logic   [55:0] */ .parser_parser_ana_s_3_from_mem        (parser_parser_ana_s_3_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_4_from_mem        (parser_parser_ana_s_4_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_5_from_mem        (parser_parser_ana_s_5_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_6_from_mem        (parser_parser_ana_s_6_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_7_from_mem        (parser_parser_ana_s_7_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_8_from_mem        (parser_parser_ana_s_8_from_mem),                  
/* input  logic   [55:0] */ .parser_parser_ana_s_9_from_mem        (parser_parser_ana_s_9_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_0_from_mem        (parser_parser_ana_w_0_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_10_from_mem       (parser_parser_ana_w_10_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_11_from_mem       (parser_parser_ana_w_11_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_12_from_mem       (parser_parser_ana_w_12_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_13_from_mem       (parser_parser_ana_w_13_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_14_from_mem       (parser_parser_ana_w_14_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_15_from_mem       (parser_parser_ana_w_15_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_16_from_mem       (parser_parser_ana_w_16_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_17_from_mem       (parser_parser_ana_w_17_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_18_from_mem       (parser_parser_ana_w_18_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_19_from_mem       (parser_parser_ana_w_19_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_1_from_mem        (parser_parser_ana_w_1_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_20_from_mem       (parser_parser_ana_w_20_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_21_from_mem       (parser_parser_ana_w_21_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_22_from_mem       (parser_parser_ana_w_22_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_23_from_mem       (parser_parser_ana_w_23_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_24_from_mem       (parser_parser_ana_w_24_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_25_from_mem       (parser_parser_ana_w_25_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_26_from_mem       (parser_parser_ana_w_26_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_27_from_mem       (parser_parser_ana_w_27_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_28_from_mem       (parser_parser_ana_w_28_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_29_from_mem       (parser_parser_ana_w_29_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_2_from_mem        (parser_parser_ana_w_2_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_30_from_mem       (parser_parser_ana_w_30_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_6_from_mem        (parser_parser_ana_w_6_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_7_from_mem        (parser_parser_ana_w_7_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_8_from_mem        (parser_parser_ana_w_8_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_9_from_mem        (parser_parser_ana_w_9_from_mem),                  
/* input  logic   [11:0] */ .parser_parser_csum_cfg_0_from_mem     (parser_parser_csum_cfg_0_from_mem),               
/* input  logic   [11:0] */ .parser_parser_csum_cfg_1_from_mem     (parser_parser_csum_cfg_1_from_mem),               
/* input  logic   [88:0] */ .parser_parser_extract_cfg_0_from_mem  (parser_parser_extract_cfg_0_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_10_from_mem (parser_parser_extract_cfg_10_from_mem),           
/* input  logic   [88:0] */ .parser_parser_extract_cfg_11_from_mem (parser_parser_extract_cfg_11_from_mem),           
/* input  logic   [88:0] */ .parser_parser_extract_cfg_12_from_mem (parser_parser_extract_cfg_12_from_mem),           
/* input  logic   [88:0] */ .parser_parser_extract_cfg_13_from_mem (parser_parser_extract_cfg_13_from_mem),           
/* input  logic   [88:0] */ .parser_parser_extract_cfg_14_from_mem (parser_parser_extract_cfg_14_from_mem),           
/* input  logic   [88:0] */ .parser_parser_extract_cfg_15_from_mem (parser_parser_extract_cfg_15_from_mem),           
/* input  logic   [88:0] */ .parser_parser_extract_cfg_1_from_mem  (parser_parser_extract_cfg_1_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_2_from_mem  (parser_parser_extract_cfg_2_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_3_from_mem  (parser_parser_extract_cfg_3_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_4_from_mem  (parser_parser_extract_cfg_4_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_5_from_mem  (parser_parser_extract_cfg_5_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_6_from_mem  (parser_parser_extract_cfg_6_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_7_from_mem  (parser_parser_extract_cfg_7_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_8_from_mem  (parser_parser_extract_cfg_8_from_mem),            
/* input  logic   [88:0] */ .parser_parser_extract_cfg_9_from_mem  (parser_parser_extract_cfg_9_from_mem),            
/* input  logic   [39:0] */ .parser_parser_key_s_0_from_mem        (parser_parser_key_s_0_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_10_from_mem       (parser_parser_key_s_10_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_11_from_mem       (parser_parser_key_s_11_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_12_from_mem       (parser_parser_key_s_12_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_13_from_mem       (parser_parser_key_s_13_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_14_from_mem       (parser_parser_key_s_14_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_15_from_mem       (parser_parser_key_s_15_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_16_from_mem       (parser_parser_key_s_16_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_17_from_mem       (parser_parser_key_s_17_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_18_from_mem       (parser_parser_key_s_18_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_19_from_mem       (parser_parser_key_s_19_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_1_from_mem        (parser_parser_key_s_1_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_20_from_mem       (parser_parser_key_s_20_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_21_from_mem       (parser_parser_key_s_21_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_22_from_mem       (parser_parser_key_s_22_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_23_from_mem       (parser_parser_key_s_23_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_24_from_mem       (parser_parser_key_s_24_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_25_from_mem       (parser_parser_key_s_25_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_26_from_mem       (parser_parser_key_s_26_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_27_from_mem       (parser_parser_key_s_27_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_28_from_mem       (parser_parser_key_s_28_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_29_from_mem       (parser_parser_key_s_29_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_2_from_mem        (parser_parser_key_s_2_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_30_from_mem       (parser_parser_key_s_30_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_31_from_mem       (parser_parser_key_s_31_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_key_s_3_from_mem        (parser_parser_key_s_3_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_4_from_mem        (parser_parser_key_s_4_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_5_from_mem        (parser_parser_key_s_5_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_6_from_mem        (parser_parser_key_s_6_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_7_from_mem        (parser_parser_key_s_7_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_8_from_mem        (parser_parser_key_s_8_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_key_s_9_from_mem        (parser_parser_key_s_9_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_0_from_mem        (parser_parser_key_w_0_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_10_from_mem       (parser_parser_key_w_10_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_11_from_mem       (parser_parser_key_w_11_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_12_from_mem       (parser_parser_key_w_12_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_13_from_mem       (parser_parser_key_w_13_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_14_from_mem       (parser_parser_key_w_14_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_15_from_mem       (parser_parser_key_w_15_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_16_from_mem       (parser_parser_key_w_16_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_17_from_mem       (parser_parser_key_w_17_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_18_from_mem       (parser_parser_key_w_18_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_19_from_mem       (parser_parser_key_w_19_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_1_from_mem        (parser_parser_key_w_1_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_20_from_mem       (parser_parser_key_w_20_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_21_from_mem       (parser_parser_key_w_21_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_22_from_mem       (parser_parser_key_w_22_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_23_from_mem       (parser_parser_key_w_23_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_24_from_mem       (parser_parser_key_w_24_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_25_from_mem       (parser_parser_key_w_25_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_26_from_mem       (parser_parser_key_w_26_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_27_from_mem       (parser_parser_key_w_27_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_28_from_mem       (parser_parser_key_w_28_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_29_from_mem       (parser_parser_key_w_29_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_2_from_mem        (parser_parser_key_w_2_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_30_from_mem       (parser_parser_key_w_30_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_31_from_mem       (parser_parser_key_w_31_from_mem),                 
/* input  logic   [72:0] */ .parser_parser_key_w_3_from_mem        (parser_parser_key_w_3_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_4_from_mem        (parser_parser_key_w_4_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_5_from_mem        (parser_parser_key_w_5_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_6_from_mem        (parser_parser_key_w_6_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_7_from_mem        (parser_parser_key_w_7_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_8_from_mem        (parser_parser_key_w_8_from_mem),                  
/* input  logic   [72:0] */ .parser_parser_key_w_9_from_mem        (parser_parser_key_w_9_from_mem),                  
/* input  logic   [69:0] */ .parser_parser_metadata_fifo_from_mem  (parser_parser_metadata_fifo_from_mem),            
/* input  logic   [72:0] */ .parser_parser_port_cfg_0_from_mem     (parser_parser_port_cfg_0_from_mem),               
/* input  logic   [72:0] */ .parser_parser_port_cfg_1_from_mem     (parser_parser_port_cfg_1_from_mem),               
/* input  logic   [20:0] */ .parser_parser_ptype_ram_from_mem      (parser_parser_ptype_ram_from_mem),                
/* input  logic          */ .parser_port_cfg_0_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_port_cfg_0_rd_adr              (),                                                
/* input  logic          */ .parser_port_cfg_0_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_port_cfg_0_wr_adr              (),                                                
/* input  logic   [63:0] */ .parser_port_cfg_0_wr_data             (),                                                
/* input  logic          */ .parser_port_cfg_0_wr_en               (),                                                
/* input  logic          */ .parser_port_cfg_1_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_port_cfg_1_rd_adr              (),                                                
/* input  logic          */ .parser_port_cfg_1_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_port_cfg_1_wr_adr              (),                                                
/* input  logic   [63:0] */ .parser_port_cfg_1_wr_data             (),                                                
/* input  logic          */ .parser_port_cfg_1_wr_en               (),                                                
/* input  logic    [5:0] */ .parser_ptype_ram_adr                  (),                                                
/* input  logic          */ .parser_ptype_ram_mem_ls_enter         (),                                                
/* input  logic          */ .parser_ptype_ram_rd_en                (),                                                
/* input  logic   [13:0] */ .parser_ptype_ram_wr_data              (),                                                
/* input  logic          */ .parser_ptype_ram_wr_en                (),                                                
/* input  logic          */ .reset_n                               (reset_n),                                         
/* input  logic          */ .unified_regs_rd                       (),                                                
/* input  logic   [31:0] */ .unified_regs_wr_data                  (),                                                
/* input  logic          */ .parser_key_w_18_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_19_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_19_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_19_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_19_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_19_wr_data               (),                                                
/* input  logic          */ .parser_key_w_19_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_1_mem_ls_enter           (),                                                
/* input  logic    [3:0] */ .parser_key_w_1_rd_adr                 (),                                                
/* input  logic          */ .parser_key_w_1_rd_en                  (),                                                
/* input  logic    [3:0] */ .parser_key_w_1_wr_adr                 (),                                                
/* input  logic          */ .PARSER_ANA_CAM_0_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_0_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_10_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_10_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_11_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_11_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_12_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_12_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_S_3_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_S_4_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_ANA_S_4_STATUS_reg_sel         (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_18_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_18_rd_en               (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_18_wr_adr              (),                                                
/* input  logic   [25:0] */ .parser_ana_ext_18_wr_data             (),                                                
/* input  logic          */ .parser_ana_ext_30_wr_en               (),                                                
/* input  logic          */ .parser_ana_ext_31_mem_ls_enter        (),                                                
/* input  logic    [4:0] */ .parser_ana_ext_31_rd_adr              (),                                                
/* input  logic          */ .parser_ana_ext_31_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_10_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_10_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_10_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_11_mem_ls_enter        (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_23_wr_adr              (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_23_wr_data             (),                                                
/* input  logic          */ .parser_ana_cam_23_wr_en               (),                                                
/* input  logic          */ .parser_ana_cam_24_mem_ls_enter        (),                                                
/* input  logic          */ .parser_ana_cam_8_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_cam_8_wr_adr               (),                                                
/* input  logic   [95:0] */ .parser_ana_cam_8_wr_data              (),                                                
/* input  logic          */ .parser_key_s_19_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_19_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_19_wr_data               (),                                                
/* input  logic          */ .parser_key_s_19_wr_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_s_31_wr_adr                (),                                                
/* input  logic   [31:0] */ .parser_key_s_31_wr_data               (),                                                
/* input  logic          */ .parser_key_s_31_wr_en                 (),                                                
/* input  logic          */ .parser_key_s_3_mem_ls_enter           (),                                                
/* input  logic  [104:0] */ .parser_parser_ana_cam_2_from_mem      (parser_parser_ana_cam_2_from_mem),                
/* input  logic  [104:0] */ .parser_parser_ana_cam_30_from_mem     (parser_parser_ana_cam_30_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_31_from_mem     (parser_parser_ana_cam_31_from_mem),               
/* input  logic  [104:0] */ .parser_parser_ana_cam_3_from_mem      (parser_parser_ana_cam_3_from_mem),                
/* input  logic          */ .parser_ana_exc_20_rd_en               (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_20_wr_adr              (),                                                
/* input  logic    [8:0] */ .parser_ana_exc_20_wr_data             (),                                                
/* input  logic          */ .parser_ana_exc_20_wr_en               (),                                                
/* input  logic          */ .parser_ana_exc_5_mem_ls_enter         (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_5_rd_adr               (),                                                
/* input  logic          */ .parser_ana_exc_5_rd_en                (),                                                
/* input  logic    [3:0] */ .parser_ana_exc_5_wr_adr               (),                                                
/* input  logic          */ .PARSER_KEY_S_6_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_7_CFG_reg_sel            (),                                                
/* input  logic          */ .PARSER_KEY_S_7_STATUS_reg_sel         (),                                                
/* input  logic          */ .PARSER_KEY_S_8_CFG_reg_sel            (),                                                
/* input  logic          */ .parser_ana_s_15_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_15_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_15_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_15_wr_adr                (),                                                
/* input  logic          */ .parser_ana_s_28_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_s_28_rd_adr                (),                                                
/* input  logic          */ .parser_ana_s_28_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_ana_s_28_wr_adr                (),                                                
/* input  logic          */ .PARSER_ANA_EXC_14_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_14_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_15_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_23_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_23_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_24_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_24_STATUS_reg_sel      (),                                                
/* input  logic          */ .parser_ana_w_11_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_12_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_12_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_12_rd_en                 (),                                                
/* input  logic          */ .parser_ana_w_24_wr_en                 (),                                                
/* input  logic          */ .parser_ana_w_25_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_ana_w_25_rd_adr                (),                                                
/* input  logic          */ .parser_ana_w_25_rd_en                 (),                                                
/* input  logic   [39:0] */ .parser_parser_ana_w_31_from_mem       (parser_parser_ana_w_31_from_mem),                 
/* input  logic   [39:0] */ .parser_parser_ana_w_3_from_mem        (parser_parser_ana_w_3_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_4_from_mem        (parser_parser_ana_w_4_from_mem),                  
/* input  logic   [39:0] */ .parser_parser_ana_w_5_from_mem        (parser_parser_ana_w_5_from_mem),                  
/* input  logic    [3:0] */ .parser_key_w_15_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_15_wr_data               (),                                                
/* input  logic          */ .parser_key_w_15_wr_en                 (),                                                
/* input  logic          */ .parser_key_w_16_mem_ls_enter          (),                                                
/* input  logic    [3:0] */ .parser_key_w_16_rd_adr                (),                                                
/* input  logic          */ .parser_key_w_16_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_16_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_16_wr_data               (),                                                
/* input  logic          */ .parser_key_w_29_rd_en                 (),                                                
/* input  logic    [3:0] */ .parser_key_w_29_wr_adr                (),                                                
/* input  logic   [63:0] */ .parser_key_w_29_wr_data               (),                                                
/* input  logic          */ .parser_key_w_29_wr_en                 (),                                                
/* input  logic   [31:0] */ .parser_ana_w_9_wr_data                (),                                                
/* input  logic          */ .parser_ana_w_9_wr_en                  (),                                                
/* input  logic          */ .parser_csum_cfg_0_mem_ls_enter        (),                                                
/* input  logic   [79:0] */ .parser_extract_cfg_5_wr_data          (),                                                
/* input  logic          */ .parser_extract_cfg_5_wr_en            (),                                                
/* input  logic          */ .parser_extract_cfg_6_mem_ls_enter     (),                                                
/* input  logic    [3:0] */ .parser_extract_cfg_6_rd_adr           (),                                                
/* input  logic          */ .PARSER_ANA_CAM_13_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_13_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_14_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_14_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_15_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_15_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_16_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_16_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_17_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_17_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_18_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_18_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_19_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_19_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_1_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_1_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_20_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_20_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_21_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_21_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_22_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_22_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_23_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_23_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_24_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_24_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_25_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_25_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_26_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_26_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_27_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_27_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_28_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_28_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_29_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_29_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_2_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_2_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_30_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_30_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_31_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_CAM_31_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_CAM_3_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_3_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_4_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_4_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_5_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_5_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_6_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_6_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_7_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_7_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_8_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_8_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_CAM_9_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_CAM_9_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_0_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_0_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_10_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_10_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_11_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_11_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_12_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_12_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_13_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_13_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_15_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_16_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_16_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_17_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_17_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_18_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_18_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_19_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_19_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_1_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_1_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_20_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_20_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_21_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_21_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_22_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_22_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_23_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_23_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_24_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_24_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_25_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_25_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_26_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_26_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_27_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_27_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_28_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_28_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_29_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_29_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_2_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_2_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_30_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_30_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_31_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXC_31_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXC_3_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_3_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_4_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_4_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_5_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_5_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_6_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_6_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_7_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_7_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_8_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_8_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXC_9_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXC_9_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_0_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_0_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_10_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_10_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_11_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_11_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_12_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_12_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_13_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_13_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_14_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_14_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_15_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_15_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_16_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_16_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_17_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_17_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_18_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_18_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_19_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_19_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_1_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_1_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_20_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_20_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_21_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_21_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_22_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_22_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_25_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_25_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_26_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_26_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_27_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_27_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_28_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_28_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_29_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_29_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_2_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_2_STATUS_reg_sel       (),                                                
/* input  logic          */ .PARSER_ANA_EXT_30_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_30_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_31_CFG_reg_sel         (),                                                
/* input  logic          */ .PARSER_ANA_EXT_31_STATUS_reg_sel      (),                                                
/* input  logic          */ .PARSER_ANA_EXT_3_CFG_reg_sel          (),                                                
/* input  logic          */ .PARSER_ANA_EXT_3_STATUS_reg_sel       (),                                                
/* output logic          */ .parser_ana_cam_0_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_0_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_0_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_0_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_10_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_10_init_done           (),                                                
/* output logic          */ .parser_ana_cam_11_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_11_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_11_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_12_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_12_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_12_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_12_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_13_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_13_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_13_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_13_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_14_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_14_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_14_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_14_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_15_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_15_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_15_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_15_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_16_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_16_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_16_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_16_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_17_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_17_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_17_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_17_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_18_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_18_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_18_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_18_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_19_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_19_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_19_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_19_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_1_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_1_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_1_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_1_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_20_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_20_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_20_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_20_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_21_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_21_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_21_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_21_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_22_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_22_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_22_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_22_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_23_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_23_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_23_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_23_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_24_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_24_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_24_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_24_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_25_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_25_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_25_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_25_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_26_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_26_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_26_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_26_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_27_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_27_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_27_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_27_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_28_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_28_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_28_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_28_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_29_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_29_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_29_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_29_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_2_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_2_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_30_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_30_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_31_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_31_init_done           (),                                                
/* output logic   [95:0] */ .parser_ana_cam_31_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_31_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_3_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_3_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_3_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_3_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_4_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_4_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_4_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_4_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_5_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_5_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_5_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_5_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_6_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_6_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_6_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_6_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_7_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_7_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_7_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_7_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_8_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_8_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_8_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_8_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_9_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_cam_9_init_done            (),                                                
/* output logic   [95:0] */ .parser_ana_cam_9_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_9_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_0_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_0_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_0_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_0_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_10_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_10_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_10_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_10_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_11_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_11_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_11_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_11_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_12_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_12_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_12_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_12_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_13_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_13_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_13_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_13_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_14_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_14_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_14_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_14_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_15_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_15_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_15_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_15_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_16_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_16_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_16_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_16_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_17_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_17_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_17_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_17_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_18_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_18_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_18_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_18_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_19_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_19_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_19_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_19_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_1_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_1_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_1_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_1_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_20_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_20_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_21_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_21_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_22_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_22_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_22_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_22_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_23_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_23_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_23_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_23_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_24_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_24_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_24_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_24_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_25_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_25_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_25_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_25_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_26_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_26_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_26_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_26_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_27_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_27_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_27_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_27_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_28_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_28_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_28_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_28_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_29_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_29_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_29_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_29_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_2_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_2_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_2_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_2_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_30_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_30_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_30_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_30_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_31_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_31_init_done           (),                                                
/* output logic    [8:0] */ .parser_ana_exc_31_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_31_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_3_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_3_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_3_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_3_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_4_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_4_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_4_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_4_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_5_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_5_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_5_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_5_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_6_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_6_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_6_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_6_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_7_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_7_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_7_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_7_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_8_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_8_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_8_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_8_rd_valid             (),                                                
/* output logic          */ .parser_ana_exc_9_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_exc_9_init_done            (),                                                
/* output logic    [8:0] */ .parser_ana_exc_9_rd_data              (),                                                
/* output logic          */ .parser_ana_exc_9_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_0_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_0_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_0_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_0_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_10_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_10_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_10_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_11_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_12_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_12_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_12_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_12_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_13_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_13_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_13_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_13_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_14_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_14_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_14_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_14_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_15_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_15_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_15_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_15_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_16_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_16_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_16_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_16_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_17_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_17_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_17_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_17_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_18_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_18_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_18_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_18_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_19_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_19_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_19_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_19_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_1_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_1_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_1_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_1_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_20_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_20_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_20_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_20_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_21_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_21_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_21_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_21_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_22_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_22_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_22_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_22_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_23_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_23_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_23_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_23_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_24_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_24_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_24_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_24_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_25_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_25_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_25_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_25_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_26_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_26_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_26_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_26_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_27_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_27_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_27_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_27_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_28_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_28_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_28_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_28_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_29_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_29_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_29_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_29_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_2_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_2_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_2_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_30_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_31_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_31_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_31_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_31_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_3_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_3_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_3_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_3_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_4_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_4_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_4_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_4_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_5_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_5_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_5_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_5_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_6_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_6_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_6_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_6_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_7_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_7_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_7_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_7_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_8_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_8_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_8_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_8_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_9_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ana_ext_9_init_done            (),                                                
/* output logic   [25:0] */ .parser_ana_ext_9_rd_data              (),                                                
/* output logic          */ .parser_ana_ext_9_rd_valid             (),                                                
/* output logic          */ .parser_ana_s_0_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_0_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_0_rd_data                (),                                                
/* output logic          */ .parser_ana_s_0_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_10_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_10_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_10_rd_data               (),                                                
/* output logic          */ .parser_ana_s_10_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_11_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_11_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_11_rd_data               (),                                                
/* output logic          */ .parser_ana_s_11_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_12_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_12_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_12_rd_data               (),                                                
/* output logic          */ .parser_ana_s_12_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_13_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_13_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_13_rd_data               (),                                                
/* output logic          */ .parser_ana_s_13_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_14_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_14_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_14_rd_data               (),                                                
/* output logic          */ .parser_ana_s_14_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_15_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_15_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_15_rd_data               (),                                                
/* output logic          */ .parser_ana_s_15_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_16_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_16_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_16_rd_data               (),                                                
/* output logic          */ .parser_ana_s_16_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_17_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_17_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_17_rd_data               (),                                                
/* output logic          */ .parser_ana_s_17_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_18_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_18_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_18_rd_data               (),                                                
/* output logic          */ .parser_ana_s_18_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_19_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_19_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_19_rd_data               (),                                                
/* output logic          */ .parser_ana_s_19_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_1_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_1_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_1_rd_data                (),                                                
/* output logic          */ .parser_ana_s_1_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_20_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_20_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_20_rd_data               (),                                                
/* output logic          */ .parser_ana_s_20_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_21_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_21_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_21_rd_data               (),                                                
/* output logic          */ .parser_ana_s_21_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_22_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_22_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_22_rd_data               (),                                                
/* output logic          */ .parser_ana_s_22_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_23_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_23_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_23_rd_data               (),                                                
/* output logic          */ .parser_ana_s_23_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_24_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_24_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_24_rd_data               (),                                                
/* output logic          */ .parser_ana_s_24_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_25_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_25_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_25_rd_data               (),                                                
/* output logic          */ .parser_ana_s_25_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_26_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_26_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_26_rd_data               (),                                                
/* output logic          */ .parser_ana_s_26_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_27_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_27_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_27_rd_data               (),                                                
/* output logic          */ .parser_ana_s_27_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_28_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_28_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_28_rd_data               (),                                                
/* output logic          */ .parser_ana_s_28_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_29_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_29_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_29_rd_data               (),                                                
/* output logic          */ .parser_ana_s_29_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_2_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_2_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_2_rd_data                (),                                                
/* output logic          */ .parser_ana_s_2_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_30_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_30_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_30_rd_data               (),                                                
/* output logic          */ .parser_ana_s_30_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_31_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_s_31_init_done             (),                                                
/* output logic   [47:0] */ .parser_ana_s_31_rd_data               (),                                                
/* output logic          */ .parser_ana_s_31_rd_valid              (),                                                
/* output logic          */ .parser_ana_s_3_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_3_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_3_rd_data                (),                                                
/* output logic          */ .parser_ana_s_3_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_4_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_4_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_4_rd_data                (),                                                
/* output logic          */ .parser_ana_s_4_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_5_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_5_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_5_rd_data                (),                                                
/* output logic          */ .parser_ana_s_5_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_6_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_6_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_6_rd_data                (),                                                
/* output logic          */ .parser_ana_s_6_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_7_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_7_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_7_rd_data                (),                                                
/* output logic          */ .parser_ana_s_7_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_8_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_8_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_8_rd_data                (),                                                
/* output logic          */ .parser_ana_s_8_rd_valid               (),                                                
/* output logic          */ .parser_ana_s_9_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_s_9_init_done              (),                                                
/* output logic   [47:0] */ .parser_ana_s_9_rd_data                (),                                                
/* output logic          */ .parser_ana_s_9_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_0_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_0_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_0_rd_data                (),                                                
/* output logic          */ .parser_ana_w_0_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_10_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_10_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_10_rd_data               (),                                                
/* output logic          */ .parser_ana_w_10_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_12_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_12_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_12_rd_data               (),                                                
/* output logic          */ .parser_ana_w_12_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_13_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_13_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_13_rd_data               (),                                                
/* output logic          */ .parser_ana_w_13_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_14_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_14_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_14_rd_data               (),                                                
/* output logic          */ .parser_ana_w_14_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_15_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_15_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_15_rd_data               (),                                                
/* output logic          */ .parser_ana_w_15_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_16_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_16_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_16_rd_data               (),                                                
/* output logic          */ .parser_ana_w_16_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_17_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_17_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_17_rd_data               (),                                                
/* output logic          */ .parser_ana_w_17_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_18_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_18_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_18_rd_data               (),                                                
/* output logic          */ .parser_ana_w_18_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_19_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_19_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_19_rd_data               (),                                                
/* output logic          */ .parser_ana_w_19_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_1_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_1_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_1_rd_data                (),                                                
/* output logic          */ .parser_ana_w_1_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_20_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_20_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_20_rd_data               (),                                                
/* output logic          */ .parser_ana_w_20_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_21_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_21_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_21_rd_data               (),                                                
/* output logic          */ .parser_ana_w_21_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_22_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_22_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_22_rd_data               (),                                                
/* output logic          */ .parser_ana_w_22_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_23_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_23_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_23_rd_data               (),                                                
/* output logic          */ .parser_ana_w_23_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_24_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_24_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_24_rd_data               (),                                                
/* output logic          */ .parser_ana_w_24_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_25_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_25_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_25_rd_data               (),                                                
/* output logic          */ .parser_ana_w_25_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_26_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_26_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_26_rd_data               (),                                                
/* output logic          */ .parser_ana_w_26_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_27_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_27_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_27_rd_data               (),                                                
/* output logic          */ .parser_ana_w_27_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_28_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_28_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_28_rd_data               (),                                                
/* output logic          */ .parser_ana_w_28_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_29_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_29_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_29_rd_data               (),                                                
/* output logic          */ .parser_ana_w_29_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_2_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_2_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_2_rd_data                (),                                                
/* output logic          */ .parser_ana_w_2_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_30_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_30_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_30_rd_data               (),                                                
/* output logic          */ .parser_ana_w_30_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_31_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_3_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_3_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_3_rd_data                (),                                                
/* output logic          */ .parser_ana_w_3_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_4_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_4_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_4_rd_data                (),                                                
/* output logic          */ .parser_ana_w_4_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_5_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_5_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_5_rd_data                (),                                                
/* output logic          */ .parser_ana_w_5_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_6_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_6_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_6_rd_data                (),                                                
/* output logic          */ .parser_ana_w_6_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_7_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_7_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_7_rd_data                (),                                                
/* output logic          */ .parser_ana_w_7_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_8_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_8_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_8_rd_data                (),                                                
/* output logic          */ .parser_ana_w_8_rd_valid               (),                                                
/* output logic          */ .parser_ana_w_9_ecc_uncor_err          (),                                                
/* output logic          */ .parser_ana_w_9_init_done              (),                                                
/* output logic   [31:0] */ .parser_ana_w_9_rd_data                (),                                                
/* output logic          */ .parser_ana_w_9_rd_valid               (),                                                
/* output logic          */ .parser_csum_cfg_0_ecc_uncor_err       (),                                                
/* output logic          */ .parser_csum_cfg_0_init_done           (),                                                
/* output logic    [5:0] */ .parser_csum_cfg_0_rd_data             (),                                                
/* output logic          */ .parser_csum_cfg_0_rd_valid            (),                                                
/* output logic          */ .parser_csum_cfg_1_ecc_uncor_err       (),                                                
/* output logic          */ .parser_csum_cfg_1_init_done           (),                                                
/* output logic    [5:0] */ .parser_csum_cfg_1_rd_data             (),                                                
/* output logic          */ .parser_csum_cfg_1_rd_valid            (),                                                
/* output logic          */ .parser_ecc_int                        (),                                                
/* output logic          */ .parser_extract_cfg_0_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_0_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_0_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_0_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_10_ecc_uncor_err   (),                                                
/* output logic          */ .parser_extract_cfg_10_init_done       (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_10_rd_data         (),                                                
/* output logic          */ .parser_extract_cfg_10_rd_valid        (),                                                
/* output logic          */ .parser_extract_cfg_11_ecc_uncor_err   (),                                                
/* output logic          */ .parser_extract_cfg_11_init_done       (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_11_rd_data         (),                                                
/* output logic          */ .parser_extract_cfg_11_rd_valid        (),                                                
/* output logic          */ .parser_extract_cfg_12_ecc_uncor_err   (),                                                
/* output logic          */ .parser_extract_cfg_12_init_done       (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_12_rd_data         (),                                                
/* output logic          */ .parser_extract_cfg_12_rd_valid        (),                                                
/* output logic          */ .parser_extract_cfg_13_ecc_uncor_err   (),                                                
/* output logic          */ .parser_extract_cfg_13_init_done       (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_13_rd_data         (),                                                
/* output logic          */ .parser_extract_cfg_13_rd_valid        (),                                                
/* output logic          */ .parser_extract_cfg_14_ecc_uncor_err   (),                                                
/* output logic          */ .parser_extract_cfg_14_init_done       (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_14_rd_data         (),                                                
/* output logic          */ .parser_extract_cfg_14_rd_valid        (),                                                
/* output logic          */ .parser_extract_cfg_15_ecc_uncor_err   (),                                                
/* output logic          */ .parser_extract_cfg_15_init_done       (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_15_rd_data         (),                                                
/* output logic          */ .parser_extract_cfg_15_rd_valid        (),                                                
/* output logic          */ .parser_extract_cfg_1_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_1_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_1_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_1_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_2_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_2_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_2_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_2_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_3_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_3_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_3_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_3_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_4_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_4_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_4_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_4_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_6_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_6_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_6_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_6_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_7_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_7_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_7_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_7_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_8_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_8_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_8_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_8_rd_valid         (),                                                
/* output logic          */ .parser_extract_cfg_9_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_9_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_9_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_9_rd_valid         (),                                                
/* output logic          */ .parser_init_done                      (),                                                
/* output logic          */ .parser_key_s_0_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_0_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_0_rd_data                (),                                                
/* output logic          */ .parser_key_s_0_rd_valid               (),                                                
/* output logic          */ .parser_key_s_10_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_10_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_10_rd_data               (),                                                
/* output logic          */ .parser_key_s_10_rd_valid              (),                                                
/* output logic          */ .parser_key_s_11_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_11_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_11_rd_data               (),                                                
/* output logic          */ .parser_key_s_11_rd_valid              (),                                                
/* output logic          */ .parser_key_s_12_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_12_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_12_rd_data               (),                                                
/* output logic          */ .parser_key_s_12_rd_valid              (),                                                
/* output logic          */ .parser_key_s_13_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_13_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_13_rd_data               (),                                                
/* output logic          */ .parser_key_s_13_rd_valid              (),                                                
/* output logic          */ .parser_key_s_14_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_14_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_14_rd_data               (),                                                
/* output logic          */ .parser_key_s_14_rd_valid              (),                                                
/* output logic          */ .parser_key_s_15_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_15_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_15_rd_data               (),                                                
/* output logic          */ .parser_key_s_15_rd_valid              (),                                                
/* output logic          */ .parser_key_s_16_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_16_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_16_rd_data               (),                                                
/* output logic          */ .parser_key_s_16_rd_valid              (),                                                
/* output logic          */ .parser_key_s_17_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_17_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_17_rd_data               (),                                                
/* output logic          */ .parser_key_s_17_rd_valid              (),                                                
/* output logic          */ .parser_key_s_18_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_18_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_18_rd_data               (),                                                
/* output logic          */ .parser_key_s_18_rd_valid              (),                                                
/* output logic          */ .parser_key_s_19_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_19_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_19_rd_data               (),                                                
/* output logic          */ .parser_key_s_19_rd_valid              (),                                                
/* output logic          */ .parser_key_s_1_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_1_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_1_rd_data                (),                                                
/* output logic          */ .parser_key_s_1_rd_valid               (),                                                
/* output logic          */ .parser_key_s_20_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_20_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_20_rd_data               (),                                                
/* output logic          */ .parser_key_s_20_rd_valid              (),                                                
/* output logic          */ .parser_key_s_21_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_21_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_21_rd_data               (),                                                
/* output logic          */ .parser_key_s_21_rd_valid              (),                                                
/* output logic          */ .parser_key_s_22_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_22_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_22_rd_data               (),                                                
/* output logic          */ .parser_key_s_22_rd_valid              (),                                                
/* output logic          */ .parser_key_s_23_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_23_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_23_rd_data               (),                                                
/* output logic          */ .parser_key_s_23_rd_valid              (),                                                
/* output logic          */ .parser_key_s_24_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_24_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_24_rd_data               (),                                                
/* output logic          */ .parser_key_s_25_rd_valid              (),                                                
/* output logic          */ .parser_key_s_26_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_26_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_26_rd_data               (),                                                
/* output logic          */ .parser_key_s_26_rd_valid              (),                                                
/* output logic          */ .parser_key_s_27_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_27_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_27_rd_data               (),                                                
/* output logic          */ .parser_key_s_27_rd_valid              (),                                                
/* output logic          */ .parser_key_s_28_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_28_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_28_rd_data               (),                                                
/* output logic          */ .parser_key_s_28_rd_valid              (),                                                
/* output logic          */ .parser_key_s_29_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_29_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_29_rd_data               (),                                                
/* output logic          */ .parser_key_s_29_rd_valid              (),                                                
/* output logic          */ .parser_key_s_2_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_2_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_2_rd_data                (),                                                
/* output logic          */ .parser_key_s_2_rd_valid               (),                                                
/* output logic          */ .parser_key_s_30_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_30_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_30_rd_data               (),                                                
/* output logic          */ .parser_key_s_30_rd_valid              (),                                                
/* output logic          */ .parser_key_s_31_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_31_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_31_rd_data               (),                                                
/* output logic          */ .parser_key_s_31_rd_valid              (),                                                
/* output logic          */ .parser_key_s_3_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_3_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_3_rd_data                (),                                                
/* output logic          */ .parser_key_s_3_rd_valid               (),                                                
/* output logic          */ .parser_key_s_4_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_4_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_4_rd_data                (),                                                
/* output logic          */ .parser_key_s_4_rd_valid               (),                                                
/* output logic          */ .parser_key_s_5_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_5_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_5_rd_data                (),                                                
/* output logic          */ .parser_key_s_5_rd_valid               (),                                                
/* output logic          */ .parser_key_s_6_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_6_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_6_rd_data                (),                                                
/* output logic          */ .parser_key_s_6_rd_valid               (),                                                
/* output logic          */ .parser_key_s_7_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_7_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_7_rd_data                (),                                                
/* output logic          */ .parser_key_s_7_rd_valid               (),                                                
/* output logic          */ .parser_key_s_8_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_8_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_8_rd_data                (),                                                
/* output logic          */ .parser_key_s_8_rd_valid               (),                                                
/* output logic          */ .parser_key_s_9_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_s_9_init_done              (),                                                
/* output logic   [31:0] */ .parser_key_s_9_rd_data                (),                                                
/* output logic          */ .parser_key_s_9_rd_valid               (),                                                
/* output logic          */ .parser_key_w_0_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_0_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_0_rd_data                (),                                                
/* output logic          */ .parser_key_w_0_rd_valid               (),                                                
/* output logic          */ .parser_key_w_10_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_10_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_10_rd_data               (),                                                
/* output logic          */ .parser_key_w_10_rd_valid              (),                                                
/* output logic          */ .parser_key_w_11_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_11_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_11_rd_data               (),                                                
/* output logic          */ .parser_key_w_11_rd_valid              (),                                                
/* output logic          */ .parser_key_w_12_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_12_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_12_rd_data               (),                                                
/* output logic          */ .parser_key_w_12_rd_valid              (),                                                
/* output logic          */ .parser_key_w_13_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_13_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_13_rd_data               (),                                                
/* output logic          */ .parser_key_w_13_rd_valid              (),                                                
/* output logic          */ .parser_key_w_14_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_14_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_14_rd_data               (),                                                
/* output logic          */ .parser_key_w_14_rd_valid              (),                                                
/* output logic          */ .parser_key_w_16_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_16_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_16_rd_data               (),                                                
/* output logic          */ .parser_key_w_16_rd_valid              (),                                                
/* output logic          */ .parser_key_w_17_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_17_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_17_rd_data               (),                                                
/* output logic          */ .parser_key_w_17_rd_valid              (),                                                
/* output logic          */ .parser_key_w_18_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_18_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_18_rd_data               (),                                                
/* output logic          */ .parser_key_w_18_rd_valid              (),                                                
/* output logic          */ .parser_key_w_19_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_19_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_19_rd_data               (),                                                
/* output logic          */ .parser_key_w_19_rd_valid              (),                                                
/* output logic          */ .parser_key_w_1_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_1_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_1_rd_data                (),                                                
/* output logic          */ .parser_key_w_1_rd_valid               (),                                                
/* output logic          */ .parser_key_w_20_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_20_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_20_rd_data               (),                                                
/* output logic          */ .parser_key_w_20_rd_valid              (),                                                
/* output logic          */ .parser_key_w_21_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_21_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_21_rd_data               (),                                                
/* output logic          */ .parser_key_w_21_rd_valid              (),                                                
/* output logic          */ .parser_key_w_22_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_22_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_22_rd_data               (),                                                
/* output logic          */ .parser_key_w_22_rd_valid              (),                                                
/* output logic          */ .parser_key_w_23_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_23_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_23_rd_data               (),                                                
/* output logic          */ .parser_key_w_23_rd_valid              (),                                                
/* output logic          */ .parser_key_w_24_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_24_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_24_rd_data               (),                                                
/* output logic          */ .parser_key_w_24_rd_valid              (),                                                
/* output logic          */ .parser_key_w_25_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_25_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_25_rd_data               (),                                                
/* output logic          */ .parser_key_w_25_rd_valid              (),                                                
/* output logic          */ .parser_key_w_26_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_26_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_26_rd_data               (),                                                
/* output logic          */ .parser_key_w_26_rd_valid              (),                                                
/* output logic          */ .parser_key_w_27_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_27_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_27_rd_data               (),                                                
/* output logic          */ .parser_key_w_27_rd_valid              (),                                                
/* output logic          */ .parser_key_w_28_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_28_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_28_rd_data               (),                                                
/* output logic          */ .parser_key_w_28_rd_valid              (),                                                
/* output logic          */ .parser_key_w_29_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_29_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_29_rd_data               (),                                                
/* output logic          */ .parser_key_w_29_rd_valid              (),                                                
/* output logic          */ .parser_key_w_2_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_2_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_2_rd_data                (),                                                
/* output logic          */ .parser_key_w_2_rd_valid               (),                                                
/* output logic          */ .parser_key_w_30_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_30_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_30_rd_data               (),                                                
/* output logic          */ .parser_key_w_30_rd_valid              (),                                                
/* output logic          */ .parser_key_w_31_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_31_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_31_rd_data               (),                                                
/* output logic          */ .parser_key_w_31_rd_valid              (),                                                
/* output logic          */ .parser_key_w_3_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_3_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_3_rd_data                (),                                                
/* output logic          */ .parser_key_w_3_rd_valid               (),                                                
/* output logic          */ .parser_key_w_4_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_4_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_4_rd_data                (),                                                
/* output logic          */ .parser_key_w_4_rd_valid               (),                                                
/* output logic          */ .parser_key_w_5_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_5_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_5_rd_data                (),                                                
/* output logic          */ .parser_key_w_5_rd_valid               (),                                                
/* output logic          */ .parser_key_w_7_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_7_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_7_rd_data                (),                                                
/* output logic          */ .parser_key_w_7_rd_valid               (),                                                
/* output logic          */ .parser_key_w_8_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_8_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_8_rd_data                (),                                                
/* output logic          */ .parser_key_w_8_rd_valid               (),                                                
/* output logic          */ .parser_key_w_9_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_9_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_9_rd_data                (),                                                
/* output logic          */ .parser_key_w_9_rd_valid               (),                                                
/* output logic          */ .parser_metadata_fifo_ecc_uncor_err    (),                                                
/* output logic          */ .parser_metadata_fifo_init_done        (),                                                
/* output logic   [60:0] */ .parser_metadata_fifo_rd_data          (),                                                
/* output logic          */ .parser_metadata_fifo_rd_valid         (),                                                
/* output logic  [119:0] */ .parser_parser_ana_cam_0_to_mem        (parser_parser_ana_cam_0_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_10_to_mem       (parser_parser_ana_cam_10_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_11_to_mem       (parser_parser_ana_cam_11_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_12_to_mem       (parser_parser_ana_cam_12_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_13_to_mem       (parser_parser_ana_cam_13_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_14_to_mem       (parser_parser_ana_cam_14_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_15_to_mem       (parser_parser_ana_cam_15_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_16_to_mem       (parser_parser_ana_cam_16_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_17_to_mem       (parser_parser_ana_cam_17_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_18_to_mem       (parser_parser_ana_cam_18_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_19_to_mem       (parser_parser_ana_cam_19_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_1_to_mem        (parser_parser_ana_cam_1_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_20_to_mem       (parser_parser_ana_cam_20_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_21_to_mem       (parser_parser_ana_cam_21_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_22_to_mem       (parser_parser_ana_cam_22_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_23_to_mem       (parser_parser_ana_cam_23_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_24_to_mem       (parser_parser_ana_cam_24_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_25_to_mem       (parser_parser_ana_cam_25_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_26_to_mem       (parser_parser_ana_cam_26_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_27_to_mem       (parser_parser_ana_cam_27_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_28_to_mem       (parser_parser_ana_cam_28_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_29_to_mem       (parser_parser_ana_cam_29_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_2_to_mem        (parser_parser_ana_cam_2_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_30_to_mem       (parser_parser_ana_cam_30_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_31_to_mem       (parser_parser_ana_cam_31_to_mem),                 
/* output logic  [119:0] */ .parser_parser_ana_cam_3_to_mem        (parser_parser_ana_cam_3_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_4_to_mem        (parser_parser_ana_cam_4_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_5_to_mem        (parser_parser_ana_cam_5_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_6_to_mem        (parser_parser_ana_cam_6_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_7_to_mem        (parser_parser_ana_cam_7_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_8_to_mem        (parser_parser_ana_cam_8_to_mem),                  
/* output logic  [119:0] */ .parser_parser_ana_cam_9_to_mem        (parser_parser_ana_cam_9_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_0_to_mem        (parser_parser_ana_exc_0_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_10_to_mem       (parser_parser_ana_exc_10_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_11_to_mem       (parser_parser_ana_exc_11_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_12_to_mem       (parser_parser_ana_exc_12_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_13_to_mem       (parser_parser_ana_exc_13_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_14_to_mem       (parser_parser_ana_exc_14_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_15_to_mem       (parser_parser_ana_exc_15_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_16_to_mem       (parser_parser_ana_exc_16_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_17_to_mem       (parser_parser_ana_exc_17_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_18_to_mem       (parser_parser_ana_exc_18_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_19_to_mem       (parser_parser_ana_exc_19_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_1_to_mem        (parser_parser_ana_exc_1_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_20_to_mem       (parser_parser_ana_exc_20_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_21_to_mem       (parser_parser_ana_exc_21_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_22_to_mem       (parser_parser_ana_exc_22_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_23_to_mem       (parser_parser_ana_exc_23_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_24_to_mem       (parser_parser_ana_exc_24_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_25_to_mem       (parser_parser_ana_exc_25_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_26_to_mem       (parser_parser_ana_exc_26_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_27_to_mem       (parser_parser_ana_exc_27_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_28_to_mem       (parser_parser_ana_exc_28_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_29_to_mem       (parser_parser_ana_exc_29_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_2_to_mem        (parser_parser_ana_exc_2_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_30_to_mem       (parser_parser_ana_exc_30_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_31_to_mem       (parser_parser_ana_exc_31_to_mem),                 
/* output logic   [29:0] */ .parser_parser_ana_exc_3_to_mem        (parser_parser_ana_exc_3_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_4_to_mem        (parser_parser_ana_exc_4_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_5_to_mem        (parser_parser_ana_exc_5_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_6_to_mem        (parser_parser_ana_exc_6_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_7_to_mem        (parser_parser_ana_exc_7_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_8_to_mem        (parser_parser_ana_exc_8_to_mem),                  
/* output logic   [29:0] */ .parser_parser_ana_exc_9_to_mem        (parser_parser_ana_exc_9_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_0_to_mem        (parser_parser_ana_ext_0_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_10_to_mem       (parser_parser_ana_ext_10_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_11_to_mem       (parser_parser_ana_ext_11_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_12_to_mem       (parser_parser_ana_ext_12_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_13_to_mem       (parser_parser_ana_ext_13_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_14_to_mem       (parser_parser_ana_ext_14_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_15_to_mem       (parser_parser_ana_ext_15_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_16_to_mem       (parser_parser_ana_ext_16_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_17_to_mem       (parser_parser_ana_ext_17_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_18_to_mem       (parser_parser_ana_ext_18_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_19_to_mem       (parser_parser_ana_ext_19_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_1_to_mem        (parser_parser_ana_ext_1_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_20_to_mem       (parser_parser_ana_ext_20_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_21_to_mem       (parser_parser_ana_ext_21_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_22_to_mem       (parser_parser_ana_ext_22_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_23_to_mem       (parser_parser_ana_ext_23_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_24_to_mem       (parser_parser_ana_ext_24_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_25_to_mem       (parser_parser_ana_ext_25_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_26_to_mem       (parser_parser_ana_ext_26_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_27_to_mem       (parser_parser_ana_ext_27_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_28_to_mem       (parser_parser_ana_ext_28_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_29_to_mem       (parser_parser_ana_ext_29_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_2_to_mem        (parser_parser_ana_ext_2_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_30_to_mem       (parser_parser_ana_ext_30_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_31_to_mem       (parser_parser_ana_ext_31_to_mem),                 
/* output logic   [49:0] */ .parser_parser_ana_ext_3_to_mem        (parser_parser_ana_ext_3_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_4_to_mem        (parser_parser_ana_ext_4_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_5_to_mem        (parser_parser_ana_ext_5_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_6_to_mem        (parser_parser_ana_ext_6_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_7_to_mem        (parser_parser_ana_ext_7_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_8_to_mem        (parser_parser_ana_ext_8_to_mem),                  
/* output logic   [49:0] */ .parser_parser_ana_ext_9_to_mem        (parser_parser_ana_ext_9_to_mem),                  
/* output logic   [70:0] */ .parser_parser_ana_s_0_to_mem          (parser_parser_ana_s_0_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_10_to_mem         (parser_parser_ana_s_10_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_11_to_mem         (parser_parser_ana_s_11_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_12_to_mem         (parser_parser_ana_s_12_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_13_to_mem         (parser_parser_ana_s_13_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_14_to_mem         (parser_parser_ana_s_14_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_15_to_mem         (parser_parser_ana_s_15_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_16_to_mem         (parser_parser_ana_s_16_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_17_to_mem         (parser_parser_ana_s_17_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_18_to_mem         (parser_parser_ana_s_18_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_19_to_mem         (parser_parser_ana_s_19_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_1_to_mem          (parser_parser_ana_s_1_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_20_to_mem         (parser_parser_ana_s_20_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_21_to_mem         (parser_parser_ana_s_21_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_22_to_mem         (parser_parser_ana_s_22_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_23_to_mem         (parser_parser_ana_s_23_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_24_to_mem         (parser_parser_ana_s_24_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_25_to_mem         (parser_parser_ana_s_25_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_26_to_mem         (parser_parser_ana_s_26_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_27_to_mem         (parser_parser_ana_s_27_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_28_to_mem         (parser_parser_ana_s_28_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_29_to_mem         (parser_parser_ana_s_29_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_2_to_mem          (parser_parser_ana_s_2_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_30_to_mem         (parser_parser_ana_s_30_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_31_to_mem         (parser_parser_ana_s_31_to_mem),                   
/* output logic   [70:0] */ .parser_parser_ana_s_3_to_mem          (parser_parser_ana_s_3_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_4_to_mem          (parser_parser_ana_s_4_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_5_to_mem          (parser_parser_ana_s_5_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_6_to_mem          (parser_parser_ana_s_6_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_7_to_mem          (parser_parser_ana_s_7_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_8_to_mem          (parser_parser_ana_s_8_to_mem),                    
/* output logic   [70:0] */ .parser_parser_ana_s_9_to_mem          (parser_parser_ana_s_9_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_0_to_mem          (parser_parser_ana_w_0_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_10_to_mem         (parser_parser_ana_w_10_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_11_to_mem         (parser_parser_ana_w_11_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_12_to_mem         (parser_parser_ana_w_12_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_13_to_mem         (parser_parser_ana_w_13_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_14_to_mem         (parser_parser_ana_w_14_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_15_to_mem         (parser_parser_ana_w_15_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_16_to_mem         (parser_parser_ana_w_16_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_17_to_mem         (parser_parser_ana_w_17_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_18_to_mem         (parser_parser_ana_w_18_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_19_to_mem         (parser_parser_ana_w_19_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_1_to_mem          (parser_parser_ana_w_1_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_20_to_mem         (parser_parser_ana_w_20_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_21_to_mem         (parser_parser_ana_w_21_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_22_to_mem         (parser_parser_ana_w_22_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_23_to_mem         (parser_parser_ana_w_23_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_24_to_mem         (parser_parser_ana_w_24_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_25_to_mem         (parser_parser_ana_w_25_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_26_to_mem         (parser_parser_ana_w_26_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_27_to_mem         (parser_parser_ana_w_27_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_28_to_mem         (parser_parser_ana_w_28_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_29_to_mem         (parser_parser_ana_w_29_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_2_to_mem          (parser_parser_ana_w_2_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_30_to_mem         (parser_parser_ana_w_30_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_31_to_mem         (parser_parser_ana_w_31_to_mem),                   
/* output logic   [54:0] */ .parser_parser_ana_w_3_to_mem          (parser_parser_ana_w_3_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_4_to_mem          (parser_parser_ana_w_4_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_5_to_mem          (parser_parser_ana_w_5_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_6_to_mem          (parser_parser_ana_w_6_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_7_to_mem          (parser_parser_ana_w_7_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_8_to_mem          (parser_parser_ana_w_8_to_mem),                    
/* output logic   [54:0] */ .parser_parser_ana_w_9_to_mem          (parser_parser_ana_w_9_to_mem),                    
/* output logic   [28:0] */ .parser_parser_csum_cfg_0_to_mem       (parser_parser_csum_cfg_0_to_mem),                 
/* output logic   [28:0] */ .parser_parser_csum_cfg_1_to_mem       (parser_parser_csum_cfg_1_to_mem),                 
/* output logic  [103:0] */ .parser_parser_extract_cfg_0_to_mem    (parser_parser_extract_cfg_0_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_10_to_mem   (parser_parser_extract_cfg_10_to_mem),             
/* output logic  [103:0] */ .parser_parser_extract_cfg_11_to_mem   (parser_parser_extract_cfg_11_to_mem),             
/* output logic  [103:0] */ .parser_parser_extract_cfg_12_to_mem   (parser_parser_extract_cfg_12_to_mem),             
/* output logic  [103:0] */ .parser_parser_extract_cfg_13_to_mem   (parser_parser_extract_cfg_13_to_mem),             
/* output logic  [103:0] */ .parser_parser_extract_cfg_14_to_mem   (parser_parser_extract_cfg_14_to_mem),             
/* output logic  [103:0] */ .parser_parser_extract_cfg_15_to_mem   (parser_parser_extract_cfg_15_to_mem),             
/* output logic  [103:0] */ .parser_parser_extract_cfg_1_to_mem    (parser_parser_extract_cfg_1_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_2_to_mem    (parser_parser_extract_cfg_2_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_3_to_mem    (parser_parser_extract_cfg_3_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_4_to_mem    (parser_parser_extract_cfg_4_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_5_to_mem    (parser_parser_extract_cfg_5_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_6_to_mem    (parser_parser_extract_cfg_6_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_7_to_mem    (parser_parser_extract_cfg_7_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_8_to_mem    (parser_parser_extract_cfg_8_to_mem),              
/* output logic  [103:0] */ .parser_parser_extract_cfg_9_to_mem    (parser_parser_extract_cfg_9_to_mem),              
/* output logic   [54:0] */ .parser_parser_key_s_0_to_mem          (parser_parser_key_s_0_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_10_to_mem         (parser_parser_key_s_10_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_11_to_mem         (parser_parser_key_s_11_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_12_to_mem         (parser_parser_key_s_12_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_13_to_mem         (parser_parser_key_s_13_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_14_to_mem         (parser_parser_key_s_14_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_15_to_mem         (parser_parser_key_s_15_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_16_to_mem         (parser_parser_key_s_16_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_17_to_mem         (parser_parser_key_s_17_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_18_to_mem         (parser_parser_key_s_18_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_19_to_mem         (parser_parser_key_s_19_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_1_to_mem          (parser_parser_key_s_1_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_20_to_mem         (parser_parser_key_s_20_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_21_to_mem         (parser_parser_key_s_21_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_22_to_mem         (parser_parser_key_s_22_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_23_to_mem         (parser_parser_key_s_23_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_24_to_mem         (parser_parser_key_s_24_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_25_to_mem         (parser_parser_key_s_25_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_26_to_mem         (parser_parser_key_s_26_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_27_to_mem         (parser_parser_key_s_27_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_28_to_mem         (parser_parser_key_s_28_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_29_to_mem         (parser_parser_key_s_29_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_2_to_mem          (parser_parser_key_s_2_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_30_to_mem         (parser_parser_key_s_30_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_31_to_mem         (parser_parser_key_s_31_to_mem),                   
/* output logic   [54:0] */ .parser_parser_key_s_3_to_mem          (parser_parser_key_s_3_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_4_to_mem          (parser_parser_key_s_4_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_5_to_mem          (parser_parser_key_s_5_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_6_to_mem          (parser_parser_key_s_6_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_7_to_mem          (parser_parser_key_s_7_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_8_to_mem          (parser_parser_key_s_8_to_mem),                    
/* output logic   [54:0] */ .parser_parser_key_s_9_to_mem          (parser_parser_key_s_9_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_0_to_mem          (parser_parser_key_w_0_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_10_to_mem         (parser_parser_key_w_10_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_11_to_mem         (parser_parser_key_w_11_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_12_to_mem         (parser_parser_key_w_12_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_13_to_mem         (parser_parser_key_w_13_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_17_to_mem         (parser_parser_key_w_17_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_18_to_mem         (parser_parser_key_w_18_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_19_to_mem         (parser_parser_key_w_19_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_1_to_mem          (parser_parser_key_w_1_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_20_to_mem         (parser_parser_key_w_20_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_21_to_mem         (parser_parser_key_w_21_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_22_to_mem         (parser_parser_key_w_22_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_23_to_mem         (parser_parser_key_w_23_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_24_to_mem         (parser_parser_key_w_24_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_25_to_mem         (parser_parser_key_w_25_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_26_to_mem         (parser_parser_key_w_26_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_27_to_mem         (parser_parser_key_w_27_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_28_to_mem         (parser_parser_key_w_28_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_29_to_mem         (parser_parser_key_w_29_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_2_to_mem          (parser_parser_key_w_2_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_30_to_mem         (parser_parser_key_w_30_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_31_to_mem         (parser_parser_key_w_31_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_3_to_mem          (parser_parser_key_w_3_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_4_to_mem          (parser_parser_key_w_4_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_5_to_mem          (parser_parser_key_w_5_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_6_to_mem          (parser_parser_key_w_6_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_7_to_mem          (parser_parser_key_w_7_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_8_to_mem          (parser_parser_key_w_8_to_mem),                    
/* output logic   [87:0] */ .parser_parser_key_w_9_to_mem          (parser_parser_key_w_9_to_mem),                    
/* output logic   [88:0] */ .parser_parser_metadata_fifo_to_mem    (parser_parser_metadata_fifo_to_mem),              
/* output logic   [89:0] */ .parser_parser_port_cfg_0_to_mem       (parser_parser_port_cfg_0_to_mem),                 
/* output logic   [89:0] */ .parser_parser_port_cfg_1_to_mem       (parser_parser_port_cfg_1_to_mem),                 
/* output logic   [34:0] */ .parser_parser_ptype_ram_to_mem        (parser_parser_ptype_ram_to_mem),                  
/* output logic          */ .parser_port_cfg_0_ecc_uncor_err       (),                                                
/* output logic          */ .parser_port_cfg_0_init_done           (),                                                
/* output logic   [63:0] */ .parser_port_cfg_0_rd_data             (),                                                
/* output logic          */ .parser_port_cfg_0_rd_valid            (),                                                
/* output logic          */ .parser_port_cfg_1_ecc_uncor_err       (),                                                
/* output logic          */ .parser_port_cfg_1_init_done           (),                                                
/* output logic   [63:0] */ .parser_port_cfg_1_rd_data             (),                                                
/* output logic          */ .parser_port_cfg_1_rd_valid            (),                                                
/* output logic          */ .parser_ptype_ram_ecc_uncor_err        (),                                                
/* output logic          */ .parser_ptype_ram_init_done            (),                                                
/* output logic   [13:0] */ .parser_ptype_ram_rd_data              (),                                                
/* output logic          */ .parser_ptype_ram_rd_valid             (),                                                
/* output logic          */ .unified_regs_ack                      (),                                                
/* output logic   [31:0] */ .unified_regs_rd_data                  (),                                                
/* output logic    [8:0] */ .parser_ana_exc_20_rd_data             (),                                                
/* output logic          */ .parser_ana_exc_20_rd_valid            (),                                                
/* output logic          */ .parser_ana_exc_21_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_exc_21_init_done           (),                                                
/* output logic          */ .parser_extract_cfg_5_ecc_uncor_err    (),                                                
/* output logic          */ .parser_extract_cfg_5_init_done        (),                                                
/* output logic   [79:0] */ .parser_extract_cfg_5_rd_data          (),                                                
/* output logic          */ .parser_extract_cfg_5_rd_valid         (),                                                
/* output logic   [95:0] */ .parser_ana_cam_2_rd_data              (),                                                
/* output logic          */ .parser_ana_cam_2_rd_valid             (),                                                
/* output logic          */ .parser_ana_cam_30_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_cam_30_init_done           (),                                                
/* output logic          */ .parser_key_w_15_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_w_15_init_done             (),                                                
/* output logic   [63:0] */ .parser_key_w_15_rd_data               (),                                                
/* output logic          */ .parser_key_w_15_rd_valid              (),                                                
/* output logic          */ .parser_key_w_6_ecc_uncor_err          (),                                                
/* output logic          */ .parser_key_w_6_init_done              (),                                                
/* output logic   [63:0] */ .parser_key_w_6_rd_data                (),                                                
/* output logic          */ .parser_key_w_6_rd_valid               (),                                                
/* output logic   [87:0] */ .parser_parser_key_w_14_to_mem         (parser_parser_key_w_14_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_15_to_mem         (parser_parser_key_w_15_to_mem),                   
/* output logic   [87:0] */ .parser_parser_key_w_16_to_mem         (parser_parser_key_w_16_to_mem),                   
/* output logic   [95:0] */ .parser_ana_cam_10_rd_data             (),                                                
/* output logic          */ .parser_ana_cam_10_rd_valid            (),                                                
/* output logic          */ .parser_ana_cam_11_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_10_rd_valid            (),                                                
/* output logic          */ .parser_ana_ext_11_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_11_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_11_rd_data             (),                                                
/* output logic          */ .parser_ana_ext_2_rd_valid             (),                                                
/* output logic          */ .parser_ana_ext_30_ecc_uncor_err       (),                                                
/* output logic          */ .parser_ana_ext_30_init_done           (),                                                
/* output logic   [25:0] */ .parser_ana_ext_30_rd_data             (),                                                
/* output logic          */ .parser_key_s_24_rd_valid              (),                                                
/* output logic          */ .parser_key_s_25_ecc_uncor_err         (),                                                
/* output logic          */ .parser_key_s_25_init_done             (),                                                
/* output logic   [31:0] */ .parser_key_s_25_rd_data               (),                                                
/* output logic          */ .parser_ana_w_11_ecc_uncor_err         (),                                                
/* output logic          */ .parser_ana_w_11_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_11_rd_data               (),                                                
/* output logic          */ .parser_ana_w_11_rd_valid              (),                                                
/* output logic          */ .parser_ana_w_31_init_done             (),                                                
/* output logic   [31:0] */ .parser_ana_w_31_rd_data               (),                                                
/* output logic          */ .parser_ana_w_31_rd_valid              ());                                                
// End of module parser_shells_wrapper from parser_shells_wrapper


// module parser_ff_mems    from parser_ff_mems using parser_ff_mems.map 
parser_ff_mems    parser_ff_mems(
/* input  logic          */ .cclk                                  (cclk),                                            
/* input  logic  [119:0] */ .parser_parser_ana_cam_10_to_mem       (parser_parser_ana_cam_10_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_0_to_mem        (parser_parser_ana_cam_0_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_11_to_mem       (parser_parser_ana_cam_11_to_mem),                 
/* input  logic          */ .car_raw_lan_power_good_with_byprst    (),                                                
/* input  logic  [119:0] */ .parser_parser_ana_cam_12_to_mem       (parser_parser_ana_cam_12_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_13_to_mem       (parser_parser_ana_cam_13_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_14_to_mem       (parser_parser_ana_cam_14_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_15_to_mem       (parser_parser_ana_cam_15_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_16_to_mem       (parser_parser_ana_cam_16_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_17_to_mem       (parser_parser_ana_cam_17_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_18_to_mem       (parser_parser_ana_cam_18_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_19_to_mem       (parser_parser_ana_cam_19_to_mem),                 
/* input  logic   [70:0] */ .parser_parser_ana_s_12_to_mem         (parser_parser_ana_s_12_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_13_to_mem         (parser_parser_ana_s_13_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_14_to_mem         (parser_parser_ana_s_14_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_15_to_mem         (parser_parser_ana_s_15_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_20_to_mem         (parser_parser_key_w_20_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_21_to_mem         (parser_parser_key_w_21_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_22_to_mem         (parser_parser_key_w_22_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_23_to_mem         (parser_parser_key_w_23_to_mem),                   
/* input  logic  [119:0] */ .parser_parser_ana_cam_1_to_mem        (parser_parser_ana_cam_1_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_20_to_mem       (parser_parser_ana_cam_20_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_21_to_mem       (parser_parser_ana_cam_21_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_22_to_mem       (parser_parser_ana_cam_22_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_23_to_mem       (parser_parser_ana_cam_23_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_24_to_mem       (parser_parser_ana_cam_24_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_25_to_mem       (parser_parser_ana_cam_25_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_26_to_mem       (parser_parser_ana_cam_26_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_27_to_mem       (parser_parser_ana_cam_27_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_28_to_mem       (parser_parser_ana_cam_28_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_29_to_mem       (parser_parser_ana_cam_29_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_2_to_mem        (parser_parser_ana_cam_2_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_30_to_mem       (parser_parser_ana_cam_30_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_31_to_mem       (parser_parser_ana_cam_31_to_mem),                 
/* input  logic  [119:0] */ .parser_parser_ana_cam_3_to_mem        (parser_parser_ana_cam_3_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_4_to_mem        (parser_parser_ana_cam_4_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_5_to_mem        (parser_parser_ana_cam_5_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_6_to_mem        (parser_parser_ana_cam_6_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_7_to_mem        (parser_parser_ana_cam_7_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_8_to_mem        (parser_parser_ana_cam_8_to_mem),                  
/* input  logic  [119:0] */ .parser_parser_ana_cam_9_to_mem        (parser_parser_ana_cam_9_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_0_to_mem        (parser_parser_ana_exc_0_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_10_to_mem       (parser_parser_ana_exc_10_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_11_to_mem       (parser_parser_ana_exc_11_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_12_to_mem       (parser_parser_ana_exc_12_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_13_to_mem       (parser_parser_ana_exc_13_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_14_to_mem       (parser_parser_ana_exc_14_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_15_to_mem       (parser_parser_ana_exc_15_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_16_to_mem       (parser_parser_ana_exc_16_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_17_to_mem       (parser_parser_ana_exc_17_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_18_to_mem       (parser_parser_ana_exc_18_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_19_to_mem       (parser_parser_ana_exc_19_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_1_to_mem        (parser_parser_ana_exc_1_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_20_to_mem       (parser_parser_ana_exc_20_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_21_to_mem       (parser_parser_ana_exc_21_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_22_to_mem       (parser_parser_ana_exc_22_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_23_to_mem       (parser_parser_ana_exc_23_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_24_to_mem       (parser_parser_ana_exc_24_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_25_to_mem       (parser_parser_ana_exc_25_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_26_to_mem       (parser_parser_ana_exc_26_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_27_to_mem       (parser_parser_ana_exc_27_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_28_to_mem       (parser_parser_ana_exc_28_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_29_to_mem       (parser_parser_ana_exc_29_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_2_to_mem        (parser_parser_ana_exc_2_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_30_to_mem       (parser_parser_ana_exc_30_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_31_to_mem       (parser_parser_ana_exc_31_to_mem),                 
/* input  logic   [29:0] */ .parser_parser_ana_exc_3_to_mem        (parser_parser_ana_exc_3_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_4_to_mem        (parser_parser_ana_exc_4_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_5_to_mem        (parser_parser_ana_exc_5_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_6_to_mem        (parser_parser_ana_exc_6_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_7_to_mem        (parser_parser_ana_exc_7_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_8_to_mem        (parser_parser_ana_exc_8_to_mem),                  
/* input  logic   [29:0] */ .parser_parser_ana_exc_9_to_mem        (parser_parser_ana_exc_9_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_0_to_mem        (parser_parser_ana_ext_0_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_10_to_mem       (parser_parser_ana_ext_10_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_11_to_mem       (parser_parser_ana_ext_11_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_12_to_mem       (parser_parser_ana_ext_12_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_13_to_mem       (parser_parser_ana_ext_13_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_14_to_mem       (parser_parser_ana_ext_14_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_15_to_mem       (parser_parser_ana_ext_15_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_16_to_mem       (parser_parser_ana_ext_16_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_17_to_mem       (parser_parser_ana_ext_17_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_18_to_mem       (parser_parser_ana_ext_18_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_19_to_mem       (parser_parser_ana_ext_19_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_1_to_mem        (parser_parser_ana_ext_1_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_20_to_mem       (parser_parser_ana_ext_20_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_21_to_mem       (parser_parser_ana_ext_21_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_22_to_mem       (parser_parser_ana_ext_22_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_23_to_mem       (parser_parser_ana_ext_23_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_24_to_mem       (parser_parser_ana_ext_24_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_25_to_mem       (parser_parser_ana_ext_25_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_26_to_mem       (parser_parser_ana_ext_26_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_27_to_mem       (parser_parser_ana_ext_27_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_28_to_mem       (parser_parser_ana_ext_28_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_29_to_mem       (parser_parser_ana_ext_29_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_2_to_mem        (parser_parser_ana_ext_2_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_30_to_mem       (parser_parser_ana_ext_30_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_31_to_mem       (parser_parser_ana_ext_31_to_mem),                 
/* input  logic   [49:0] */ .parser_parser_ana_ext_3_to_mem        (parser_parser_ana_ext_3_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_4_to_mem        (parser_parser_ana_ext_4_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_5_to_mem        (parser_parser_ana_ext_5_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_6_to_mem        (parser_parser_ana_ext_6_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_7_to_mem        (parser_parser_ana_ext_7_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_8_to_mem        (parser_parser_ana_ext_8_to_mem),                  
/* input  logic   [49:0] */ .parser_parser_ana_ext_9_to_mem        (parser_parser_ana_ext_9_to_mem),                  
/* input  logic   [70:0] */ .parser_parser_ana_s_0_to_mem          (parser_parser_ana_s_0_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_10_to_mem         (parser_parser_ana_s_10_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_11_to_mem         (parser_parser_ana_s_11_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_16_to_mem         (parser_parser_ana_s_16_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_17_to_mem         (parser_parser_ana_s_17_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_18_to_mem         (parser_parser_ana_s_18_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_19_to_mem         (parser_parser_ana_s_19_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_1_to_mem          (parser_parser_ana_s_1_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_20_to_mem         (parser_parser_ana_s_20_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_21_to_mem         (parser_parser_ana_s_21_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_22_to_mem         (parser_parser_ana_s_22_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_23_to_mem         (parser_parser_ana_s_23_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_24_to_mem         (parser_parser_ana_s_24_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_25_to_mem         (parser_parser_ana_s_25_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_26_to_mem         (parser_parser_ana_s_26_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_27_to_mem         (parser_parser_ana_s_27_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_28_to_mem         (parser_parser_ana_s_28_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_29_to_mem         (parser_parser_ana_s_29_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_2_to_mem          (parser_parser_ana_s_2_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_30_to_mem         (parser_parser_ana_s_30_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_31_to_mem         (parser_parser_ana_s_31_to_mem),                   
/* input  logic   [70:0] */ .parser_parser_ana_s_3_to_mem          (parser_parser_ana_s_3_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_4_to_mem          (parser_parser_ana_s_4_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_5_to_mem          (parser_parser_ana_s_5_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_6_to_mem          (parser_parser_ana_s_6_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_7_to_mem          (parser_parser_ana_s_7_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_8_to_mem          (parser_parser_ana_s_8_to_mem),                    
/* input  logic   [70:0] */ .parser_parser_ana_s_9_to_mem          (parser_parser_ana_s_9_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_0_to_mem          (parser_parser_ana_w_0_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_10_to_mem         (parser_parser_ana_w_10_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_11_to_mem         (parser_parser_ana_w_11_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_12_to_mem         (parser_parser_ana_w_12_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_13_to_mem         (parser_parser_ana_w_13_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_14_to_mem         (parser_parser_ana_w_14_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_15_to_mem         (parser_parser_ana_w_15_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_16_to_mem         (parser_parser_ana_w_16_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_17_to_mem         (parser_parser_ana_w_17_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_18_to_mem         (parser_parser_ana_w_18_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_19_to_mem         (parser_parser_ana_w_19_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_1_to_mem          (parser_parser_ana_w_1_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_20_to_mem         (parser_parser_ana_w_20_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_21_to_mem         (parser_parser_ana_w_21_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_22_to_mem         (parser_parser_ana_w_22_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_23_to_mem         (parser_parser_ana_w_23_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_24_to_mem         (parser_parser_ana_w_24_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_25_to_mem         (parser_parser_ana_w_25_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_26_to_mem         (parser_parser_ana_w_26_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_27_to_mem         (parser_parser_ana_w_27_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_28_to_mem         (parser_parser_ana_w_28_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_29_to_mem         (parser_parser_ana_w_29_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_2_to_mem          (parser_parser_ana_w_2_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_30_to_mem         (parser_parser_ana_w_30_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_31_to_mem         (parser_parser_ana_w_31_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_ana_w_3_to_mem          (parser_parser_ana_w_3_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_4_to_mem          (parser_parser_ana_w_4_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_5_to_mem          (parser_parser_ana_w_5_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_6_to_mem          (parser_parser_ana_w_6_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_7_to_mem          (parser_parser_ana_w_7_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_8_to_mem          (parser_parser_ana_w_8_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_ana_w_9_to_mem          (parser_parser_ana_w_9_to_mem),                    
/* input  logic   [28:0] */ .parser_parser_csum_cfg_0_to_mem       (parser_parser_csum_cfg_0_to_mem),                 
/* input  logic   [28:0] */ .parser_parser_csum_cfg_1_to_mem       (parser_parser_csum_cfg_1_to_mem),                 
/* input  logic  [103:0] */ .parser_parser_extract_cfg_0_to_mem    (parser_parser_extract_cfg_0_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_10_to_mem   (parser_parser_extract_cfg_10_to_mem),             
/* input  logic  [103:0] */ .parser_parser_extract_cfg_11_to_mem   (parser_parser_extract_cfg_11_to_mem),             
/* input  logic  [103:0] */ .parser_parser_extract_cfg_12_to_mem   (parser_parser_extract_cfg_12_to_mem),             
/* input  logic  [103:0] */ .parser_parser_extract_cfg_13_to_mem   (parser_parser_extract_cfg_13_to_mem),             
/* input  logic  [103:0] */ .parser_parser_extract_cfg_14_to_mem   (parser_parser_extract_cfg_14_to_mem),             
/* input  logic  [103:0] */ .parser_parser_extract_cfg_15_to_mem   (parser_parser_extract_cfg_15_to_mem),             
/* input  logic  [103:0] */ .parser_parser_extract_cfg_1_to_mem    (parser_parser_extract_cfg_1_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_2_to_mem    (parser_parser_extract_cfg_2_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_3_to_mem    (parser_parser_extract_cfg_3_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_4_to_mem    (parser_parser_extract_cfg_4_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_5_to_mem    (parser_parser_extract_cfg_5_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_6_to_mem    (parser_parser_extract_cfg_6_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_7_to_mem    (parser_parser_extract_cfg_7_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_8_to_mem    (parser_parser_extract_cfg_8_to_mem),              
/* input  logic  [103:0] */ .parser_parser_extract_cfg_9_to_mem    (parser_parser_extract_cfg_9_to_mem),              
/* input  logic   [54:0] */ .parser_parser_key_s_0_to_mem          (parser_parser_key_s_0_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_10_to_mem         (parser_parser_key_s_10_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_11_to_mem         (parser_parser_key_s_11_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_12_to_mem         (parser_parser_key_s_12_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_13_to_mem         (parser_parser_key_s_13_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_14_to_mem         (parser_parser_key_s_14_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_15_to_mem         (parser_parser_key_s_15_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_16_to_mem         (parser_parser_key_s_16_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_17_to_mem         (parser_parser_key_s_17_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_18_to_mem         (parser_parser_key_s_18_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_19_to_mem         (parser_parser_key_s_19_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_1_to_mem          (parser_parser_key_s_1_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_20_to_mem         (parser_parser_key_s_20_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_21_to_mem         (parser_parser_key_s_21_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_22_to_mem         (parser_parser_key_s_22_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_23_to_mem         (parser_parser_key_s_23_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_24_to_mem         (parser_parser_key_s_24_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_25_to_mem         (parser_parser_key_s_25_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_26_to_mem         (parser_parser_key_s_26_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_27_to_mem         (parser_parser_key_s_27_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_28_to_mem         (parser_parser_key_s_28_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_29_to_mem         (parser_parser_key_s_29_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_2_to_mem          (parser_parser_key_s_2_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_30_to_mem         (parser_parser_key_s_30_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_31_to_mem         (parser_parser_key_s_31_to_mem),                   
/* input  logic   [54:0] */ .parser_parser_key_s_3_to_mem          (parser_parser_key_s_3_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_4_to_mem          (parser_parser_key_s_4_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_5_to_mem          (parser_parser_key_s_5_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_6_to_mem          (parser_parser_key_s_6_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_7_to_mem          (parser_parser_key_s_7_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_8_to_mem          (parser_parser_key_s_8_to_mem),                    
/* input  logic   [54:0] */ .parser_parser_key_s_9_to_mem          (parser_parser_key_s_9_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_0_to_mem          (parser_parser_key_w_0_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_10_to_mem         (parser_parser_key_w_10_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_11_to_mem         (parser_parser_key_w_11_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_12_to_mem         (parser_parser_key_w_12_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_13_to_mem         (parser_parser_key_w_13_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_14_to_mem         (parser_parser_key_w_14_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_15_to_mem         (parser_parser_key_w_15_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_16_to_mem         (parser_parser_key_w_16_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_17_to_mem         (parser_parser_key_w_17_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_18_to_mem         (parser_parser_key_w_18_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_19_to_mem         (parser_parser_key_w_19_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_1_to_mem          (parser_parser_key_w_1_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_24_to_mem         (parser_parser_key_w_24_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_25_to_mem         (parser_parser_key_w_25_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_26_to_mem         (parser_parser_key_w_26_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_27_to_mem         (parser_parser_key_w_27_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_28_to_mem         (parser_parser_key_w_28_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_29_to_mem         (parser_parser_key_w_29_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_2_to_mem          (parser_parser_key_w_2_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_30_to_mem         (parser_parser_key_w_30_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_31_to_mem         (parser_parser_key_w_31_to_mem),                   
/* input  logic   [87:0] */ .parser_parser_key_w_3_to_mem          (parser_parser_key_w_3_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_4_to_mem          (parser_parser_key_w_4_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_5_to_mem          (parser_parser_key_w_5_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_6_to_mem          (parser_parser_key_w_6_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_7_to_mem          (parser_parser_key_w_7_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_8_to_mem          (parser_parser_key_w_8_to_mem),                    
/* input  logic   [87:0] */ .parser_parser_key_w_9_to_mem          (parser_parser_key_w_9_to_mem),                    
/* input  logic   [88:0] */ .parser_parser_metadata_fifo_to_mem    (parser_parser_metadata_fifo_to_mem),              
/* input  logic   [89:0] */ .parser_parser_port_cfg_0_to_mem       (parser_parser_port_cfg_0_to_mem),                 
/* input  logic   [89:0] */ .parser_parser_port_cfg_1_to_mem       (parser_parser_port_cfg_1_to_mem),                 
/* input  logic   [34:0] */ .parser_parser_ptype_ram_to_mem        (parser_parser_ptype_ram_to_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_13_from_mem       (parser_parser_key_w_13_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_14_from_mem       (parser_parser_key_w_14_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_15_from_mem       (parser_parser_key_w_15_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_16_from_mem       (parser_parser_key_w_16_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_17_from_mem       (parser_parser_key_w_17_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_18_from_mem       (parser_parser_key_w_18_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_19_from_mem       (parser_parser_key_w_19_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_1_from_mem        (parser_parser_key_w_1_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_20_from_mem       (parser_parser_key_w_20_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_21_from_mem       (parser_parser_key_w_21_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_22_from_mem       (parser_parser_key_w_22_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_23_from_mem       (parser_parser_key_w_23_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_24_from_mem       (parser_parser_key_w_24_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_25_from_mem       (parser_parser_key_w_25_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_26_from_mem       (parser_parser_key_w_26_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_30_from_mem       (parser_parser_key_w_30_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_31_from_mem       (parser_parser_key_w_31_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_3_from_mem        (parser_parser_key_w_3_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_4_from_mem        (parser_parser_key_w_4_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_5_from_mem        (parser_parser_key_w_5_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_6_from_mem        (parser_parser_key_w_6_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_7_from_mem        (parser_parser_key_w_7_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_8_from_mem        (parser_parser_key_w_8_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_9_from_mem        (parser_parser_key_w_9_from_mem),                  
/* output logic   [69:0] */ .parser_parser_metadata_fifo_from_mem  (parser_parser_metadata_fifo_from_mem),            
/* output logic   [72:0] */ .parser_parser_port_cfg_0_from_mem     (parser_parser_port_cfg_0_from_mem),               
/* output logic   [72:0] */ .parser_parser_port_cfg_1_from_mem     (parser_parser_port_cfg_1_from_mem),               
/* output logic   [20:0] */ .parser_parser_ptype_ram_from_mem      (parser_parser_ptype_ram_from_mem),                
/* output logic   [55:0] */ .parser_parser_ana_s_16_from_mem       (parser_parser_ana_s_16_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_17_from_mem       (parser_parser_ana_s_17_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_18_from_mem       (parser_parser_ana_s_18_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_27_from_mem       (parser_parser_key_w_27_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_28_from_mem       (parser_parser_key_w_28_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_29_from_mem       (parser_parser_key_w_29_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_2_from_mem        (parser_parser_key_w_2_from_mem),                  
/* output logic  [104:0] */ .parser_parser_ana_cam_0_from_mem      (parser_parser_ana_cam_0_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_10_from_mem     (parser_parser_ana_cam_10_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_11_from_mem     (parser_parser_ana_cam_11_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_12_from_mem     (parser_parser_ana_cam_12_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_13_from_mem     (parser_parser_ana_cam_13_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_14_from_mem     (parser_parser_ana_cam_14_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_15_from_mem     (parser_parser_ana_cam_15_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_16_from_mem     (parser_parser_ana_cam_16_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_17_from_mem     (parser_parser_ana_cam_17_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_18_from_mem     (parser_parser_ana_cam_18_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_19_from_mem     (parser_parser_ana_cam_19_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_1_from_mem      (parser_parser_ana_cam_1_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_20_from_mem     (parser_parser_ana_cam_20_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_21_from_mem     (parser_parser_ana_cam_21_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_22_from_mem     (parser_parser_ana_cam_22_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_23_from_mem     (parser_parser_ana_cam_23_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_24_from_mem     (parser_parser_ana_cam_24_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_25_from_mem     (parser_parser_ana_cam_25_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_26_from_mem     (parser_parser_ana_cam_26_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_27_from_mem     (parser_parser_ana_cam_27_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_28_from_mem     (parser_parser_ana_cam_28_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_29_from_mem     (parser_parser_ana_cam_29_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_2_from_mem      (parser_parser_ana_cam_2_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_30_from_mem     (parser_parser_ana_cam_30_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_31_from_mem     (parser_parser_ana_cam_31_from_mem),               
/* output logic  [104:0] */ .parser_parser_ana_cam_3_from_mem      (parser_parser_ana_cam_3_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_4_from_mem      (parser_parser_ana_cam_4_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_5_from_mem      (parser_parser_ana_cam_5_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_6_from_mem      (parser_parser_ana_cam_6_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_7_from_mem      (parser_parser_ana_cam_7_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_8_from_mem      (parser_parser_ana_cam_8_from_mem),                
/* output logic  [104:0] */ .parser_parser_ana_cam_9_from_mem      (parser_parser_ana_cam_9_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_0_from_mem      (parser_parser_ana_exc_0_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_10_from_mem     (parser_parser_ana_exc_10_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_11_from_mem     (parser_parser_ana_exc_11_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_12_from_mem     (parser_parser_ana_exc_12_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_13_from_mem     (parser_parser_ana_exc_13_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_14_from_mem     (parser_parser_ana_exc_14_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_15_from_mem     (parser_parser_ana_exc_15_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_16_from_mem     (parser_parser_ana_exc_16_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_17_from_mem     (parser_parser_ana_exc_17_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_18_from_mem     (parser_parser_ana_exc_18_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_19_from_mem     (parser_parser_ana_exc_19_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_1_from_mem      (parser_parser_ana_exc_1_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_20_from_mem     (parser_parser_ana_exc_20_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_21_from_mem     (parser_parser_ana_exc_21_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_22_from_mem     (parser_parser_ana_exc_22_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_23_from_mem     (parser_parser_ana_exc_23_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_24_from_mem     (parser_parser_ana_exc_24_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_25_from_mem     (parser_parser_ana_exc_25_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_26_from_mem     (parser_parser_ana_exc_26_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_27_from_mem     (parser_parser_ana_exc_27_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_28_from_mem     (parser_parser_ana_exc_28_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_29_from_mem     (parser_parser_ana_exc_29_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_2_from_mem      (parser_parser_ana_exc_2_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_30_from_mem     (parser_parser_ana_exc_30_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_31_from_mem     (parser_parser_ana_exc_31_from_mem),               
/* output logic   [14:0] */ .parser_parser_ana_exc_3_from_mem      (parser_parser_ana_exc_3_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_4_from_mem      (parser_parser_ana_exc_4_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_5_from_mem      (parser_parser_ana_exc_5_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_6_from_mem      (parser_parser_ana_exc_6_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_7_from_mem      (parser_parser_ana_exc_7_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_8_from_mem      (parser_parser_ana_exc_8_from_mem),                
/* output logic   [14:0] */ .parser_parser_ana_exc_9_from_mem      (parser_parser_ana_exc_9_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_0_from_mem      (parser_parser_ana_ext_0_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_10_from_mem     (parser_parser_ana_ext_10_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_11_from_mem     (parser_parser_ana_ext_11_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_12_from_mem     (parser_parser_ana_ext_12_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_13_from_mem     (parser_parser_ana_ext_13_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_14_from_mem     (parser_parser_ana_ext_14_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_15_from_mem     (parser_parser_ana_ext_15_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_16_from_mem     (parser_parser_ana_ext_16_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_17_from_mem     (parser_parser_ana_ext_17_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_18_from_mem     (parser_parser_ana_ext_18_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_19_from_mem     (parser_parser_ana_ext_19_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_1_from_mem      (parser_parser_ana_ext_1_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_20_from_mem     (parser_parser_ana_ext_20_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_21_from_mem     (parser_parser_ana_ext_21_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_22_from_mem     (parser_parser_ana_ext_22_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_23_from_mem     (parser_parser_ana_ext_23_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_24_from_mem     (parser_parser_ana_ext_24_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_25_from_mem     (parser_parser_ana_ext_25_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_26_from_mem     (parser_parser_ana_ext_26_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_27_from_mem     (parser_parser_ana_ext_27_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_28_from_mem     (parser_parser_ana_ext_28_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_29_from_mem     (parser_parser_ana_ext_29_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_2_from_mem      (parser_parser_ana_ext_2_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_30_from_mem     (parser_parser_ana_ext_30_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_31_from_mem     (parser_parser_ana_ext_31_from_mem),               
/* output logic   [32:0] */ .parser_parser_ana_ext_3_from_mem      (parser_parser_ana_ext_3_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_4_from_mem      (parser_parser_ana_ext_4_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_5_from_mem      (parser_parser_ana_ext_5_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_6_from_mem      (parser_parser_ana_ext_6_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_7_from_mem      (parser_parser_ana_ext_7_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_8_from_mem      (parser_parser_ana_ext_8_from_mem),                
/* output logic   [32:0] */ .parser_parser_ana_ext_9_from_mem      (parser_parser_ana_ext_9_from_mem),                
/* output logic   [55:0] */ .parser_parser_ana_s_0_from_mem        (parser_parser_ana_s_0_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_10_from_mem       (parser_parser_ana_s_10_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_11_from_mem       (parser_parser_ana_s_11_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_12_from_mem       (parser_parser_ana_s_12_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_13_from_mem       (parser_parser_ana_s_13_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_14_from_mem       (parser_parser_ana_s_14_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_15_from_mem       (parser_parser_ana_s_15_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_19_from_mem       (parser_parser_ana_s_19_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_1_from_mem        (parser_parser_ana_s_1_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_20_from_mem       (parser_parser_ana_s_20_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_21_from_mem       (parser_parser_ana_s_21_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_22_from_mem       (parser_parser_ana_s_22_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_23_from_mem       (parser_parser_ana_s_23_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_24_from_mem       (parser_parser_ana_s_24_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_25_from_mem       (parser_parser_ana_s_25_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_26_from_mem       (parser_parser_ana_s_26_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_27_from_mem       (parser_parser_ana_s_27_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_28_from_mem       (parser_parser_ana_s_28_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_29_from_mem       (parser_parser_ana_s_29_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_2_from_mem        (parser_parser_ana_s_2_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_30_from_mem       (parser_parser_ana_s_30_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_31_from_mem       (parser_parser_ana_s_31_from_mem),                 
/* output logic   [55:0] */ .parser_parser_ana_s_3_from_mem        (parser_parser_ana_s_3_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_4_from_mem        (parser_parser_ana_s_4_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_5_from_mem        (parser_parser_ana_s_5_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_6_from_mem        (parser_parser_ana_s_6_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_7_from_mem        (parser_parser_ana_s_7_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_8_from_mem        (parser_parser_ana_s_8_from_mem),                  
/* output logic   [55:0] */ .parser_parser_ana_s_9_from_mem        (parser_parser_ana_s_9_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_0_from_mem        (parser_parser_ana_w_0_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_10_from_mem       (parser_parser_ana_w_10_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_11_from_mem       (parser_parser_ana_w_11_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_12_from_mem       (parser_parser_ana_w_12_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_13_from_mem       (parser_parser_ana_w_13_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_14_from_mem       (parser_parser_ana_w_14_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_15_from_mem       (parser_parser_ana_w_15_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_16_from_mem       (parser_parser_ana_w_16_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_17_from_mem       (parser_parser_ana_w_17_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_18_from_mem       (parser_parser_ana_w_18_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_19_from_mem       (parser_parser_ana_w_19_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_1_from_mem        (parser_parser_ana_w_1_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_20_from_mem       (parser_parser_ana_w_20_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_21_from_mem       (parser_parser_ana_w_21_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_22_from_mem       (parser_parser_ana_w_22_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_23_from_mem       (parser_parser_ana_w_23_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_24_from_mem       (parser_parser_ana_w_24_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_25_from_mem       (parser_parser_ana_w_25_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_26_from_mem       (parser_parser_ana_w_26_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_27_from_mem       (parser_parser_ana_w_27_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_28_from_mem       (parser_parser_ana_w_28_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_29_from_mem       (parser_parser_ana_w_29_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_2_from_mem        (parser_parser_ana_w_2_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_30_from_mem       (parser_parser_ana_w_30_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_31_from_mem       (parser_parser_ana_w_31_from_mem),                 
/* output logic   [39:0] */ .parser_parser_ana_w_3_from_mem        (parser_parser_ana_w_3_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_4_from_mem        (parser_parser_ana_w_4_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_5_from_mem        (parser_parser_ana_w_5_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_6_from_mem        (parser_parser_ana_w_6_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_7_from_mem        (parser_parser_ana_w_7_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_8_from_mem        (parser_parser_ana_w_8_from_mem),                  
/* output logic   [39:0] */ .parser_parser_ana_w_9_from_mem        (parser_parser_ana_w_9_from_mem),                  
/* output logic   [11:0] */ .parser_parser_csum_cfg_0_from_mem     (parser_parser_csum_cfg_0_from_mem),               
/* output logic   [11:0] */ .parser_parser_csum_cfg_1_from_mem     (parser_parser_csum_cfg_1_from_mem),               
/* output logic   [88:0] */ .parser_parser_extract_cfg_0_from_mem  (parser_parser_extract_cfg_0_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_10_from_mem (parser_parser_extract_cfg_10_from_mem),           
/* output logic   [88:0] */ .parser_parser_extract_cfg_11_from_mem (parser_parser_extract_cfg_11_from_mem),           
/* output logic   [88:0] */ .parser_parser_extract_cfg_12_from_mem (parser_parser_extract_cfg_12_from_mem),           
/* output logic   [88:0] */ .parser_parser_extract_cfg_13_from_mem (parser_parser_extract_cfg_13_from_mem),           
/* output logic   [88:0] */ .parser_parser_extract_cfg_14_from_mem (parser_parser_extract_cfg_14_from_mem),           
/* output logic   [88:0] */ .parser_parser_extract_cfg_15_from_mem (parser_parser_extract_cfg_15_from_mem),           
/* output logic   [88:0] */ .parser_parser_extract_cfg_1_from_mem  (parser_parser_extract_cfg_1_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_2_from_mem  (parser_parser_extract_cfg_2_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_3_from_mem  (parser_parser_extract_cfg_3_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_4_from_mem  (parser_parser_extract_cfg_4_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_5_from_mem  (parser_parser_extract_cfg_5_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_6_from_mem  (parser_parser_extract_cfg_6_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_7_from_mem  (parser_parser_extract_cfg_7_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_8_from_mem  (parser_parser_extract_cfg_8_from_mem),            
/* output logic   [88:0] */ .parser_parser_extract_cfg_9_from_mem  (parser_parser_extract_cfg_9_from_mem),            
/* output logic   [39:0] */ .parser_parser_key_s_0_from_mem        (parser_parser_key_s_0_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_10_from_mem       (parser_parser_key_s_10_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_11_from_mem       (parser_parser_key_s_11_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_12_from_mem       (parser_parser_key_s_12_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_13_from_mem       (parser_parser_key_s_13_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_14_from_mem       (parser_parser_key_s_14_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_15_from_mem       (parser_parser_key_s_15_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_16_from_mem       (parser_parser_key_s_16_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_17_from_mem       (parser_parser_key_s_17_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_18_from_mem       (parser_parser_key_s_18_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_19_from_mem       (parser_parser_key_s_19_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_1_from_mem        (parser_parser_key_s_1_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_20_from_mem       (parser_parser_key_s_20_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_21_from_mem       (parser_parser_key_s_21_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_22_from_mem       (parser_parser_key_s_22_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_23_from_mem       (parser_parser_key_s_23_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_24_from_mem       (parser_parser_key_s_24_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_25_from_mem       (parser_parser_key_s_25_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_26_from_mem       (parser_parser_key_s_26_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_27_from_mem       (parser_parser_key_s_27_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_28_from_mem       (parser_parser_key_s_28_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_29_from_mem       (parser_parser_key_s_29_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_2_from_mem        (parser_parser_key_s_2_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_30_from_mem       (parser_parser_key_s_30_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_31_from_mem       (parser_parser_key_s_31_from_mem),                 
/* output logic   [39:0] */ .parser_parser_key_s_3_from_mem        (parser_parser_key_s_3_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_4_from_mem        (parser_parser_key_s_4_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_5_from_mem        (parser_parser_key_s_5_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_6_from_mem        (parser_parser_key_s_6_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_7_from_mem        (parser_parser_key_s_7_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_8_from_mem        (parser_parser_key_s_8_from_mem),                  
/* output logic   [39:0] */ .parser_parser_key_s_9_from_mem        (parser_parser_key_s_9_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_0_from_mem        (parser_parser_key_w_0_from_mem),                  
/* output logic   [72:0] */ .parser_parser_key_w_10_from_mem       (parser_parser_key_w_10_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_11_from_mem       (parser_parser_key_w_11_from_mem),                 
/* output logic   [72:0] */ .parser_parser_key_w_12_from_mem       (parser_parser_key_w_12_from_mem));                 
// End of module parser_ff_mems from parser_ff_mems

endmodule // parser_top
