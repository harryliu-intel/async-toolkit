magic
tech scmos
timestamp 988943070
<< nselect >>
rect -60 -75 0 16
<< pselect >>
rect 0 -68 40 8
<< ndiffusion >>
rect -40 4 -8 5
rect -40 0 -8 1
rect -40 -8 -28 0
rect -40 -9 -8 -8
rect -40 -13 -8 -12
rect -40 -22 -8 -21
rect -40 -26 -8 -25
rect -40 -34 -28 -26
rect -40 -35 -8 -34
rect -40 -39 -8 -38
rect -40 -48 -8 -47
rect -40 -52 -8 -51
rect -40 -60 -28 -52
rect -40 -61 -8 -60
rect -40 -65 -8 -64
<< pdiffusion >>
rect 8 -6 28 -5
rect 8 -14 28 -9
rect 8 -22 28 -17
rect 8 -26 28 -25
rect 8 -35 28 -34
rect 8 -43 28 -38
rect 8 -51 28 -46
rect 8 -55 28 -54
<< ntransistor >>
rect -40 1 -8 4
rect -40 -12 -8 -9
rect -40 -25 -8 -22
rect -40 -38 -8 -35
rect -40 -51 -8 -48
rect -40 -64 -8 -61
<< ptransistor >>
rect 8 -9 28 -6
rect 8 -17 28 -14
rect 8 -25 28 -22
rect 8 -38 28 -35
rect 8 -46 28 -43
rect 8 -54 28 -51
<< polysilicon >>
rect -52 1 -40 4
rect -8 1 6 4
rect 3 -6 6 1
rect 3 -9 8 -6
rect 28 -9 32 -6
rect -44 -12 -40 -9
rect -8 -12 -3 -9
rect -6 -14 -3 -12
rect -6 -17 8 -14
rect 28 -17 32 -14
rect -44 -25 -40 -22
rect -8 -25 8 -22
rect 28 -25 32 -22
rect -52 -38 -40 -35
rect -8 -38 8 -35
rect 28 -38 32 -35
rect -6 -46 8 -43
rect 28 -46 32 -43
rect -6 -48 -3 -46
rect -44 -51 -40 -48
rect -8 -51 -3 -48
rect 3 -54 8 -51
rect 28 -54 32 -51
rect 3 -61 6 -54
rect -44 -64 -40 -61
rect -8 -64 6 -61
<< ndcontact >>
rect -40 5 -8 13
rect -28 -8 -8 0
rect -40 -21 -8 -13
rect -28 -34 -8 -26
rect -40 -47 -8 -39
rect -28 -60 -8 -52
rect -40 -73 -8 -65
<< pdcontact >>
rect 8 -5 28 3
rect 8 -34 28 -26
rect 8 -63 28 -55
<< polycontact >>
rect -60 -4 -52 4
rect -52 -17 -44 -9
rect -60 -38 -52 -30
rect 32 -30 40 -22
rect -52 -56 -44 -48
rect 32 -59 40 -51
<< metal1 >>
rect -40 5 -8 13
rect -60 -4 -52 4
rect -60 -30 -56 -4
rect -52 -17 -44 -9
rect -60 -38 -52 -30
rect -48 -48 -44 -17
rect -52 -56 -44 -48
rect -40 -13 -32 5
rect -28 -8 4 0
rect 8 -5 28 3
rect -40 -21 -8 -13
rect -40 -39 -32 -21
rect -4 -26 4 -8
rect -28 -34 28 -26
rect -40 -47 -8 -39
rect -40 -65 -32 -47
rect -4 -52 4 -34
rect -28 -60 4 -52
rect 8 -63 28 -55
rect 32 -59 40 -22
rect -40 -73 -8 -65
<< labels >>
rlabel metal1 32 -59 40 -22 7 a
rlabel metal1 -48 -56 -44 -9 1 b
rlabel metal1 -60 -38 -56 4 3 c
rlabel space -61 -75 -28 16 7 ^n
rlabel space 28 -68 41 8 3 ^p
rlabel metal1 -40 -47 -8 -39 1 GND!|pin|s|0
rlabel metal1 -40 -73 -32 13 1 GND!|pin|s|0
rlabel metal1 8 -5 28 3 1 Vdd!|pin|s|1
rlabel metal1 -4 -60 4 0 1 x|pin|s|2
rlabel metal1 -28 -8 4 0 1 x|pin|s|2
rlabel metal1 -28 -60 4 -52 1 x|pin|s|2
rlabel metal1 -28 -34 28 -26 1 x|pin|s|2
rlabel metal1 -40 5 -8 13 1 GND!|pin|s|0
rlabel metal1 -40 -21 -8 -13 1 GND!|pin|s|0
rlabel metal1 -40 -73 -8 -65 1 GND!|pin|s|0
rlabel metal1 8 -63 28 -55 1 Vdd!|pin|s|0
<< end >>
