// vim: noai : ts=3 : sw=3 : expandtab : ft=systemverilog

//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors.  The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//=======================================================================
// COPYRIGHT (C)  2012 SYNOPSYS INC.
// This software and the associated documentation are confidential and
// proprietary to Synopsys, Inc. Your use or disclosure of this software
// is subject to the terms and conditions of a written license agreement
// between you, or your company, and Synopsys, Inc. In the event of
// publications, the following notice is applicable:
//
// ALL RIGHTS RESERVED
//
// The entire notice above must be reproduced on all authorized copies.
//
//------------------------------------------------------------------------------
//   Author        : Dhivya Sankar
//   Project       : Madison Bay
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Class : ahb_master_directed_sequence 
// ahb_master_directed_sequence is used by test to provide initiator
// scenario information to the Master agent present in the System Env.
// This class defines a sequence in which a AHB WRITE followed by a AHB READ
// sequence is generated by assigning values to the transactions rather than
// randomization, and then transmitted using `uvm_send.
//------------------------------------------------------------------------------

`ifndef GUARD_AHB_MASTER_DIRECTED_SEQUENCE_SV
`define GUARD_AHB_MASTER_DIRECTED_SEQUENCE_SV

class ahb_master_directed_sequence extends svt_ahb_master_transaction_base_sequence;

   `uvm_object_utils(ahb_master_directed_sequence)

  svt_ahb_master_transaction write_tran, read_tran;
  svt_configuration get_cfg;
  bit status;

  /** Class Constructor */
  function new(string name="ahb_master_directed_sequence");
    super.new(name);
  endfunction
  
  virtual task body();
    
    `uvm_info("body", "Entered ...", UVM_LOW)

    super.body();

    /** Obtain a handle to the port configuration */
    p_sequencer.get_cfg(get_cfg);
    if (!$cast(cfg, get_cfg)) begin
      `uvm_fatal("body", "Unable to $cast the configuration to a svt_ahb_port_configuration class");
    end

      /** Set up the write transaction */
      `uvm_create(write_tran)
      write_tran.randomize()with {
      write_tran.lock         == 0;
      write_tran.cfg          == cfg;
      write_tran.xact_type    == svt_ahb_transaction::WRITE;
      write_tran.addr         == (32'h0000_0000 | ('h10 * 1));
      write_tran.burst_type   == svt_ahb_transaction::INCR4;
      write_tran.burst_size   == svt_ahb_transaction::BURST_SIZE_32BIT;
      write_tran.data[0] == 1;
      };
       
      `uvm_send(write_tran)
      get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm write sequence received:\n%s",rsp.sprint()));
 

    `uvm_info("body", "Exiting...", UVM_LOW)
  endtask: body

endclass: ahb_master_directed_sequence

`endif // GUARD_AHB_MASTER_DIRECTED_SEQUENCE_SV
