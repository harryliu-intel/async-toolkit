magic
tech scmos
timestamp 988943070
<< nselect >>
rect -52 -21 0 35
<< pselect >>
rect 0 -21 75 35
<< ndiffusion >>
rect -25 22 -13 23
rect -25 14 -13 19
rect -25 10 -13 11
rect -25 2 -23 10
rect -25 1 -13 2
rect -47 -7 -39 -6
rect -25 -7 -13 -2
rect -47 -11 -39 -10
rect -25 -11 -13 -10
<< pdiffusion >>
rect 8 22 28 23
rect 59 21 63 24
rect 8 14 28 19
rect 8 10 28 11
rect 8 1 28 2
rect 59 15 63 18
rect 8 -7 28 -2
rect 57 -7 65 -6
rect 8 -11 28 -10
rect 57 -11 65 -10
<< ntransistor >>
rect -25 19 -13 22
rect -25 11 -13 14
rect -25 -2 -13 1
rect -47 -10 -39 -7
rect -25 -10 -13 -7
<< ptransistor >>
rect 8 19 28 22
rect 8 11 28 14
rect 59 18 63 21
rect 8 -2 28 1
rect 8 -10 28 -7
rect 57 -10 65 -7
<< polysilicon >>
rect -29 19 -25 22
rect -13 19 -4 22
rect 4 19 8 22
rect 28 19 40 22
rect -30 11 -25 14
rect -13 11 -9 14
rect -4 11 8 14
rect 28 11 32 14
rect -52 -7 -49 10
rect -30 6 -27 11
rect -27 -2 -25 1
rect -13 -2 -9 1
rect -4 -7 -1 11
rect 37 1 40 19
rect 55 18 59 21
rect 63 18 67 21
rect 4 -2 8 1
rect 28 -2 40 1
rect 50 -7 53 2
rect -52 -10 -47 -7
rect -39 -10 -35 -7
rect -29 -10 -25 -7
rect -13 -10 8 -7
rect 28 -10 32 -7
rect 50 -10 57 -7
rect 65 -10 69 -7
<< ndcontact >>
rect -25 23 -13 31
rect -47 -6 -39 2
rect -23 2 -13 10
rect -47 -19 -39 -11
rect -25 -19 -13 -11
<< pdcontact >>
rect 8 23 28 31
rect 55 24 63 32
rect 8 2 28 10
rect 55 7 63 15
rect 57 -6 65 2
rect 8 -19 28 -11
rect 57 -19 65 -11
<< polycontact >>
rect -4 19 4 27
rect -52 10 -44 18
rect -35 -2 -27 6
rect 45 2 53 10
rect 67 13 75 21
rect -4 -18 4 -10
<< metal1 >>
rect 55 31 63 32
rect -25 23 -13 31
rect -4 19 4 27
rect 8 23 63 31
rect -52 10 -15 18
rect 55 11 63 15
rect 48 10 63 11
rect -23 7 63 10
rect 67 13 75 21
rect -35 2 -27 6
rect -23 2 53 7
rect 67 2 71 13
rect -47 -2 -27 2
rect 57 -2 71 2
rect -47 -6 -39 -2
rect -31 -6 65 -2
rect -47 -19 -13 -11
rect -4 -18 4 -10
rect 8 -19 65 -11
<< labels >>
rlabel space 28 -21 76 35 3 ^p
rlabel metal1 8 23 63 31 1 Vdd!|pin|s|1
rlabel metal1 -25 23 -13 31 1 GND!|pin|s|0
rlabel metal1 -47 -19 -13 -11 1 GND!|pin|s|1
rlabel metal1 8 -19 65 -11 1 Vdd!|pin|s|0
rlabel metal1 -4 -18 4 -10 1 a
rlabel metal1 -4 19 4 27 1 b
rlabel metal1 -23 2 53 10 1 x
rlabel metal1 -52 10 -15 18 1 x
rlabel metal1 55 24 63 32 1 Vdd!|pin|s|1
<< end >>
