// -----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Raghu P Gudla
// Created On   :  09/22/2018
// Description  :  SVT_BFM level Defines, Typedefs, or PARAMETERS.
// -----------------------------------------------------------------------------


//   `define SVT_AXI_USER_DEFINES_SVI

