magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -220 -724 -214 -723
rect -220 -730 -214 -726
rect -220 -736 -214 -732
rect -220 -742 -214 -738
rect -220 -748 -214 -744
rect -220 -754 -214 -750
rect -220 -757 -214 -756
rect -220 -761 -218 -757
rect -220 -762 -214 -761
rect -220 -768 -214 -764
rect -220 -774 -214 -770
rect -220 -780 -214 -776
rect -220 -786 -214 -782
rect -220 -792 -214 -788
rect -220 -795 -214 -794
<< pdiffusion >>
rect -195 -712 -187 -709
rect -199 -713 -187 -712
rect -199 -717 -187 -715
rect -199 -721 -193 -717
rect -199 -722 -187 -721
rect -199 -725 -187 -724
rect -189 -729 -187 -725
rect -199 -730 -187 -729
rect -199 -733 -187 -732
rect -199 -737 -193 -733
rect -199 -738 -187 -737
rect -199 -741 -187 -740
rect -189 -745 -187 -741
rect -199 -746 -187 -745
rect -199 -749 -187 -748
rect -199 -753 -193 -749
rect -199 -754 -187 -753
rect -199 -757 -187 -756
rect -189 -761 -187 -757
rect -199 -762 -187 -761
rect -199 -765 -187 -764
rect -199 -769 -193 -765
rect -199 -770 -187 -769
rect -199 -773 -187 -772
rect -189 -777 -187 -773
rect -199 -778 -187 -777
rect -199 -781 -187 -780
rect -199 -785 -193 -781
rect -199 -786 -187 -785
rect -199 -789 -187 -788
rect -189 -793 -187 -789
rect -199 -794 -187 -793
rect -199 -797 -187 -796
<< ntransistor >>
rect -220 -726 -214 -724
rect -220 -732 -214 -730
rect -220 -738 -214 -736
rect -220 -744 -214 -742
rect -220 -750 -214 -748
rect -220 -756 -214 -754
rect -220 -764 -214 -762
rect -220 -770 -214 -768
rect -220 -776 -214 -774
rect -220 -782 -214 -780
rect -220 -788 -214 -786
rect -220 -794 -214 -792
<< ptransistor >>
rect -199 -715 -187 -713
rect -199 -724 -187 -722
rect -199 -732 -187 -730
rect -199 -740 -187 -738
rect -199 -748 -187 -746
rect -199 -756 -187 -754
rect -199 -764 -187 -762
rect -199 -772 -187 -770
rect -199 -780 -187 -778
rect -199 -788 -187 -786
rect -199 -796 -187 -794
<< polysilicon >>
rect -202 -715 -199 -713
rect -187 -715 -184 -713
rect -203 -724 -199 -722
rect -187 -724 -184 -722
rect -223 -726 -220 -724
rect -214 -726 -211 -724
rect -203 -730 -201 -724
rect -223 -732 -220 -730
rect -214 -732 -199 -730
rect -187 -732 -184 -730
rect -223 -738 -220 -736
rect -214 -738 -211 -736
rect -208 -740 -199 -738
rect -187 -740 -184 -738
rect -208 -742 -206 -740
rect -223 -744 -220 -742
rect -214 -744 -206 -742
rect -203 -748 -199 -746
rect -187 -748 -184 -746
rect -223 -750 -220 -748
rect -214 -750 -201 -748
rect -203 -754 -201 -750
rect -223 -756 -220 -754
rect -214 -756 -211 -754
rect -203 -756 -199 -754
rect -187 -756 -184 -754
rect -223 -764 -220 -762
rect -214 -764 -211 -762
rect -203 -764 -199 -762
rect -187 -764 -184 -762
rect -203 -768 -201 -764
rect -223 -770 -220 -768
rect -214 -770 -201 -768
rect -203 -772 -199 -770
rect -187 -772 -184 -770
rect -223 -776 -220 -774
rect -214 -776 -206 -774
rect -208 -778 -206 -776
rect -208 -780 -199 -778
rect -187 -780 -184 -778
rect -223 -782 -220 -780
rect -214 -782 -211 -780
rect -223 -788 -220 -786
rect -214 -788 -199 -786
rect -187 -788 -184 -786
rect -223 -794 -220 -792
rect -214 -794 -211 -792
rect -203 -794 -201 -788
rect -203 -796 -199 -794
rect -187 -796 -184 -794
<< ndcontact >>
rect -220 -723 -214 -719
rect -218 -761 -214 -757
rect -220 -799 -214 -795
<< pdcontact >>
rect -199 -712 -195 -708
rect -193 -721 -187 -717
rect -199 -729 -189 -725
rect -193 -737 -187 -733
rect -199 -745 -189 -741
rect -193 -753 -187 -749
rect -199 -761 -189 -757
rect -193 -769 -187 -765
rect -199 -777 -189 -773
rect -193 -785 -187 -781
rect -199 -793 -189 -789
rect -199 -801 -187 -797
<< metal1 >>
rect -199 -712 -195 -708
rect -220 -723 -214 -719
rect -199 -725 -196 -712
rect -193 -721 -187 -717
rect -199 -729 -189 -725
rect -199 -741 -196 -729
rect -193 -737 -187 -733
rect -199 -745 -189 -741
rect -199 -757 -196 -745
rect -193 -753 -187 -749
rect -218 -761 -189 -757
rect -199 -773 -196 -761
rect -193 -769 -187 -765
rect -199 -777 -189 -773
rect -199 -789 -196 -777
rect -193 -785 -187 -781
rect -199 -793 -189 -789
rect -220 -799 -214 -795
rect -199 -801 -187 -797
<< labels >>
rlabel polysilicon -186 -723 -186 -723 3 e
rlabel polysilicon -186 -731 -186 -731 3 e
rlabel polysilicon -186 -739 -186 -739 3 c
rlabel polysilicon -186 -755 -186 -755 3 b
rlabel polysilicon -186 -747 -186 -747 3 b
rlabel polysilicon -186 -771 -186 -771 3 d
rlabel polysilicon -186 -763 -186 -763 3 d
rlabel polysilicon -186 -779 -186 -779 3 c
rlabel polysilicon -186 -795 -186 -795 3 a
rlabel polysilicon -186 -787 -186 -787 3 a
rlabel space -191 -802 -184 -718 3 ^p
rlabel polysilicon -221 -793 -221 -793 3 _SReset!
rlabel polysilicon -221 -725 -221 -725 3 _SReset!
rlabel polysilicon -221 -787 -221 -787 3 a
rlabel polysilicon -221 -781 -221 -781 3 b
rlabel polysilicon -221 -775 -221 -775 3 c
rlabel polysilicon -221 -769 -221 -769 3 d
rlabel polysilicon -221 -763 -221 -763 3 e
rlabel polysilicon -221 -755 -221 -755 3 a
rlabel polysilicon -221 -749 -221 -749 3 b
rlabel polysilicon -221 -743 -221 -743 3 c
rlabel polysilicon -221 -737 -221 -737 3 d
rlabel polysilicon -221 -731 -221 -731 3 e
rlabel space -223 -800 -217 -718 7 ^n
rlabel polysilicon -186 -714 -186 -714 1 _PReset!
rlabel pdcontact -197 -791 -197 -791 1 x
rlabel pdcontact -197 -775 -197 -775 1 x
rlabel pdcontact -197 -759 -197 -759 1 x
rlabel pdcontact -197 -743 -197 -743 1 x
rlabel pdcontact -197 -727 -197 -727 1 x
rlabel pdcontact -190 -719 -190 -719 1 Vdd!
rlabel pdcontact -190 -735 -190 -735 1 Vdd!
rlabel pdcontact -190 -751 -190 -751 1 Vdd!
rlabel pdcontact -190 -767 -190 -767 1 Vdd!
rlabel pdcontact -190 -783 -190 -783 1 Vdd!
rlabel pdcontact -190 -799 -190 -799 1 Vdd!
rlabel ndcontact -216 -759 -216 -759 1 x
rlabel ndcontact -217 -797 -217 -797 1 GND!
rlabel ndcontact -217 -721 -217 -721 5 GND!
rlabel pdcontact -197 -710 -197 -710 1 x
<< end >>
