// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

`define pargpio 		 `soc.pargpio
`define pmu_wrapper1 		 `pargpio.pmu_wrapper1

