magic
tech scmos
timestamp 965070451
<< ndiffusion >>
rect 198 645 206 646
rect 198 637 206 642
rect 198 633 206 634
rect 198 624 206 625
rect 198 616 206 621
rect 198 612 206 613
rect 198 603 206 604
rect 198 595 206 600
rect 198 591 206 592
rect 198 582 206 583
rect 198 574 206 579
rect 198 570 206 571
<< pdiffusion >>
rect 222 655 230 656
rect 222 651 230 652
rect 222 642 230 643
rect 222 638 230 639
rect 222 629 230 630
rect 222 625 230 626
rect 222 616 230 617
rect 222 612 230 613
rect 222 603 230 604
rect 222 599 230 600
rect 222 590 230 591
rect 222 586 230 587
rect 222 577 230 578
rect 222 573 230 574
rect 222 564 230 565
rect 222 560 230 561
<< ntransistor >>
rect 198 642 206 645
rect 198 634 206 637
rect 198 621 206 624
rect 198 613 206 616
rect 198 600 206 603
rect 198 592 206 595
rect 198 579 206 582
rect 198 571 206 574
<< ptransistor >>
rect 222 652 230 655
rect 222 639 230 642
rect 222 626 230 629
rect 222 613 230 616
rect 222 600 230 603
rect 222 587 230 590
rect 222 574 230 577
rect 222 561 230 564
<< polysilicon >>
rect 208 652 222 655
rect 230 652 234 655
rect 208 645 211 652
rect 194 642 198 645
rect 206 642 211 645
rect 217 639 222 642
rect 230 639 234 642
rect 217 637 220 639
rect 194 634 198 637
rect 206 634 220 637
rect 217 626 222 629
rect 230 626 234 629
rect 217 624 220 626
rect 194 621 198 624
rect 206 621 220 624
rect 194 613 198 616
rect 206 613 222 616
rect 230 613 234 616
rect 194 600 198 603
rect 206 600 222 603
rect 230 600 234 603
rect 194 592 198 595
rect 206 592 220 595
rect 217 590 220 592
rect 217 587 222 590
rect 230 587 234 590
rect 194 579 198 582
rect 206 579 220 582
rect 217 577 220 579
rect 217 574 222 577
rect 230 574 234 577
rect 194 571 198 574
rect 206 571 211 574
rect 208 564 211 571
rect 208 561 222 564
rect 230 561 234 564
<< ndcontact >>
rect 198 646 206 654
rect 198 625 206 633
rect 198 604 206 612
rect 198 583 206 591
rect 198 562 206 570
<< pdcontact >>
rect 222 656 230 664
rect 222 643 230 651
rect 222 630 230 638
rect 222 617 230 625
rect 222 604 230 612
rect 222 591 230 599
rect 222 578 230 586
rect 222 565 230 573
rect 222 552 230 560
<< polycontact >>
rect 234 647 242 655
rect 186 629 194 637
rect 234 621 242 629
rect 186 608 194 616
rect 234 600 242 608
rect 186 587 194 595
rect 234 574 242 582
rect 186 566 194 574
<< metal1 >>
rect 222 656 230 664
rect 198 646 206 654
rect 210 643 230 651
rect 234 647 242 655
rect 186 629 194 637
rect 210 633 218 643
rect 187 616 192 629
rect 198 625 218 633
rect 222 630 230 638
rect 235 629 240 647
rect 210 617 230 625
rect 234 621 242 629
rect 186 608 194 616
rect 187 595 192 608
rect 198 604 206 612
rect 210 599 218 617
rect 222 604 230 612
rect 235 608 240 621
rect 234 600 242 608
rect 186 587 194 595
rect 210 591 230 599
rect 187 574 192 587
rect 198 583 218 591
rect 186 566 194 574
rect 210 573 218 583
rect 222 578 230 586
rect 235 582 240 600
rect 234 574 242 582
rect 198 562 206 570
rect 210 565 230 573
rect 222 552 230 560
<< labels >>
rlabel metal1 226 595 226 595 1 x
rlabel metal1 226 608 226 608 5 Vdd!
rlabel metal1 226 582 226 582 1 Vdd!
rlabel polysilicon 231 601 231 601 1 b
rlabel metal1 226 556 226 556 1 Vdd!
rlabel polysilicon 231 575 231 575 1 b
rlabel metal1 226 647 226 647 1 x
rlabel metal1 226 660 226 660 5 Vdd!
rlabel metal1 226 634 226 634 1 Vdd!
rlabel polysilicon 231 653 231 653 1 b
rlabel metal1 226 621 226 621 5 x
rlabel polysilicon 231 627 231 627 1 b
rlabel metal1 202 608 202 608 5 GND!
rlabel polysilicon 197 593 197 593 3 a
rlabel polysilicon 197 572 197 572 3 a
rlabel metal1 202 587 202 587 5 x
rlabel metal1 202 566 202 566 1 GND!
rlabel polysilicon 197 614 197 614 3 a
rlabel polysilicon 197 635 197 635 3 a
rlabel metal1 202 650 202 650 5 GND!
rlabel metal1 202 629 202 629 5 x
rlabel metal1 226 569 226 569 5 x
rlabel space 185 561 199 655 7 ^n
rlabel space 229 551 243 665 3 ^p
rlabel polysilicon 231 562 231 562 1 a
rlabel polysilicon 231 588 231 588 1 a
rlabel polysilicon 231 614 231 614 1 a
rlabel polysilicon 231 640 231 640 1 a
rlabel polysilicon 197 643 197 643 3 b
rlabel polysilicon 197 622 197 622 3 b
rlabel polysilicon 197 601 197 601 3 b
rlabel polysilicon 197 580 197 580 3 b
<< end >>
