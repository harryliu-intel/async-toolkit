//There will be a TB here
