magic
tech scmos
timestamp 970024428
<< ndiffusion >>
rect -24 564 -8 565
rect -24 556 -8 561
rect -24 552 -8 553
<< pdiffusion >>
rect 8 564 24 565
rect 8 560 24 561
rect 8 551 24 552
rect 8 547 24 548
<< ntransistor >>
rect -24 561 -8 564
rect -24 553 -8 556
<< ptransistor >>
rect 8 561 24 564
rect 8 548 24 551
<< polysilicon >>
rect -28 561 -24 564
rect -8 561 -4 564
rect 4 561 8 564
rect 24 561 28 564
rect -28 553 -24 556
rect -8 553 -1 556
rect -4 551 -1 553
rect -4 548 8 551
rect 24 548 28 551
<< ndcontact >>
rect -24 565 -8 573
rect -24 544 -8 552
<< pdcontact >>
rect 8 565 24 573
rect 8 552 24 560
rect 8 539 24 547
<< psubstratepcontact >>
rect -41 557 -33 565
<< nsubstratencontact >>
rect 33 557 41 565
<< polycontact >>
rect -4 561 4 569
rect -4 540 4 548
<< metal1 >>
rect -21 573 -8 575
rect -41 565 -8 573
rect 8 573 21 575
rect -41 557 -33 565
rect 8 565 41 573
rect -4 561 4 563
rect 8 557 24 560
rect 33 557 41 565
rect -24 551 -21 552
rect 21 552 24 557
rect -24 544 -8 551
rect -4 545 4 548
rect 8 545 24 547
rect 8 539 9 545
rect 21 539 24 545
<< m2contact >>
rect -21 575 -3 581
rect 3 575 21 581
rect -4 563 4 569
rect -21 551 -8 557
rect 8 551 21 557
rect -4 539 4 545
rect 9 539 21 545
<< metal2 >>
rect -6 563 6 569
rect -21 551 21 557
rect -27 539 4 545
<< m3contact >>
rect -21 575 -3 581
rect 3 575 21 581
rect 9 539 21 545
<< metal3 >>
rect -21 536 -3 584
rect 3 536 21 584
<< labels >>
rlabel metal1 12 569 12 569 5 Vdd!
rlabel m2contact 12 543 12 543 1 Vdd!
rlabel polysilicon 25 562 25 562 1 b
rlabel polysilicon 25 549 25 549 1 a
rlabel metal1 -12 569 -12 569 5 GND!
rlabel polysilicon -25 562 -25 562 3 b
rlabel polysilicon -25 554 -25 554 3 a
rlabel metal2 0 566 0 566 1 b
rlabel metal2 -27 539 -25 545 3 ^n
rlabel metal2 -26 542 -26 542 3 a
rlabel metal2 0 551 0 557 1 x
rlabel metal1 -37 561 -37 561 3 GND!
rlabel space -42 538 -23 574 7 ^n
rlabel metal1 37 561 37 561 7 Vdd!
rlabel space 23 538 42 574 3 ^p
<< end >>
