// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

`define CCU_TOP soc.parcgu.ccu_top
`define CGU soc.parcgu.cgu
`define CLTAP_WRAPPER_DFT soc.pargpio.cltap_wrapper_dft
`define DFXAGG_TOP soc.pargpio.dfxagg_top
`define EC_TOP soc.parmain.ec_top
`define FUSE_HIP soc.parfuse.fuse_hip
`define FUSE_TOP soc.parfuse.fuse_top
`define GPCOMGPIOCOM0UNIT_WRAPPER soc.pargpio.gpcomgpiocom0unit_wrapper
`define GPIOHIP_STUB soc.pargpio.gpiohip_stub
`define MPHY_0 soc.parpcie.mphy_0
`define NORTHPEAK soc.parmain.northpeak
`define P2SB soc.parmain.p2sb
`define PMSRVR_UPMAS soc.pargpio.pmsrvr_upmas
`define PMU_WRAPPER1 soc.pargpio.pmu_wrapper1
`define PSF0 soc.parmain.psf0
`define PSF1 soc.parmain.psf1
`define SBR_GP0 soc.parmain.sbr_gp0
`define SBR_GP1 soc.parmain.sbr_gp1
`define SBR_GP2 soc.parmain.sbr_gp2
`define SBR_PM0 soc.parmain.sbr_pm0
`define SBR_PM1 soc.parmain.sbr_pm1
`define SIP_IOSF_TAM_TOP_WRAPPER1 soc.parmain.sip_iosf_tam_top_wrapper1
`define TAP2IOSFSB_0 soc.pargpio.tap2iosfsb_0
`define TAP2IOSFSB_1 soc.parmain.tap2iosfsb_1
`define TAPLINK_0_WRAPPER soc.pargpio.taplink_0_wrapper
`define TSANADIGLDO_0 soc.parmain.tsanadigldo_0
`define TSANADIGLDO_1 soc.parmain.tsanadigldo_1
`define TSANADIGLDO_2 soc.parmain.tsanadigldo_2
`define TSANADIGLDO_3 soc.parmain.tsanadigldo_3
`define USP_0_PIPELINE soc.parchannel.usp_0_pipeline
`define USP_1_PIPELINE soc.parchannel.usp_1_pipeline
`define USP_LL soc.parpcie.usp_ll
`define USP_MM soc.parpcie.usp_mm
`define USP_TT soc.parpcie.usp_tt
`define VSP0_TT soc.parmain.vsp0_tt
`define VSP1_TT soc.parmain.vsp1_tt
`define VSP2_TT soc.parmain.vsp2_tt
`define VSP3_TT soc.parmain.vsp3_tt
