//-----------------------------------------------------------------------------
// Title         : Ingress sequence library
// Project       : Madison Bay
//-----------------------------------------------------------------------------
// File          : ingress_seqlib.sv
// Author        : jose.j.godinez.carrillo  <jjgodine@ichips.intel.com>
// Created       : 21.08.2018
// Last modified : 21.08.2018
//-----------------------------------------------------------------------------
// Description :
//
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by Intel Corporation This model is the confidential and
// proprietary property of Intel Corporation and the possession or use of this
// file requires a written license from Intel Corporation.
//------------------------------------------------------------------------------
// Modification history :
// 21.08.2018 : created
//-----------------------------------------------------------------------------

`include "mby_igr_env_base_seq.sv"
`include "mby_igr_extended_base_seq.sv"
`include "mby_igr_hard_reset_seq.sv"
