magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -83 304 -79 305
rect -83 298 -79 302
rect -83 295 -79 296
<< pdiffusion >>
rect -67 304 -63 305
rect -67 298 -63 302
rect -67 295 -63 296
<< ntransistor >>
rect -83 302 -79 304
rect -83 296 -79 298
<< ptransistor >>
rect -67 302 -63 304
rect -67 296 -63 298
<< polysilicon >>
rect -86 302 -83 304
rect -79 302 -67 304
rect -63 302 -60 304
rect -86 296 -83 298
rect -79 296 -67 298
rect -63 296 -60 298
<< ndcontact >>
rect -83 305 -79 309
rect -83 291 -79 295
<< pdcontact >>
rect -67 305 -63 309
rect -67 291 -63 295
<< metal1 >>
rect -83 305 -63 309
rect -83 291 -79 295
rect -67 291 -63 295
<< labels >>
rlabel polysilicon -84 297 -84 297 3 a
rlabel polysilicon -84 303 -84 303 3 b
rlabel space -87 290 -83 310 7 ^n
rlabel space -63 290 -59 310 3 ^p
rlabel polysilicon -62 297 -62 297 3 a
rlabel polysilicon -62 303 -62 303 3 b
rlabel ndcontact -81 307 -81 307 1 x
rlabel ndcontact -81 293 -81 293 1 GND!
rlabel pdcontact -65 307 -65 307 1 x
rlabel pdcontact -65 293 -65 293 1 Vdd!
<< end >>
