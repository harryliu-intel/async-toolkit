///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
// ---------------------------------------------------------------------------------------------------------------------
// -- Author : Jim McCormick <jim.mccormick@intel.com>
// -- Project Name : ??? 
// -- Description  : The top-level-module in this tesbench 
//
// -- Instantiation Hierarchy:                                  definition file
//                                                              ---------------
//          module  top                                         top.sv
//              msh_dut_if dut_if                               msh_dut_if.sv
//              msh_node    dut                                 $(CLONE_ROOT)/src/msh/rtl/mby_msh_node.sv
//                  ...                                         (see mby_msh.sv)
//              testcase    test                                tests/<testcase>.sv
//                  env     env                                 env.sv
//                      system_driver   sys_drvr                system_driver.sv
//                      configuration   cfg                     configuration.sv
//                      id_generator    id_gen                  ig_generator.sv
//                      inp_driver      inp_driver              inp_driver.sv
//                          stimulus        stim                stimulus.sv
//                      monitor         mntr                    monitor.sv
//                      scoreboard      sb                      scoreboard.sv
//                  `include "test_loop_include"                test_loop_include.sv
//
//  FIXME:  change these to mesh assertions
//          bind tmpl_arb                                       $(CLONE_ROOT)/src/rtl/template/sva/template_binds.svh
//              tmpl_arb_assert a__tmpl_arb_assert              $(CLONE_ROOT)/src/rtl/template/sva/tmpl_arb_asert.sv
//
//  note:  verilog/msh_sim_pkg.sv is included on the compilation command line so that it can be used widely
//         without being included everywhere.
// ---------------------------------------------------------------------------------------------------------------------

// A module is a top-level-module if is defined but never instantiated

module top 
import mby_msh_pkg::*;
import msh_sim_pkg::*;
();

    logic clk = 0;                              // declare clock


    // define clock
    initial                                     // "initial" procedures are executed at the beginning of simulation
        forever                                 // "forever" is just a type of loop that executes forever 
            #(10/2)                             //  #<n> means wait <n> clocks
                clk = ~clk;                     //  invert the clock

    // instantiate DUT interface
    msh_dut_if #(
        .NUM_MSH_ROWS(NUM_MSH_ROWS),
        .NUM_MSH_COLS(NUM_MSH_COLS)
    ) dut_if (
        .mclk(clk)                               // pass clock into this interface to make it part of the interface
    );

logic reset;

    // start firing reset immediately to protect reset guarded assertions
    initial dut_if.chreset = 1'b1;
    initial dut_if.csreset = 1'b1;
    initial dut_if.mhreset = 1'b1;
    initial dut_if.msreset = 1'b1;
    initial reset = 1'b1;

    // instantiate DUT (Design Under Test)
//    mby_msh dut (
//
//        // DUT inputs
//        .mclk       (dut_if.mclk          ),      // The interface instantiated above is connected to the DUT 
//        .i_reset    (dut_if.i_reset       )      // Note the naming convention i_<???> for inputs.
//       
//    );

mby_msh #(

    .NUM_MSH_ROWS(NUM_MSH_ROWS),
    .NUM_MSH_COLS(NUM_MSH_COLS)

) msh (

    
    .cclk(clk),                                // core clock
    .chreset(dut_if.chreset),                  // core hard reset
    .csreset(dut_if.csreset),                  // core soft reset

    .mclk(clk),                                // mesh clock
    .mhreset(dut_if.mhreset),                  // mesh hard reset
    .msreset(dut_if.msreset),                  // mesh soft reset


     .i_igr_eb_wreq_valid   (dut_if.i_igr_eb_wreq_valid),
     .i_igr_eb_wr_seg_ptr   (dut_if.i_igr_eb_wr_seg_ptr),
     .i_igr_eb_wr_sema      (dut_if.i_igr_eb_wr_sema),
     .i_igr_eb_wr_wd_sel    (dut_if.i_igr_eb_wr_wd_sel),
     .i_igr_eb_wreq_id      (dut_if.i_igr_eb_wreq_id),
     .i_igr_eb_wr_data      (dut_if.i_igr_eb_wr_data),
     .o_igr_wb_wreq_credits (dut_if.o_igr_wb_wreq_credits),
     .i_igr_wb_wreq_valid   (dut_if.i_igr_wb_wreq_valid),
     .i_igr_wb_wr_seg_ptr   (dut_if.i_igr_wb_wr_seg_ptr),
     .i_igr_wb_wr_sema      (dut_if.i_igr_wb_wr_sema),
     .i_igr_wb_wr_wd_sel    (dut_if.i_igr_wb_wr_wd_sel),
     .i_igr_wb_wreq_id      (dut_if.i_igr_wb_wreq_id),
     .i_igr_wb_wr_data      (dut_if.i_igr_wb_wr_data),
     .o_igr_eb_wreq_credits (dut_if.o_igr_eb_wreq_credits),
     .i_egr_eb_rreq_valid   (dut_if.i_egr_eb_rreq_valid),
     .i_egr_eb_seg_ptr      (dut_if.i_egr_eb_seg_ptr),
     .i_egr_eb_sema         (dut_if.i_egr_eb_sema),
     .i_egr_eb_wd_sel       (dut_if.i_egr_eb_wd_sel),
     .i_egr_eb_req_id       (dut_if.i_egr_eb_req_id),
     .o_egr_wb_rreq_credits (dut_if.o_egr_wb_rreq_credits),
     .i_egr_wb_rreq_valid   (dut_if.i_egr_wb_rreq_valid),
     .i_egr_wb_seg_ptr      (dut_if.i_egr_wb_seg_ptr),
     .i_egr_wb_sema         (dut_if.i_egr_wb_sema),
     .i_egr_wb_wd_sel       (dut_if.i_egr_wb_wd_sel),
     .i_egr_wb_req_id       (dut_if.i_egr_wb_req_id),
     .o_egr_eb_rreq_credits (dut_if.o_egr_eb_rreq_credits),
     .o_egr_wb_rrsp_valid   (dut_if.o_egr_wb_rrsp_valid),
     .o_egr_wb_rrsp_dest_block  (dut_if.o_egr_wb_rrsp_dest_block),
     .o_egr_wb_rrsp_req_id  (dut_if.o_egr_wb_rrsp_req_id),
     .o_egr_wb_rd_data      (dut_if.o_egr_wb_rd_data),
     .o_egr_eb_rrsp_valid   (dut_if.o_egr_eb_rrsp_valid),
     .o_egr_eb_rrsp_dest_block  (dut_if.o_egr_eb_rrsp_dest_block),
     .o_egr_eb_rrsp_req_id  (dut_if.o_egr_eb_rrsp_req_id),
     .o_egr_eb_rd_data      (dut_if.o_egr_eb_rd_data),
     .i_sb_wreq_valid       (dut_if.i_sb_wreq_valid),
     .i_sb_wr_seg_ptr       (dut_if.i_sb_wr_seg_ptr),
     .i_sb_wr_sema          (dut_if.i_sb_wr_sema),
     .i_sb_wr_wd_sel        (dut_if.i_sb_wr_wd_sel),
     .i_sb_wreq_id          (dut_if.i_sb_wreq_id),
     .i_sb_wr_data          (dut_if.i_sb_wr_data),
     .o_nb_wreq_credits     (dut_if.o_nb_wreq_credits),
     .i_nb_wreq_valid       (dut_if.i_nb_wreq_valid),
     .i_nb_wr_seg_ptr       (dut_if.i_nb_wr_seg_ptr),
     .i_nb_wr_sema          (dut_if.i_nb_wr_sema),
     .i_nb_wr_wd_sel        (dut_if.i_nb_wr_wd_sel),
     .i_nb_wreq_id          (dut_if.i_nb_wreq_id),
     .i_nb_wr_data          (dut_if.i_nb_wr_data),
     .o_sb_wreq_credits     (dut_if.o_sb_wreq_credits),
     .i_sb_rreq_valid       (dut_if.i_sb_rreq_valid),
     .i_sb_rreq_seg_ptr     (dut_if.i_sb_rreq_seg_ptr),
     .i_sb_rreq_sema        (dut_if.i_sb_rreq_sema),
     .i_sb_rreq_wd_sel      (dut_if.i_sb_rreq_wd_sel),
     .i_sb_rreq_id          (dut_if.i_sb_rreq_id),
     .o_nb_rreq_credits     (dut_if.o_nb_rreq_credits),
     .i_nb_rreq_valid       (dut_if.i_nb_rreq_valid),
     .i_nb_rreq_seg_ptr     (dut_if.i_nb_rreq_seg_ptr),
     .i_nb_rreq_sema        (dut_if.i_nb_rreq_sema),
     .i_nb_rreq_wd_sel      (dut_if.i_nb_rreq_wd_sel),
     .i_nb_rreq_id          (dut_if.i_nb_rreq_id),
     .o_sb_rreq_credits     (dut_if.o_sb_rreq_credits),
     .o_nb_rrsp_valid       (dut_if.o_nb_rrsp_valid),
     .o_nb_rrsp_dest_block  (dut_if.o_nb_rrsp_dest_block),
     .o_nb_rrsp_req_id      (dut_if.o_nb_rrsp_req_id),
     .o_nb_rd_data          (dut_if.o_nb_rd_data),
     .o_sb_rrsp_valid       (dut_if.o_sb_rrsp_valid),
     .o_sb_rrsp_dest_block  (dut_if.o_sb_rrsp_dest_block),
     .o_sb_rrsp_req_id      (dut_if.o_sb_rrsp_req_id),
     .o_sb_rd_data          (dut_if.o_sb_rd_data)
    
);

    // instantiate testcase
    testcase test(
        dut_if                                    // pass interface dut_if into testcase
    );

endmodule

