magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 127 76 130 78
rect 143 76 144 80
rect 143 75 149 76
rect 127 68 130 72
rect 143 72 149 73
rect 143 67 149 68
rect 127 64 130 66
rect 143 64 149 65
<< pdiffusion >>
rect 107 77 115 78
rect 94 73 98 74
rect 107 74 115 75
rect 94 67 98 71
rect 111 71 115 74
rect 161 75 165 76
rect 107 68 110 70
rect 94 64 98 65
rect 107 64 110 66
rect 161 72 165 73
rect 161 67 165 68
rect 161 64 165 65
<< ntransistor >>
rect 127 72 130 76
rect 143 73 149 75
rect 127 66 130 68
rect 143 65 149 67
<< ptransistor >>
rect 107 75 115 77
rect 94 71 98 73
rect 161 73 165 75
rect 94 65 98 67
rect 107 66 110 68
rect 161 65 165 67
<< polysilicon >>
rect 104 75 107 77
rect 115 76 124 77
rect 115 75 127 76
rect 122 74 127 75
rect 91 71 94 73
rect 98 71 101 73
rect 124 72 127 74
rect 130 72 133 76
rect 139 73 143 75
rect 149 73 161 75
rect 165 73 169 75
rect 91 65 94 67
rect 98 65 101 67
rect 104 66 107 68
rect 110 66 116 68
rect 120 66 127 68
rect 130 66 133 68
rect 139 67 141 73
rect 167 67 169 73
rect 139 65 143 67
rect 149 65 161 67
rect 165 65 169 67
<< ndcontact >>
rect 127 78 131 82
rect 144 76 149 80
rect 143 68 149 72
rect 127 60 131 64
rect 143 60 149 64
<< pdcontact >>
rect 107 78 115 82
rect 94 74 98 78
rect 107 70 111 74
rect 161 76 165 80
rect 94 60 98 64
rect 161 68 165 72
rect 107 60 111 64
rect 161 60 165 64
<< polycontact >>
rect 137 75 141 79
rect 116 65 120 69
<< metal1 >>
rect 107 78 115 82
rect 127 81 131 82
rect 127 79 140 81
rect 127 78 141 79
rect 94 74 98 78
rect 137 75 141 78
rect 144 76 149 80
rect 161 76 165 80
rect 95 73 98 74
rect 107 73 111 74
rect 95 70 111 73
rect 143 71 165 72
rect 117 69 165 71
rect 116 68 165 69
rect 116 65 120 68
rect 94 60 111 64
rect 127 60 149 64
rect 161 60 165 64
<< labels >>
rlabel polysilicon 93 66 93 66 3 a
rlabel polysilicon 93 72 93 72 3 b
rlabel space 91 59 95 79 7 ^p1
rlabel polysilicon 116 76 116 76 5 _PReset!
rlabel space 164 59 169 81 3 ^p2
rlabel space 148 58 170 82 3 ^n2
rlabel ndcontact 129 62 129 62 1 GND!
rlabel ndcontact 129 80 129 80 5 _x
rlabel pdcontact 96 62 96 62 1 Vdd!
rlabel pdcontact 96 76 96 76 1 _x
rlabel pdcontact 111 80 111 80 1 Vdd!
rlabel pdcontact 109 72 109 72 5 _x
rlabel pdcontact 109 62 109 62 1 Vdd!
rlabel ndcontact 147 62 147 62 1 GND!
rlabel ndcontact 147 78 147 78 5 GND!
rlabel pdcontact 163 70 163 70 1 x
rlabel ndcontact 147 70 147 70 1 x
rlabel pdcontact 163 78 163 78 5 Vdd!
rlabel pdcontact 163 62 163 62 1 Vdd!
<< end >>
