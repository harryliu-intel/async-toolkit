// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

//-----------------------------------------------------------------------------
// Title         : Ingress Testbench Config Object
// Project       : Madison Bay
//-----------------------------------------------------------------------------
// File          : mby_egr_tb_cfg.svh
// Author        : paul.j.pladsen <paul.j.pladsen@intel.com>
// Created       : 22.10.2018
// Last modified : 22.10.2018
//-----------------------------------------------------------------------------
// Description :
// This is the testbench configuration object which contains an instance of the dut configuration object and the env
// configuration object.  The dut configuration object holds all variable necessary to configure the design.  The env
// configuration object holds all variables and switches necessary to configure the simulation environment including
// BFMs, scoreboards, and test command line arguments.
//
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by Intel Corporation This model is the confidential and
// proprietary property of Intel Corporation and the possession or use of this
// file requires a written license from Intel Corporation.
//-----------------------------------------------------------------------------
// Modification history :
// 22.10.2018 : created
//-----------------------------------------------------------------------------

//-----------------------------------------------------------------------------
// Class: mby_egr_tb_cfg
//-----------------------------------------------------------------------------
class mby_egr_tb_cfg extends shdv_base_config;

   mby_egr_env_cfg env_cfg;
   mby_egr_dut_cfg dut_cfg;
   rand mesh_status_e mesh_status = NO_CONGESTION;
   rand eth_bfm_pkg::speed_e speed_cfg[4]; 
   bit randomize_speed_cfg = $test$plusargs("RAND_SPEED_CFG"); 
       
   constraint allowed_cfg{
      if(randomize_speed_cfg) 
         foreach(speed_cfg[i]) (i==0) ? speed_cfg[i] inside {eth_bfm_pkg::SPEED_400G,eth_bfm_pkg::SPEED_200G,eth_bfm_pkg::SPEED_100G} : speed_cfg[i] == eth_bfm_pkg::SPEED_OFF;
      else 
         foreach(speed_cfg[i]) (i==0) ? speed_cfg[i] inside {eth_bfm_pkg::SPEED_400G} : speed_cfg[i] == eth_bfm_pkg::SPEED_OFF;
   } 

   constraint mesh_status_c{
      (mesh_status == NO_CONGESTION)      -> (env_cfg.smm_bfm_cfg.delay_profile == IDEAL_DELAY);
      (mesh_status == MEDIUM_CONGESTION)  -> (env_cfg.smm_bfm_cfg.delay_profile == MEDIUM_DELAY);
      (mesh_status == HIGH_CONGESTION)    -> (env_cfg.smm_bfm_cfg.delay_profile == HIGH_DELAY);
      solve mesh_status before env_cfg.smm_bfm_cfg.delay_profile;
   }


   `uvm_object_utils_begin(mby_egr_tb_cfg)
      `uvm_field_object( env_cfg, UVM_ALL_ON )
      `uvm_field_object( dut_cfg, UVM_ALL_ON )
   `uvm_object_utils_end

   //--------------------------------------------------------------------------
   // Function: new
   //--------------------------------------------------------------------------
   function new (string name = "mby_egr_tb_cfg");
      super.new(name);
      
      env_cfg = new();
      dut_cfg = new();
   endfunction : new

endclass : mby_egr_tb_cfg
