module gmm_top(
    input   cclk,       // system clock
    input   arst,       // Asynchronous reset
    gmm_if.gmm    gmm_intf
);
 

endmodule
