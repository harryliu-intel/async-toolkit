magic
tech scmos
timestamp 965071540
<< ndiffusion >>
rect -214 -706 -206 -705
rect -214 -714 -206 -709
rect -214 -722 -206 -717
rect -214 -730 -206 -725
rect -214 -734 -206 -733
rect -214 -743 -206 -742
rect -214 -751 -206 -746
rect -214 -759 -206 -754
rect -214 -767 -206 -762
rect -214 -771 -206 -770
<< pdiffusion >>
rect -184 -691 -176 -690
rect -184 -695 -176 -694
rect -184 -704 -176 -703
rect -184 -708 -176 -707
rect -184 -717 -176 -716
rect -184 -721 -176 -720
rect -184 -730 -176 -729
rect -184 -734 -176 -733
rect -184 -743 -176 -742
rect -184 -747 -176 -746
rect -184 -756 -176 -755
rect -184 -760 -176 -759
rect -184 -769 -176 -768
rect -184 -773 -176 -772
rect -184 -782 -176 -781
rect -184 -786 -176 -785
<< ntransistor >>
rect -214 -709 -206 -706
rect -214 -717 -206 -714
rect -214 -725 -206 -722
rect -214 -733 -206 -730
rect -214 -746 -206 -743
rect -214 -754 -206 -751
rect -214 -762 -206 -759
rect -214 -770 -206 -767
<< ptransistor >>
rect -184 -694 -176 -691
rect -184 -707 -176 -704
rect -184 -720 -176 -717
rect -184 -733 -176 -730
rect -184 -746 -176 -743
rect -184 -759 -176 -756
rect -184 -772 -176 -769
rect -184 -785 -176 -782
<< polysilicon >>
rect -189 -694 -184 -691
rect -176 -694 -172 -691
rect -189 -704 -186 -694
rect -189 -706 -184 -704
rect -218 -709 -214 -706
rect -206 -707 -184 -706
rect -176 -707 -172 -704
rect -206 -709 -186 -707
rect -218 -717 -214 -714
rect -206 -717 -186 -714
rect -189 -720 -184 -717
rect -176 -720 -172 -717
rect -218 -725 -214 -722
rect -206 -725 -194 -722
rect -197 -730 -194 -725
rect -218 -733 -214 -730
rect -206 -733 -202 -730
rect -197 -733 -184 -730
rect -176 -733 -172 -730
rect -218 -746 -214 -743
rect -206 -746 -202 -743
rect -197 -746 -184 -743
rect -176 -746 -172 -743
rect -197 -751 -194 -746
rect -218 -754 -214 -751
rect -206 -754 -194 -751
rect -189 -759 -184 -756
rect -176 -759 -172 -756
rect -218 -762 -214 -759
rect -206 -762 -186 -759
rect -218 -770 -214 -767
rect -206 -769 -186 -767
rect -206 -770 -184 -769
rect -189 -772 -184 -770
rect -176 -772 -172 -769
rect -189 -782 -186 -772
rect -189 -785 -184 -782
rect -176 -785 -172 -782
<< ndcontact >>
rect -214 -705 -206 -697
rect -214 -742 -206 -734
rect -214 -779 -206 -771
<< pdcontact >>
rect -184 -690 -176 -682
rect -184 -703 -176 -695
rect -184 -716 -176 -708
rect -184 -729 -176 -721
rect -184 -742 -176 -734
rect -184 -755 -176 -747
rect -184 -768 -176 -760
rect -184 -781 -176 -773
rect -184 -794 -176 -786
<< metal1 >>
rect -184 -690 -176 -682
rect -214 -705 -206 -697
rect -196 -703 -176 -695
rect -196 -721 -188 -703
rect -184 -716 -176 -708
rect -196 -729 -176 -721
rect -196 -734 -188 -729
rect -214 -742 -188 -734
rect -184 -742 -176 -734
rect -196 -747 -188 -742
rect -196 -755 -176 -747
rect -214 -779 -206 -771
rect -196 -773 -188 -755
rect -184 -768 -176 -760
rect -196 -781 -176 -773
rect -184 -794 -176 -786
<< labels >>
rlabel metal1 -180 -724 -180 -724 1 x
rlabel metal1 -180 -790 -180 -790 1 Vdd!
rlabel metal1 -180 -699 -180 -699 5 x
rlabel polysilicon -175 -784 -175 -784 7 a
rlabel polysilicon -175 -693 -175 -693 7 d
rlabel metal1 -180 -712 -180 -712 5 Vdd!
rlabel metal1 -180 -738 -180 -738 5 Vdd!
rlabel metal1 -180 -764 -180 -764 1 Vdd!
rlabel metal1 -180 -777 -180 -777 1 x
rlabel metal1 -180 -751 -180 -751 5 x
rlabel metal1 -180 -686 -180 -686 1 Vdd!
rlabel polysilicon -175 -758 -175 -758 7 b
rlabel polysilicon -175 -706 -175 -706 7 d
rlabel polysilicon -175 -771 -175 -771 7 a
rlabel polysilicon -175 -745 -175 -745 7 c
rlabel polysilicon -175 -732 -175 -732 7 b
rlabel polysilicon -175 -719 -175 -719 7 c
rlabel space -176 -794 -171 -682 3 ^p
rlabel polysilicon -215 -732 -215 -732 3 a
rlabel polysilicon -215 -724 -215 -724 3 b
rlabel polysilicon -215 -716 -215 -716 3 c
rlabel metal1 -210 -738 -210 -738 5 x
rlabel metal1 -210 -701 -210 -701 5 GND!
rlabel metal1 -210 -775 -210 -775 1 GND!
rlabel polysilicon -215 -708 -215 -708 1 d
rlabel polysilicon -215 -761 -215 -761 3 b
rlabel polysilicon -215 -769 -215 -769 3 a
rlabel polysilicon -215 -753 -215 -753 1 c
rlabel space -219 -779 -214 -697 7 ^n
rlabel polysilicon -215 -745 -215 -745 3 d
<< end >>
