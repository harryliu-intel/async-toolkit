// File: mby_test_pack.sv

package mby_test_pack;
    
`ifdef XVM
   import ovm_pkg::*;
   import xvm_pkg::*;
   `include "ovm_macros.svh"
   `include "sla_macros.svh"
`endif

import sla_pkg::*;
    import uvm_pkg::*;
    import mby_env_pkg::*;
  
    `include "uvm_macros.svh"
    `include "slu_macros.svh"

    `include "mby_base_test.svh"
    `include "mby_alive_test/mby_alive_test.svh"
endpackage
