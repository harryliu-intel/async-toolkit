magic
tech scmos
timestamp 962519057
<< ndiffusion >>
rect -70 26 -66 27
rect -84 21 -80 24
rect -88 20 -80 21
rect -70 23 -66 24
rect -70 18 -66 19
rect -88 14 -80 18
rect -88 11 -80 12
rect -84 8 -80 11
rect -70 15 -66 16
rect -70 10 -66 11
rect -70 7 -66 8
rect -70 2 -66 3
rect -70 -1 -66 0
<< pdiffusion >>
rect -120 26 -114 27
rect -120 23 -114 24
rect -120 18 -114 19
rect -54 26 -50 27
rect -120 15 -114 16
rect -116 11 -114 15
rect -120 10 -114 11
rect -54 23 -50 24
rect -54 18 -50 19
rect -104 14 -100 15
rect -120 7 -114 8
rect -120 2 -114 3
rect -104 8 -100 12
rect -54 15 -50 16
rect -54 10 -50 11
rect -54 7 -50 8
rect -54 2 -50 3
rect -120 -1 -114 0
rect -54 -1 -50 0
<< ntransistor >>
rect -70 24 -66 26
rect -88 18 -80 20
rect -70 16 -66 18
rect -88 12 -80 14
rect -70 8 -66 10
rect -70 0 -66 2
<< ptransistor >>
rect -120 24 -114 26
rect -54 24 -50 26
rect -120 16 -114 18
rect -54 16 -50 18
rect -104 12 -100 14
rect -120 8 -114 10
rect -54 8 -50 10
rect -120 0 -114 2
rect -54 0 -50 2
<< polysilicon >>
rect -123 24 -120 26
rect -114 24 -110 26
rect -112 23 -110 24
rect -112 21 -90 23
rect -112 18 -110 21
rect -92 20 -90 21
rect -74 24 -70 26
rect -66 24 -54 26
rect -50 24 -46 26
rect -123 16 -120 18
rect -114 16 -110 18
rect -112 10 -110 16
rect -92 18 -88 20
rect -80 18 -77 20
rect -74 18 -72 24
rect -48 18 -46 24
rect -74 16 -70 18
rect -66 16 -54 18
rect -50 16 -46 18
rect -107 12 -104 14
rect -100 12 -95 14
rect -123 8 -120 10
rect -114 8 -110 10
rect -112 2 -110 8
rect -91 12 -88 14
rect -80 12 -77 14
rect -74 10 -72 16
rect -48 10 -46 16
rect -74 8 -70 10
rect -66 8 -54 10
rect -50 8 -46 10
rect -123 0 -120 2
rect -114 0 -110 2
rect -74 2 -72 8
rect -48 2 -46 8
rect -74 0 -70 2
rect -66 0 -54 2
rect -50 0 -46 2
<< ndcontact >>
rect -88 21 -84 25
rect -70 27 -66 31
rect -70 19 -66 23
rect -88 7 -84 11
rect -70 11 -66 15
rect -70 3 -66 7
rect -70 -5 -66 -1
<< pdcontact >>
rect -120 27 -114 31
rect -120 19 -114 23
rect -54 27 -50 31
rect -120 11 -116 15
rect -104 15 -100 19
rect -54 19 -50 23
rect -120 3 -114 7
rect -104 4 -100 8
rect -54 11 -50 15
rect -54 3 -50 7
rect -120 -5 -114 -1
rect -54 -5 -50 -1
<< polycontact >>
rect -78 24 -74 28
rect -95 10 -91 14
<< metal1 >>
rect -120 27 -114 31
rect -78 27 -74 28
rect -70 27 -66 31
rect -54 27 -50 31
rect -87 25 -74 27
rect -88 24 -74 25
rect -120 22 -114 23
rect -120 19 -110 22
rect -88 21 -84 24
rect -103 19 -85 21
rect -70 19 -50 23
rect -113 18 -85 19
rect -113 16 -100 18
rect -120 11 -116 15
rect -113 7 -110 16
rect -104 15 -100 16
rect -70 14 -66 15
rect -95 10 -91 14
rect -87 11 -66 14
rect -120 4 -110 7
rect -120 3 -114 4
rect -104 -1 -100 8
rect -94 4 -91 10
rect -88 7 -84 11
rect -62 7 -58 19
rect -54 11 -50 15
rect -70 6 -50 7
rect -78 4 -50 6
rect -94 3 -50 4
rect -94 1 -75 3
rect -120 -5 -100 -1
rect -70 -5 -66 -1
rect -54 -5 -50 -1
<< labels >>
rlabel polysilicon -79 19 -79 19 1 a
rlabel space -123 -6 -119 32 7 ^p1
rlabel polysilicon -121 17 -121 17 3 a
rlabel polysilicon -121 25 -121 25 3 a
rlabel polysilicon -121 9 -121 9 3 a
rlabel polysilicon -121 1 -121 1 3 a
rlabel space -51 -6 -46 32 3 ^p2
rlabel space -67 -7 -45 33 3 ^n2
rlabel polycontact -93 12 -93 12 1 x
rlabel pdcontact -102 17 -102 17 4 _x
rlabel pdcontact -102 6 -102 6 1 Vdd!
rlabel ndcontact -86 9 -86 9 1 GND!
rlabel ndcontact -86 23 -86 23 5 _x
rlabel pdcontact -118 29 -118 29 5 Vdd!
rlabel pdcontact -118 -3 -118 -3 1 Vdd!
rlabel pdcontact -118 13 -118 13 5 Vdd!
rlabel pdcontact -118 5 -118 5 1 _x
rlabel pdcontact -118 21 -118 21 5 _x
rlabel ndcontact -68 -3 -68 -3 1 GND!
rlabel ndcontact -68 13 -68 13 5 GND!
rlabel ndcontact -68 5 -68 5 1 x
rlabel ndcontact -68 21 -68 21 5 x
rlabel ndcontact -68 29 -68 29 5 GND!
rlabel pdcontact -52 29 -52 29 5 Vdd!
rlabel pdcontact -52 21 -52 21 5 x
rlabel pdcontact -52 13 -52 13 5 Vdd!
rlabel pdcontact -52 5 -52 5 1 x
rlabel pdcontact -52 -3 -52 -3 1 Vdd!
<< end >>
