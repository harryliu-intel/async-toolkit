// import files at global scope to resolve issues with collage generated content using package contents but not importing the packages
import mby_gmm_pkg::*;

