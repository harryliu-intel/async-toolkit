///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_modify_map_pkg.vh                                  
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_MODIFY_MAP_PKG_VH
`define MBY_PPE_MODIFY_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_modify_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_modify_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_modify_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_modify_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [23:0] CMD_1;  // RW
    logic [23:0] CMD_0;  // RW
} MOD_PROFILE_COMMAND_t;

localparam MOD_PROFILE_COMMAND_REG_STRIDE = 48'h8;
localparam MOD_PROFILE_COMMAND_REG_ENTRIES = 16;
localparam MOD_PROFILE_COMMAND_REGFILE_STRIDE = 48'h80;
localparam MOD_PROFILE_COMMAND_REGFILE_ENTRIES = 64;
localparam MOD_PROFILE_COMMAND_CR_ADDR = 48'h0;
localparam MOD_PROFILE_COMMAND_SIZE = 64;
localparam MOD_PROFILE_COMMAND_CMD_1_LO = 24;
localparam MOD_PROFILE_COMMAND_CMD_1_HI = 47;
localparam MOD_PROFILE_COMMAND_CMD_1_RESET = 24'h0;
localparam MOD_PROFILE_COMMAND_CMD_0_LO = 0;
localparam MOD_PROFILE_COMMAND_CMD_0_HI = 23;
localparam MOD_PROFILE_COMMAND_CMD_0_RESET = 24'h0;
localparam MOD_PROFILE_COMMAND_USEMASK = 64'hFFFFFFFFFFFF;
localparam MOD_PROFILE_COMMAND_RO_MASK = 64'h0;
localparam MOD_PROFILE_COMMAND_WO_MASK = 64'h0;
localparam MOD_PROFILE_COMMAND_RESET = 64'h0;

typedef struct packed {
    logic [12:0] reserved0;  // RSVD
    logic  [8:0] OFFSET_2;  // RW
    logic  [7:0] PROTOCOL_ID_2;  // RW
    logic  [8:0] OFFSET_1;  // RW
    logic  [7:0] PROTOCOL_ID_1;  // RW
    logic  [8:0] OFFSET_0;  // RW
    logic  [7:0] PROTOCOL_ID_0;  // RW
} MOD_PROFILE_FIELD_t;

localparam MOD_PROFILE_FIELD_REG_STRIDE = 48'h8;
localparam MOD_PROFILE_FIELD_REG_ENTRIES = 8;
localparam MOD_PROFILE_FIELD_REGFILE_STRIDE = 48'h40;
localparam MOD_PROFILE_FIELD_REGFILE_ENTRIES = 64;
localparam MOD_PROFILE_FIELD_CR_ADDR = 48'h2000;
localparam MOD_PROFILE_FIELD_SIZE = 64;
localparam MOD_PROFILE_FIELD_OFFSET_2_LO = 42;
localparam MOD_PROFILE_FIELD_OFFSET_2_HI = 50;
localparam MOD_PROFILE_FIELD_OFFSET_2_RESET = 9'h0;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_2_LO = 34;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_2_HI = 41;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_2_RESET = 8'hff;
localparam MOD_PROFILE_FIELD_OFFSET_1_LO = 25;
localparam MOD_PROFILE_FIELD_OFFSET_1_HI = 33;
localparam MOD_PROFILE_FIELD_OFFSET_1_RESET = 9'h0;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_1_LO = 17;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_1_HI = 24;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_1_RESET = 8'hff;
localparam MOD_PROFILE_FIELD_OFFSET_0_LO = 8;
localparam MOD_PROFILE_FIELD_OFFSET_0_HI = 16;
localparam MOD_PROFILE_FIELD_OFFSET_0_RESET = 9'h0;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_0_LO = 0;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_0_HI = 7;
localparam MOD_PROFILE_FIELD_PROTOCOL_ID_0_RESET = 8'hff;
localparam MOD_PROFILE_FIELD_USEMASK = 64'h7FFFFFFFFFFFF;
localparam MOD_PROFILE_FIELD_RO_MASK = 64'h0;
localparam MOD_PROFILE_FIELD_WO_MASK = 64'h0;
localparam MOD_PROFILE_FIELD_RESET = 64'h3FC01FE00FF;

typedef struct packed {
    logic  [7:0] VALUE7;  // RW
    logic  [7:0] VALUE6;  // RW
    logic  [7:0] VALUE5;  // RW
    logic  [7:0] VALUE4;  // RW
    logic  [7:0] VALUE3;  // RW
    logic  [7:0] VALUE2;  // RW
    logic  [7:0] VALUE1;  // RW
    logic  [7:0] VALUE0;  // RW
} MOD_MAP_DUAL_t;

localparam MOD_MAP_DUAL_REG_STRIDE = 48'h8;
localparam MOD_MAP_DUAL_REG_ENTRIES = 8;
localparam MOD_MAP_DUAL_REGFILE_STRIDE = 48'h40;
localparam MOD_MAP_DUAL_REGFILE_ENTRIES = 1024;
localparam MOD_MAP_DUAL_CR_ADDR = 48'h10000;
localparam MOD_MAP_DUAL_SIZE = 64;
localparam MOD_MAP_DUAL_VALUE7_LO = 56;
localparam MOD_MAP_DUAL_VALUE7_HI = 63;
localparam MOD_MAP_DUAL_VALUE7_RESET = 8'h0;
localparam MOD_MAP_DUAL_VALUE6_LO = 48;
localparam MOD_MAP_DUAL_VALUE6_HI = 55;
localparam MOD_MAP_DUAL_VALUE6_RESET = 8'h0;
localparam MOD_MAP_DUAL_VALUE5_LO = 40;
localparam MOD_MAP_DUAL_VALUE5_HI = 47;
localparam MOD_MAP_DUAL_VALUE5_RESET = 8'h0;
localparam MOD_MAP_DUAL_VALUE4_LO = 32;
localparam MOD_MAP_DUAL_VALUE4_HI = 39;
localparam MOD_MAP_DUAL_VALUE4_RESET = 8'h0;
localparam MOD_MAP_DUAL_VALUE3_LO = 24;
localparam MOD_MAP_DUAL_VALUE3_HI = 31;
localparam MOD_MAP_DUAL_VALUE3_RESET = 8'h0;
localparam MOD_MAP_DUAL_VALUE2_LO = 16;
localparam MOD_MAP_DUAL_VALUE2_HI = 23;
localparam MOD_MAP_DUAL_VALUE2_RESET = 8'h0;
localparam MOD_MAP_DUAL_VALUE1_LO = 8;
localparam MOD_MAP_DUAL_VALUE1_HI = 15;
localparam MOD_MAP_DUAL_VALUE1_RESET = 8'h0;
localparam MOD_MAP_DUAL_VALUE0_LO = 0;
localparam MOD_MAP_DUAL_VALUE0_HI = 7;
localparam MOD_MAP_DUAL_VALUE0_RESET = 8'h0;
localparam MOD_MAP_DUAL_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam MOD_MAP_DUAL_RO_MASK = 64'h0;
localparam MOD_MAP_DUAL_WO_MASK = 64'h0;
localparam MOD_MAP_DUAL_RESET = 64'h0;

typedef struct packed {
    logic [15:0] VALUE3;  // RW
    logic [15:0] VALUE2;  // RW
    logic [15:0] VALUE1;  // RW
    logic [15:0] VALUE0;  // RW
} MOD_MAP_t;

localparam MOD_MAP_REG_STRIDE = 48'h8;
localparam MOD_MAP_REG_ENTRIES = 512;
localparam MOD_MAP_REGFILE_STRIDE = 48'h1000;
localparam MOD_MAP_REGFILE_ENTRIES = 4;
localparam MOD_MAP_CR_ADDR = 48'h20000;
localparam MOD_MAP_SIZE = 64;
localparam MOD_MAP_VALUE3_LO = 48;
localparam MOD_MAP_VALUE3_HI = 63;
localparam MOD_MAP_VALUE3_RESET = 16'h0;
localparam MOD_MAP_VALUE2_LO = 32;
localparam MOD_MAP_VALUE2_HI = 47;
localparam MOD_MAP_VALUE2_RESET = 16'h0;
localparam MOD_MAP_VALUE1_LO = 16;
localparam MOD_MAP_VALUE1_HI = 31;
localparam MOD_MAP_VALUE1_RESET = 16'h0;
localparam MOD_MAP_VALUE0_LO = 0;
localparam MOD_MAP_VALUE0_HI = 15;
localparam MOD_MAP_VALUE0_RESET = 16'h0;
localparam MOD_MAP_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam MOD_MAP_RO_MASK = 64'h0;
localparam MOD_MAP_WO_MASK = 64'h0;
localparam MOD_MAP_RESET = 64'h0;

typedef struct packed {
    logic  [0:0] reserved0;  // RSVD
    logic  [8:0] GROUP_7;  // RW
    logic  [8:0] GROUP_6;  // RW
    logic  [8:0] GROUP_5;  // RW
    logic  [8:0] GROUP_4;  // RW
    logic  [8:0] GROUP_3;  // RW
    logic  [8:0] GROUP_2;  // RW
    logic  [8:0] GROUP_1;  // RW
} MOD_PROFILE_GROUP_t;

localparam MOD_PROFILE_GROUP_REG_STRIDE = 48'h8;
localparam MOD_PROFILE_GROUP_REG_ENTRIES = 64;
localparam MOD_PROFILE_GROUP_CR_ADDR = 48'h24000;
localparam MOD_PROFILE_GROUP_SIZE = 64;
localparam MOD_PROFILE_GROUP_GROUP_7_LO = 54;
localparam MOD_PROFILE_GROUP_GROUP_7_HI = 62;
localparam MOD_PROFILE_GROUP_GROUP_7_RESET = 9'h0;
localparam MOD_PROFILE_GROUP_GROUP_6_LO = 45;
localparam MOD_PROFILE_GROUP_GROUP_6_HI = 53;
localparam MOD_PROFILE_GROUP_GROUP_6_RESET = 9'h0;
localparam MOD_PROFILE_GROUP_GROUP_5_LO = 36;
localparam MOD_PROFILE_GROUP_GROUP_5_HI = 44;
localparam MOD_PROFILE_GROUP_GROUP_5_RESET = 9'h0;
localparam MOD_PROFILE_GROUP_GROUP_4_LO = 27;
localparam MOD_PROFILE_GROUP_GROUP_4_HI = 35;
localparam MOD_PROFILE_GROUP_GROUP_4_RESET = 9'h0;
localparam MOD_PROFILE_GROUP_GROUP_3_LO = 18;
localparam MOD_PROFILE_GROUP_GROUP_3_HI = 26;
localparam MOD_PROFILE_GROUP_GROUP_3_RESET = 9'h0;
localparam MOD_PROFILE_GROUP_GROUP_2_LO = 9;
localparam MOD_PROFILE_GROUP_GROUP_2_HI = 17;
localparam MOD_PROFILE_GROUP_GROUP_2_RESET = 9'h0;
localparam MOD_PROFILE_GROUP_GROUP_1_LO = 0;
localparam MOD_PROFILE_GROUP_GROUP_1_HI = 8;
localparam MOD_PROFILE_GROUP_GROUP_1_RESET = 9'h0;
localparam MOD_PROFILE_GROUP_USEMASK = 64'h7FFFFFFFFFFFFFFF;
localparam MOD_PROFILE_GROUP_RO_MASK = 64'h0;
localparam MOD_PROFILE_GROUP_WO_MASK = 64'h0;
localparam MOD_PROFILE_GROUP_RESET = 64'h0;

typedef struct packed {
    logic  [0:0] reserved0;  // RSVD
    logic  [0:0] STORE_PORT;  // RW
    logic  [0:0] STORE_VSI;  // RW
    logic  [4:0] METADATA_TYPE0;  // RW
    logic  [7:0] METADATA_BYTE_OFFSET0;  // RW
    logic [15:0] METADATA_VALUE0;  // RW
    logic [15:0] METADATA_MASK0;  // RW
    logic  [0:0] AUTO_LEARN;  // RW
    logic  [0:0] RECIRCULATE;  // RW
    logic  [0:0] PRE_MOD;  // RW
    logic  [0:0] TRUNC;  // RW
    logic [11:0] MIRROR_DST;  // RW
} MOD_MIRROR_PROFILE_TABLE0_t;

localparam MOD_MIRROR_PROFILE_TABLE0_REG_STRIDE = 48'h8;
localparam MOD_MIRROR_PROFILE_TABLE0_REG_ENTRIES = 64;
localparam MOD_MIRROR_PROFILE_TABLE0_CR_ADDR = 48'h24200;
localparam MOD_MIRROR_PROFILE_TABLE0_SIZE = 64;
localparam MOD_MIRROR_PROFILE_TABLE0_STORE_PORT_LO = 62;
localparam MOD_MIRROR_PROFILE_TABLE0_STORE_PORT_HI = 62;
localparam MOD_MIRROR_PROFILE_TABLE0_STORE_PORT_RESET = 1'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_STORE_VSI_LO = 61;
localparam MOD_MIRROR_PROFILE_TABLE0_STORE_VSI_HI = 61;
localparam MOD_MIRROR_PROFILE_TABLE0_STORE_VSI_RESET = 1'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_TYPE0_LO = 56;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_TYPE0_HI = 60;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_TYPE0_RESET = 5'h1f;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_BYTE_OFFSET0_LO = 48;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_BYTE_OFFSET0_HI = 55;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_BYTE_OFFSET0_RESET = 8'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_VALUE0_LO = 32;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_VALUE0_HI = 47;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_VALUE0_RESET = 16'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_MASK0_LO = 16;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_MASK0_HI = 31;
localparam MOD_MIRROR_PROFILE_TABLE0_METADATA_MASK0_RESET = 16'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_AUTO_LEARN_LO = 15;
localparam MOD_MIRROR_PROFILE_TABLE0_AUTO_LEARN_HI = 15;
localparam MOD_MIRROR_PROFILE_TABLE0_AUTO_LEARN_RESET = 1'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_RECIRCULATE_LO = 14;
localparam MOD_MIRROR_PROFILE_TABLE0_RECIRCULATE_HI = 14;
localparam MOD_MIRROR_PROFILE_TABLE0_RECIRCULATE_RESET = 1'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_PRE_MOD_LO = 13;
localparam MOD_MIRROR_PROFILE_TABLE0_PRE_MOD_HI = 13;
localparam MOD_MIRROR_PROFILE_TABLE0_PRE_MOD_RESET = 1'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_TRUNC_LO = 12;
localparam MOD_MIRROR_PROFILE_TABLE0_TRUNC_HI = 12;
localparam MOD_MIRROR_PROFILE_TABLE0_TRUNC_RESET = 1'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_MIRROR_DST_LO = 0;
localparam MOD_MIRROR_PROFILE_TABLE0_MIRROR_DST_HI = 11;
localparam MOD_MIRROR_PROFILE_TABLE0_MIRROR_DST_RESET = 12'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_USEMASK = 64'h7FFFFFFFFFFFFFFF;
localparam MOD_MIRROR_PROFILE_TABLE0_RO_MASK = 64'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_WO_MASK = 64'h0;
localparam MOD_MIRROR_PROFILE_TABLE0_RESET = 64'h1F00000000000000;

typedef struct packed {
    logic [18:0] reserved0;  // RSVD
    logic  [4:0] METADATA_TYPE1;  // RW
    logic  [7:0] METADATA_BYTE_OFFSET1;  // RW
    logic [15:0] METADATA_VALUE1;  // RW
    logic [15:0] METADATA_MASK1;  // RW
} MOD_MIRROR_PROFILE_TABLE1_t;

localparam MOD_MIRROR_PROFILE_TABLE1_REG_STRIDE = 48'h8;
localparam MOD_MIRROR_PROFILE_TABLE1_REG_ENTRIES = 64;
localparam MOD_MIRROR_PROFILE_TABLE1_CR_ADDR = 48'h24400;
localparam MOD_MIRROR_PROFILE_TABLE1_SIZE = 64;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_TYPE1_LO = 40;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_TYPE1_HI = 44;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_TYPE1_RESET = 5'h1f;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_BYTE_OFFSET1_LO = 32;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_BYTE_OFFSET1_HI = 39;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_BYTE_OFFSET1_RESET = 8'h0;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_VALUE1_LO = 16;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_VALUE1_HI = 31;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_VALUE1_RESET = 16'h0;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_MASK1_LO = 0;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_MASK1_HI = 15;
localparam MOD_MIRROR_PROFILE_TABLE1_METADATA_MASK1_RESET = 16'h0;
localparam MOD_MIRROR_PROFILE_TABLE1_USEMASK = 64'h1FFFFFFFFFFF;
localparam MOD_MIRROR_PROFILE_TABLE1_RO_MASK = 64'h0;
localparam MOD_MIRROR_PROFILE_TABLE1_WO_MASK = 64'h0;
localparam MOD_MIRROR_PROFILE_TABLE1_RESET = 64'h1F0000000000;

typedef struct packed {
    logic [25:0] reserved0;  // RSVD
    logic [13:0] DST_Q;  // RW
    logic  [0:0] FUNC_VALID;  // RW
    logic  [0:0] reserved1;  // RSVD
    logic  [5:0] PF_NUM;  // RW
    logic  [1:0] reserved2;  // RSVD
    logic  [1:0] FUNCTION_TYPE;  // RW
    logic [11:0] FUNCTION_NUM;  // RW
} MOD_MIRROR_PROFILE_TABLE2_t;

localparam MOD_MIRROR_PROFILE_TABLE2_REG_STRIDE = 48'h8;
localparam MOD_MIRROR_PROFILE_TABLE2_REG_ENTRIES = 64;
localparam MOD_MIRROR_PROFILE_TABLE2_CR_ADDR = 48'h24600;
localparam MOD_MIRROR_PROFILE_TABLE2_SIZE = 64;
localparam MOD_MIRROR_PROFILE_TABLE2_DST_Q_LO = 24;
localparam MOD_MIRROR_PROFILE_TABLE2_DST_Q_HI = 37;
localparam MOD_MIRROR_PROFILE_TABLE2_DST_Q_RESET = 14'h0;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNC_VALID_LO = 23;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNC_VALID_HI = 23;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNC_VALID_RESET = 1'h0;
localparam MOD_MIRROR_PROFILE_TABLE2_PF_NUM_LO = 16;
localparam MOD_MIRROR_PROFILE_TABLE2_PF_NUM_HI = 21;
localparam MOD_MIRROR_PROFILE_TABLE2_PF_NUM_RESET = 6'h0;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNCTION_TYPE_LO = 12;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNCTION_TYPE_HI = 13;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNCTION_TYPE_RESET = 2'h0;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNCTION_NUM_LO = 0;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNCTION_NUM_HI = 11;
localparam MOD_MIRROR_PROFILE_TABLE2_FUNCTION_NUM_RESET = 12'h0;
localparam MOD_MIRROR_PROFILE_TABLE2_USEMASK = 64'h3FFFBF3FFF;
localparam MOD_MIRROR_PROFILE_TABLE2_RO_MASK = 64'h0;
localparam MOD_MIRROR_PROFILE_TABLE2_WO_MASK = 64'h0;
localparam MOD_MIRROR_PROFILE_TABLE2_RESET = 64'h0;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic  [3:0] OUTPUT_SHIFT;  // RW
    logic [15:0] OUTPUT_MASK;  // RW
    logic  [3:0] BASE_MASK_LEN;  // RW
    logic  [3:0] BASE_SHIFT_RIGHT;  // RW
    logic  [3:0] IDX_MASK_LEN;  // RW
    logic  [3:0] IDX_SHIFT_RIGHT;  // RW
} MOD_MAP_CFG_t;

localparam MOD_MAP_CFG_REG_STRIDE = 48'h8;
localparam MOD_MAP_CFG_REG_ENTRIES = 4;
localparam MOD_MAP_CFG_CR_ADDR = 48'h24800;
localparam MOD_MAP_CFG_SIZE = 64;
localparam MOD_MAP_CFG_OUTPUT_SHIFT_LO = 32;
localparam MOD_MAP_CFG_OUTPUT_SHIFT_HI = 35;
localparam MOD_MAP_CFG_OUTPUT_SHIFT_RESET = 4'h0;
localparam MOD_MAP_CFG_OUTPUT_MASK_LO = 16;
localparam MOD_MAP_CFG_OUTPUT_MASK_HI = 31;
localparam MOD_MAP_CFG_OUTPUT_MASK_RESET = 16'h0;
localparam MOD_MAP_CFG_BASE_MASK_LEN_LO = 12;
localparam MOD_MAP_CFG_BASE_MASK_LEN_HI = 15;
localparam MOD_MAP_CFG_BASE_MASK_LEN_RESET = 4'h0;
localparam MOD_MAP_CFG_BASE_SHIFT_RIGHT_LO = 8;
localparam MOD_MAP_CFG_BASE_SHIFT_RIGHT_HI = 11;
localparam MOD_MAP_CFG_BASE_SHIFT_RIGHT_RESET = 4'h0;
localparam MOD_MAP_CFG_IDX_MASK_LEN_LO = 4;
localparam MOD_MAP_CFG_IDX_MASK_LEN_HI = 7;
localparam MOD_MAP_CFG_IDX_MASK_LEN_RESET = 4'h0;
localparam MOD_MAP_CFG_IDX_SHIFT_RIGHT_LO = 0;
localparam MOD_MAP_CFG_IDX_SHIFT_RIGHT_HI = 3;
localparam MOD_MAP_CFG_IDX_SHIFT_RIGHT_RESET = 4'h0;
localparam MOD_MAP_CFG_USEMASK = 64'hFFFFFFFFF;
localparam MOD_MAP_CFG_RO_MASK = 64'h0;
localparam MOD_MAP_CFG_WO_MASK = 64'h0;
localparam MOD_MAP_CFG_RESET = 64'h0;

typedef struct packed {
    logic [29:0] reserved0;  // RSVD
    logic  [3:0] OUTPUT_SHIFT;  // RW
    logic [15:0] OUTPUT_MASK;  // RW
    logic  [2:0] IDX1_MASK_LEN;  // RW
    logic  [2:0] IDX1_SHIFT_RIGHT;  // RW
    logic  [3:0] IDX0_MASK_LEN;  // RW
    logic  [3:0] IDX0_SHIFT_RIGHT;  // RW
} MOD_MAP_DUAL_CFG_t;

localparam MOD_MAP_DUAL_CFG_REG_STRIDE = 48'h8;
localparam MOD_MAP_DUAL_CFG_REG_ENTRIES = 1;
localparam MOD_MAP_DUAL_CFG_CR_ADDR = 48'h24820;
localparam MOD_MAP_DUAL_CFG_SIZE = 64;
localparam MOD_MAP_DUAL_CFG_OUTPUT_SHIFT_LO = 30;
localparam MOD_MAP_DUAL_CFG_OUTPUT_SHIFT_HI = 33;
localparam MOD_MAP_DUAL_CFG_OUTPUT_SHIFT_RESET = 4'h0;
localparam MOD_MAP_DUAL_CFG_OUTPUT_MASK_LO = 14;
localparam MOD_MAP_DUAL_CFG_OUTPUT_MASK_HI = 29;
localparam MOD_MAP_DUAL_CFG_OUTPUT_MASK_RESET = 16'h0;
localparam MOD_MAP_DUAL_CFG_IDX1_MASK_LEN_LO = 11;
localparam MOD_MAP_DUAL_CFG_IDX1_MASK_LEN_HI = 13;
localparam MOD_MAP_DUAL_CFG_IDX1_MASK_LEN_RESET = 3'h0;
localparam MOD_MAP_DUAL_CFG_IDX1_SHIFT_RIGHT_LO = 8;
localparam MOD_MAP_DUAL_CFG_IDX1_SHIFT_RIGHT_HI = 10;
localparam MOD_MAP_DUAL_CFG_IDX1_SHIFT_RIGHT_RESET = 3'h0;
localparam MOD_MAP_DUAL_CFG_IDX0_MASK_LEN_LO = 4;
localparam MOD_MAP_DUAL_CFG_IDX0_MASK_LEN_HI = 7;
localparam MOD_MAP_DUAL_CFG_IDX0_MASK_LEN_RESET = 4'h0;
localparam MOD_MAP_DUAL_CFG_IDX0_SHIFT_RIGHT_LO = 0;
localparam MOD_MAP_DUAL_CFG_IDX0_SHIFT_RIGHT_HI = 3;
localparam MOD_MAP_DUAL_CFG_IDX0_SHIFT_RIGHT_RESET = 4'h0;
localparam MOD_MAP_DUAL_CFG_USEMASK = 64'h3FFFFFFFF;
localparam MOD_MAP_DUAL_CFG_RO_MASK = 64'h0;
localparam MOD_MAP_DUAL_CFG_WO_MASK = 64'h0;
localparam MOD_MAP_DUAL_CFG_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic  [7:0] IPV6_2;  // RW
    logic  [7:0] IPV6_1;  // RW
    logic  [7:0] IPV6_0;  // RW
    logic  [7:0] IPV4_2;  // RW
    logic  [7:0] IPV4_1;  // RW
    logic  [7:0] IPV4_0;  // RW
} MOD_CSUM_CFG1_t;

localparam MOD_CSUM_CFG1_REG_STRIDE = 48'h8;
localparam MOD_CSUM_CFG1_REG_ENTRIES = 1;
localparam MOD_CSUM_CFG1_CR_ADDR = 48'h24828;
localparam MOD_CSUM_CFG1_SIZE = 64;
localparam MOD_CSUM_CFG1_IPV6_2_LO = 40;
localparam MOD_CSUM_CFG1_IPV6_2_HI = 47;
localparam MOD_CSUM_CFG1_IPV6_2_RESET = 8'hff;
localparam MOD_CSUM_CFG1_IPV6_1_LO = 32;
localparam MOD_CSUM_CFG1_IPV6_1_HI = 39;
localparam MOD_CSUM_CFG1_IPV6_1_RESET = 8'hff;
localparam MOD_CSUM_CFG1_IPV6_0_LO = 24;
localparam MOD_CSUM_CFG1_IPV6_0_HI = 31;
localparam MOD_CSUM_CFG1_IPV6_0_RESET = 8'hff;
localparam MOD_CSUM_CFG1_IPV4_2_LO = 16;
localparam MOD_CSUM_CFG1_IPV4_2_HI = 23;
localparam MOD_CSUM_CFG1_IPV4_2_RESET = 8'hff;
localparam MOD_CSUM_CFG1_IPV4_1_LO = 8;
localparam MOD_CSUM_CFG1_IPV4_1_HI = 15;
localparam MOD_CSUM_CFG1_IPV4_1_RESET = 8'hff;
localparam MOD_CSUM_CFG1_IPV4_0_LO = 0;
localparam MOD_CSUM_CFG1_IPV4_0_HI = 7;
localparam MOD_CSUM_CFG1_IPV4_0_RESET = 8'hff;
localparam MOD_CSUM_CFG1_USEMASK = 64'hFFFFFFFFFFFF;
localparam MOD_CSUM_CFG1_RO_MASK = 64'h0;
localparam MOD_CSUM_CFG1_WO_MASK = 64'h0;
localparam MOD_CSUM_CFG1_RESET = 64'hFFFFFFFFFFFF;

typedef struct packed {
    logic  [7:0] reserved0;  // RSVD
    logic  [7:0] SCTP;  // RW
    logic  [7:0] TCP_2;  // RW
    logic  [7:0] TCP_1;  // RW
    logic  [7:0] TCP_0;  // RW
    logic  [7:0] UDP_2;  // RW
    logic  [7:0] UDP_1;  // RW
    logic  [7:0] UDP_0;  // RW
} MOD_CSUM_CFG2_t;

localparam MOD_CSUM_CFG2_REG_STRIDE = 48'h8;
localparam MOD_CSUM_CFG2_REG_ENTRIES = 1;
localparam MOD_CSUM_CFG2_CR_ADDR = 48'h24830;
localparam MOD_CSUM_CFG2_SIZE = 64;
localparam MOD_CSUM_CFG2_SCTP_LO = 48;
localparam MOD_CSUM_CFG2_SCTP_HI = 55;
localparam MOD_CSUM_CFG2_SCTP_RESET = 8'hff;
localparam MOD_CSUM_CFG2_TCP_2_LO = 40;
localparam MOD_CSUM_CFG2_TCP_2_HI = 47;
localparam MOD_CSUM_CFG2_TCP_2_RESET = 8'hff;
localparam MOD_CSUM_CFG2_TCP_1_LO = 32;
localparam MOD_CSUM_CFG2_TCP_1_HI = 39;
localparam MOD_CSUM_CFG2_TCP_1_RESET = 8'hff;
localparam MOD_CSUM_CFG2_TCP_0_LO = 24;
localparam MOD_CSUM_CFG2_TCP_0_HI = 31;
localparam MOD_CSUM_CFG2_TCP_0_RESET = 8'hff;
localparam MOD_CSUM_CFG2_UDP_2_LO = 16;
localparam MOD_CSUM_CFG2_UDP_2_HI = 23;
localparam MOD_CSUM_CFG2_UDP_2_RESET = 8'hff;
localparam MOD_CSUM_CFG2_UDP_1_LO = 8;
localparam MOD_CSUM_CFG2_UDP_1_HI = 15;
localparam MOD_CSUM_CFG2_UDP_1_RESET = 8'hff;
localparam MOD_CSUM_CFG2_UDP_0_LO = 0;
localparam MOD_CSUM_CFG2_UDP_0_HI = 7;
localparam MOD_CSUM_CFG2_UDP_0_RESET = 8'hff;
localparam MOD_CSUM_CFG2_USEMASK = 64'hFFFFFFFFFFFFFF;
localparam MOD_CSUM_CFG2_RO_MASK = 64'h0;
localparam MOD_CSUM_CFG2_WO_MASK = 64'h0;
localparam MOD_CSUM_CFG2_RESET = 64'hFFFFFFFFFFFFFF;

typedef struct packed {
    logic [52:0] reserved0;  // RSVD
    logic  [0:0] SCTP_EN;  // RW
    logic  [0:0] D1_TCP_EN;  // RW
    logic  [0:0] D0_TCP_EN;  // RW
    logic  [0:0] D1_UDP_EN;  // RW
    logic  [0:0] D0_UDP_EN;  // RW
    logic  [0:0] D2_IPV6_EN;  // RW
    logic  [0:0] D1_IPV6_EN;  // RW
    logic  [0:0] D0_IPV6_EN;  // RW
    logic  [0:0] D2_IPV4_EN;  // RW
    logic  [0:0] D1_IPV4_EN;  // RW
    logic  [0:0] D0_IPV4_EN;  // RW
} MOD_CSUM_EN_CFG_t;

localparam MOD_CSUM_EN_CFG_REG_STRIDE = 48'h8;
localparam MOD_CSUM_EN_CFG_REG_ENTRIES = 1;
localparam [47:0] MOD_CSUM_EN_CFG_CR_ADDR = 48'h24838;
localparam MOD_CSUM_EN_CFG_SIZE = 64;
localparam MOD_CSUM_EN_CFG_SCTP_EN_LO = 10;
localparam MOD_CSUM_EN_CFG_SCTP_EN_HI = 10;
localparam MOD_CSUM_EN_CFG_SCTP_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D1_TCP_EN_LO = 9;
localparam MOD_CSUM_EN_CFG_D1_TCP_EN_HI = 9;
localparam MOD_CSUM_EN_CFG_D1_TCP_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D0_TCP_EN_LO = 8;
localparam MOD_CSUM_EN_CFG_D0_TCP_EN_HI = 8;
localparam MOD_CSUM_EN_CFG_D0_TCP_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D1_UDP_EN_LO = 7;
localparam MOD_CSUM_EN_CFG_D1_UDP_EN_HI = 7;
localparam MOD_CSUM_EN_CFG_D1_UDP_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D0_UDP_EN_LO = 6;
localparam MOD_CSUM_EN_CFG_D0_UDP_EN_HI = 6;
localparam MOD_CSUM_EN_CFG_D0_UDP_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D2_IPV6_EN_LO = 5;
localparam MOD_CSUM_EN_CFG_D2_IPV6_EN_HI = 5;
localparam MOD_CSUM_EN_CFG_D2_IPV6_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D1_IPV6_EN_LO = 4;
localparam MOD_CSUM_EN_CFG_D1_IPV6_EN_HI = 4;
localparam MOD_CSUM_EN_CFG_D1_IPV6_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D0_IPV6_EN_LO = 3;
localparam MOD_CSUM_EN_CFG_D0_IPV6_EN_HI = 3;
localparam MOD_CSUM_EN_CFG_D0_IPV6_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D2_IPV4_EN_LO = 2;
localparam MOD_CSUM_EN_CFG_D2_IPV4_EN_HI = 2;
localparam MOD_CSUM_EN_CFG_D2_IPV4_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D1_IPV4_EN_LO = 1;
localparam MOD_CSUM_EN_CFG_D1_IPV4_EN_HI = 1;
localparam MOD_CSUM_EN_CFG_D1_IPV4_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_D0_IPV4_EN_LO = 0;
localparam MOD_CSUM_EN_CFG_D0_IPV4_EN_HI = 0;
localparam MOD_CSUM_EN_CFG_D0_IPV4_EN_RESET = 1'h1;
localparam MOD_CSUM_EN_CFG_USEMASK = 64'h7FF;
localparam MOD_CSUM_EN_CFG_RO_MASK = 64'h0;
localparam MOD_CSUM_EN_CFG_WO_MASK = 64'h0;
localparam MOD_CSUM_EN_CFG_RESET = 64'h7FF;

typedef struct packed {
    MOD_CSUM_EN_CFG_t  MOD_CSUM_EN_CFG;
} mby_ppe_modify_map_registers_t;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_MOD_PROFILE_COMMAND_t;

typedef logic [7:0] we_MOD_PROFILE_FIELD_t;

typedef logic [7:0] we_MOD_MAP_DUAL_t;

typedef logic [7:0] we_MOD_MAP_t;

typedef logic [7:0] we_MOD_PROFILE_GROUP_t;

typedef logic [7:0] we_MOD_MIRROR_PROFILE_TABLE0_t;

typedef logic [7:0] we_MOD_MIRROR_PROFILE_TABLE1_t;

typedef logic [7:0] we_MOD_MIRROR_PROFILE_TABLE2_t;

typedef logic [7:0] we_MOD_MAP_CFG_t;

typedef logic [7:0] we_MOD_MAP_DUAL_CFG_t;

typedef logic [7:0] we_MOD_CSUM_CFG1_t;

typedef logic [7:0] we_MOD_CSUM_CFG2_t;

typedef struct packed {
    we_MOD_PROFILE_COMMAND_t MOD_PROFILE_COMMAND;
    we_MOD_PROFILE_FIELD_t MOD_PROFILE_FIELD;
    we_MOD_MAP_DUAL_t MOD_MAP_DUAL;
    we_MOD_MAP_t MOD_MAP;
    we_MOD_PROFILE_GROUP_t MOD_PROFILE_GROUP;
    we_MOD_MIRROR_PROFILE_TABLE0_t MOD_MIRROR_PROFILE_TABLE0;
    we_MOD_MIRROR_PROFILE_TABLE1_t MOD_MIRROR_PROFILE_TABLE1;
    we_MOD_MIRROR_PROFILE_TABLE2_t MOD_MIRROR_PROFILE_TABLE2;
    we_MOD_MAP_CFG_t MOD_MAP_CFG;
    we_MOD_MAP_DUAL_CFG_t MOD_MAP_DUAL_CFG;
    we_MOD_CSUM_CFG1_t MOD_CSUM_CFG1;
    we_MOD_CSUM_CFG2_t MOD_CSUM_CFG2;
} mby_ppe_modify_map_handcoded_t;

typedef logic [7:0] re_MOD_PROFILE_COMMAND_t;

typedef logic [7:0] re_MOD_PROFILE_FIELD_t;

typedef logic [7:0] re_MOD_MAP_DUAL_t;

typedef logic [7:0] re_MOD_MAP_t;

typedef logic [7:0] re_MOD_PROFILE_GROUP_t;

typedef logic [7:0] re_MOD_MIRROR_PROFILE_TABLE0_t;

typedef logic [7:0] re_MOD_MIRROR_PROFILE_TABLE1_t;

typedef logic [7:0] re_MOD_MIRROR_PROFILE_TABLE2_t;

typedef logic [7:0] re_MOD_MAP_CFG_t;

typedef logic [7:0] re_MOD_MAP_DUAL_CFG_t;

typedef logic [7:0] re_MOD_CSUM_CFG1_t;

typedef logic [7:0] re_MOD_CSUM_CFG2_t;

typedef struct packed {
    re_MOD_PROFILE_COMMAND_t MOD_PROFILE_COMMAND;
    re_MOD_PROFILE_FIELD_t MOD_PROFILE_FIELD;
    re_MOD_MAP_DUAL_t MOD_MAP_DUAL;
    re_MOD_MAP_t MOD_MAP;
    re_MOD_PROFILE_GROUP_t MOD_PROFILE_GROUP;
    re_MOD_MIRROR_PROFILE_TABLE0_t MOD_MIRROR_PROFILE_TABLE0;
    re_MOD_MIRROR_PROFILE_TABLE1_t MOD_MIRROR_PROFILE_TABLE1;
    re_MOD_MIRROR_PROFILE_TABLE2_t MOD_MIRROR_PROFILE_TABLE2;
    re_MOD_MAP_CFG_t MOD_MAP_CFG;
    re_MOD_MAP_DUAL_CFG_t MOD_MAP_DUAL_CFG;
    re_MOD_CSUM_CFG1_t MOD_CSUM_CFG1;
    re_MOD_CSUM_CFG2_t MOD_CSUM_CFG2;
} mby_ppe_modify_map_hc_re_t;

typedef logic handcode_rvalid_MOD_PROFILE_COMMAND_t;

typedef logic handcode_rvalid_MOD_PROFILE_FIELD_t;

typedef logic handcode_rvalid_MOD_MAP_DUAL_t;

typedef logic handcode_rvalid_MOD_MAP_t;

typedef logic handcode_rvalid_MOD_PROFILE_GROUP_t;

typedef logic handcode_rvalid_MOD_MIRROR_PROFILE_TABLE0_t;

typedef logic handcode_rvalid_MOD_MIRROR_PROFILE_TABLE1_t;

typedef logic handcode_rvalid_MOD_MIRROR_PROFILE_TABLE2_t;

typedef logic handcode_rvalid_MOD_MAP_CFG_t;

typedef logic handcode_rvalid_MOD_MAP_DUAL_CFG_t;

typedef logic handcode_rvalid_MOD_CSUM_CFG1_t;

typedef logic handcode_rvalid_MOD_CSUM_CFG2_t;

typedef struct packed {
    handcode_rvalid_MOD_PROFILE_COMMAND_t MOD_PROFILE_COMMAND;
    handcode_rvalid_MOD_PROFILE_FIELD_t MOD_PROFILE_FIELD;
    handcode_rvalid_MOD_MAP_DUAL_t MOD_MAP_DUAL;
    handcode_rvalid_MOD_MAP_t MOD_MAP;
    handcode_rvalid_MOD_PROFILE_GROUP_t MOD_PROFILE_GROUP;
    handcode_rvalid_MOD_MIRROR_PROFILE_TABLE0_t MOD_MIRROR_PROFILE_TABLE0;
    handcode_rvalid_MOD_MIRROR_PROFILE_TABLE1_t MOD_MIRROR_PROFILE_TABLE1;
    handcode_rvalid_MOD_MIRROR_PROFILE_TABLE2_t MOD_MIRROR_PROFILE_TABLE2;
    handcode_rvalid_MOD_MAP_CFG_t MOD_MAP_CFG;
    handcode_rvalid_MOD_MAP_DUAL_CFG_t MOD_MAP_DUAL_CFG;
    handcode_rvalid_MOD_CSUM_CFG1_t MOD_CSUM_CFG1;
    handcode_rvalid_MOD_CSUM_CFG2_t MOD_CSUM_CFG2;
} mby_ppe_modify_map_hc_rvalid_t;

typedef logic handcode_wvalid_MOD_PROFILE_COMMAND_t;

typedef logic handcode_wvalid_MOD_PROFILE_FIELD_t;

typedef logic handcode_wvalid_MOD_MAP_DUAL_t;

typedef logic handcode_wvalid_MOD_MAP_t;

typedef logic handcode_wvalid_MOD_PROFILE_GROUP_t;

typedef logic handcode_wvalid_MOD_MIRROR_PROFILE_TABLE0_t;

typedef logic handcode_wvalid_MOD_MIRROR_PROFILE_TABLE1_t;

typedef logic handcode_wvalid_MOD_MIRROR_PROFILE_TABLE2_t;

typedef logic handcode_wvalid_MOD_MAP_CFG_t;

typedef logic handcode_wvalid_MOD_MAP_DUAL_CFG_t;

typedef logic handcode_wvalid_MOD_CSUM_CFG1_t;

typedef logic handcode_wvalid_MOD_CSUM_CFG2_t;

typedef struct packed {
    handcode_wvalid_MOD_PROFILE_COMMAND_t MOD_PROFILE_COMMAND;
    handcode_wvalid_MOD_PROFILE_FIELD_t MOD_PROFILE_FIELD;
    handcode_wvalid_MOD_MAP_DUAL_t MOD_MAP_DUAL;
    handcode_wvalid_MOD_MAP_t MOD_MAP;
    handcode_wvalid_MOD_PROFILE_GROUP_t MOD_PROFILE_GROUP;
    handcode_wvalid_MOD_MIRROR_PROFILE_TABLE0_t MOD_MIRROR_PROFILE_TABLE0;
    handcode_wvalid_MOD_MIRROR_PROFILE_TABLE1_t MOD_MIRROR_PROFILE_TABLE1;
    handcode_wvalid_MOD_MIRROR_PROFILE_TABLE2_t MOD_MIRROR_PROFILE_TABLE2;
    handcode_wvalid_MOD_MAP_CFG_t MOD_MAP_CFG;
    handcode_wvalid_MOD_MAP_DUAL_CFG_t MOD_MAP_DUAL_CFG;
    handcode_wvalid_MOD_CSUM_CFG1_t MOD_CSUM_CFG1;
    handcode_wvalid_MOD_CSUM_CFG2_t MOD_CSUM_CFG2;
} mby_ppe_modify_map_hc_wvalid_t;

typedef logic handcode_error_MOD_PROFILE_COMMAND_t;

typedef logic handcode_error_MOD_PROFILE_FIELD_t;

typedef logic handcode_error_MOD_MAP_DUAL_t;

typedef logic handcode_error_MOD_MAP_t;

typedef logic handcode_error_MOD_PROFILE_GROUP_t;

typedef logic handcode_error_MOD_MIRROR_PROFILE_TABLE0_t;

typedef logic handcode_error_MOD_MIRROR_PROFILE_TABLE1_t;

typedef logic handcode_error_MOD_MIRROR_PROFILE_TABLE2_t;

typedef logic handcode_error_MOD_MAP_CFG_t;

typedef logic handcode_error_MOD_MAP_DUAL_CFG_t;

typedef logic handcode_error_MOD_CSUM_CFG1_t;

typedef logic handcode_error_MOD_CSUM_CFG2_t;

typedef struct packed {
    handcode_error_MOD_PROFILE_COMMAND_t MOD_PROFILE_COMMAND;
    handcode_error_MOD_PROFILE_FIELD_t MOD_PROFILE_FIELD;
    handcode_error_MOD_MAP_DUAL_t MOD_MAP_DUAL;
    handcode_error_MOD_MAP_t MOD_MAP;
    handcode_error_MOD_PROFILE_GROUP_t MOD_PROFILE_GROUP;
    handcode_error_MOD_MIRROR_PROFILE_TABLE0_t MOD_MIRROR_PROFILE_TABLE0;
    handcode_error_MOD_MIRROR_PROFILE_TABLE1_t MOD_MIRROR_PROFILE_TABLE1;
    handcode_error_MOD_MIRROR_PROFILE_TABLE2_t MOD_MIRROR_PROFILE_TABLE2;
    handcode_error_MOD_MAP_CFG_t MOD_MAP_CFG;
    handcode_error_MOD_MAP_DUAL_CFG_t MOD_MAP_DUAL_CFG;
    handcode_error_MOD_CSUM_CFG1_t MOD_CSUM_CFG1;
    handcode_error_MOD_CSUM_CFG2_t MOD_CSUM_CFG2;
} mby_ppe_modify_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    MOD_PROFILE_COMMAND_t MOD_PROFILE_COMMAND;
    MOD_PROFILE_FIELD_t MOD_PROFILE_FIELD;
    MOD_MAP_DUAL_t MOD_MAP_DUAL;
    MOD_MAP_t MOD_MAP;
    MOD_PROFILE_GROUP_t MOD_PROFILE_GROUP;
    MOD_MIRROR_PROFILE_TABLE0_t MOD_MIRROR_PROFILE_TABLE0;
    MOD_MIRROR_PROFILE_TABLE1_t MOD_MIRROR_PROFILE_TABLE1;
    MOD_MIRROR_PROFILE_TABLE2_t MOD_MIRROR_PROFILE_TABLE2;
    MOD_MAP_CFG_t MOD_MAP_CFG;
    MOD_MAP_DUAL_CFG_t MOD_MAP_DUAL_CFG;
    MOD_CSUM_CFG1_t MOD_CSUM_CFG1;
    MOD_CSUM_CFG2_t MOD_CSUM_CFG2;
} mby_ppe_modify_map_hc_reg_read_t;

typedef struct packed {
    MOD_PROFILE_COMMAND_t MOD_PROFILE_COMMAND;
    MOD_PROFILE_FIELD_t MOD_PROFILE_FIELD;
    MOD_MAP_DUAL_t MOD_MAP_DUAL;
    MOD_MAP_t MOD_MAP;
    MOD_PROFILE_GROUP_t MOD_PROFILE_GROUP;
    MOD_MIRROR_PROFILE_TABLE0_t MOD_MIRROR_PROFILE_TABLE0;
    MOD_MIRROR_PROFILE_TABLE1_t MOD_MIRROR_PROFILE_TABLE1;
    MOD_MIRROR_PROFILE_TABLE2_t MOD_MIRROR_PROFILE_TABLE2;
    MOD_MAP_CFG_t MOD_MAP_CFG;
    MOD_MAP_DUAL_CFG_t MOD_MAP_DUAL_CFG;
    MOD_CSUM_CFG1_t MOD_CSUM_CFG1;
    MOD_CSUM_CFG2_t MOD_CSUM_CFG2;
} mby_ppe_modify_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_modify_map_pkg

`endif // MBY_PPE_MODIFY_MAP_PKG_VH
