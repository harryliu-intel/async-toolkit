magic
tech scmos
timestamp 970030226
<< ndiffusion >>
rect -16 118 -8 119
rect -16 114 -8 115
rect -64 99 -61 103
rect -56 99 -51 103
rect -48 99 -45 103
rect -25 81 -8 82
rect -48 73 -32 74
rect -25 73 -8 78
rect -48 65 -32 70
rect -25 65 -8 70
rect -48 57 -32 62
rect -25 57 -8 62
rect -48 49 -32 54
rect -25 49 -8 54
rect -48 41 -32 46
rect -25 45 -8 46
rect -48 37 -32 38
<< pdiffusion >>
rect 8 118 16 119
rect 8 114 16 115
rect 23 110 27 119
rect 46 116 58 117
rect 46 107 58 108
rect 23 103 27 106
rect 46 103 58 104
rect 54 98 58 103
rect 14 81 40 82
rect 14 77 40 78
rect 14 68 40 69
rect 14 64 40 65
rect 28 56 40 64
rect 14 55 40 56
rect 14 51 40 52
rect 14 42 40 43
rect 14 38 40 39
<< ntransistor >>
rect -16 115 -8 118
rect -61 99 -56 103
rect -51 99 -48 103
rect -25 78 -8 81
rect -48 70 -32 73
rect -25 70 -8 73
rect -48 62 -32 65
rect -25 62 -8 65
rect -48 54 -32 57
rect -25 54 -8 57
rect -48 46 -32 49
rect -25 46 -8 49
rect -48 38 -32 41
<< ptransistor >>
rect 8 115 16 118
rect 23 106 27 110
rect 46 104 58 107
rect 14 78 40 81
rect 14 65 40 68
rect 14 52 40 55
rect 14 39 40 42
<< polysilicon >>
rect -61 103 -56 117
rect -20 115 -16 118
rect -8 115 -4 118
rect -51 105 -33 108
rect -51 103 -48 105
rect 4 115 8 118
rect 16 115 20 118
rect 18 106 23 110
rect 27 107 29 110
rect 27 106 31 107
rect 18 104 21 106
rect -61 95 -56 99
rect -51 95 -48 99
rect -28 101 21 104
rect 42 104 46 107
rect 58 104 62 107
rect -52 84 -27 87
rect -30 81 -27 84
rect -30 78 -25 81
rect -8 78 -4 81
rect 1 78 14 81
rect 40 78 44 81
rect 1 73 4 78
rect -52 70 -48 73
rect -32 70 -25 73
rect -8 70 4 73
rect 9 65 14 68
rect 40 65 44 68
rect -52 62 -48 65
rect -32 62 -25 65
rect -8 62 12 65
rect -52 54 -48 57
rect -32 54 -25 57
rect -8 55 12 57
rect -8 54 14 55
rect 9 52 14 54
rect 40 52 44 55
rect -52 46 -48 49
rect -32 46 -25 49
rect -8 47 4 49
rect -8 46 -4 47
rect -52 38 -48 41
rect -32 38 -28 41
rect 4 39 14 42
rect 40 39 44 42
<< ndcontact >>
rect -16 119 -8 127
rect -16 106 -8 114
rect -72 95 -64 103
rect -45 95 -37 103
rect -48 74 -32 82
rect -25 82 -8 90
rect -25 37 -8 45
rect -48 29 -32 37
<< pdcontact >>
rect 8 119 16 127
rect 22 119 30 127
rect 8 106 16 114
rect 46 108 58 116
rect 23 95 31 103
rect 46 95 54 103
rect 14 82 40 90
rect 14 69 40 77
rect 14 56 28 64
rect 14 43 40 51
rect 14 30 40 38
<< psubstratepcontact >>
rect -46 112 -38 120
<< nsubstratencontact >>
rect 46 117 58 125
<< polycontact >>
rect -64 117 -56 125
rect -33 104 -25 112
rect -4 110 4 118
rect 29 107 37 115
rect 62 104 70 112
rect -60 79 -52 87
rect 44 73 52 81
rect 44 60 52 68
rect -60 33 -52 41
rect -4 39 4 47
rect 44 47 52 55
<< metal1 >>
rect -64 117 -56 121
rect -45 121 -21 127
rect -45 120 -8 121
rect -46 119 -8 120
rect 21 121 58 127
rect 8 119 58 121
rect -46 113 -38 119
rect -69 112 -38 113
rect -16 112 -8 114
rect -69 107 -39 112
rect -33 108 -8 112
rect -69 103 -64 107
rect -33 104 -25 108
rect -16 106 -8 108
rect -4 103 4 118
rect 8 112 16 114
rect 29 112 37 115
rect 8 108 37 112
rect 46 108 58 119
rect 8 106 16 108
rect 29 107 37 108
rect 62 104 70 121
rect -72 95 -64 103
rect -45 99 -37 103
rect -45 97 -4 99
rect 23 99 31 103
rect 46 99 54 103
rect 4 97 54 99
rect -45 95 54 97
rect -60 31 -52 87
rect -25 85 -21 90
rect -25 82 -8 85
rect -48 74 -32 82
rect -40 64 -32 74
rect -4 64 4 95
rect 21 85 40 90
rect 14 82 40 85
rect 44 79 52 81
rect 14 69 40 77
rect -40 56 28 64
rect -16 45 -8 56
rect 32 51 40 69
rect 44 67 52 68
rect 44 60 52 61
rect -25 37 -8 45
rect -4 43 4 47
rect 14 43 40 51
rect 44 47 52 49
rect -48 31 -32 37
rect 14 31 40 38
rect -48 25 -21 31
rect 21 30 40 31
<< m2contact >>
rect -64 121 -56 127
rect -21 121 -8 127
rect 8 121 21 127
rect 62 121 70 127
rect -4 97 4 103
rect -21 85 -8 91
rect 8 85 21 91
rect 44 73 52 79
rect 44 61 52 67
rect 44 49 52 55
rect -4 37 4 43
rect -60 25 -52 31
rect -21 25 -3 31
rect 3 25 21 31
<< metal2 >>
rect -64 121 -27 127
rect 27 121 70 127
rect -6 97 6 103
rect 0 73 52 79
rect 0 61 52 67
rect 0 49 52 55
rect -6 37 6 43
rect -60 25 -26 31
<< m3contact >>
rect -21 121 -8 127
rect 8 121 21 127
rect -21 85 -3 91
rect 4 85 21 91
rect -21 25 -3 31
rect 3 25 21 31
<< metal3 >>
rect -21 22 -3 130
rect 3 22 21 130
<< labels >>
rlabel metal1 -68 99 -68 99 3 GND!
rlabel polysilicon -60 104 -60 104 3 _SReset!
rlabel metal1 27 98 27 98 5 x
rlabel metal1 -41 99 -41 99 3 x
rlabel metal2 -60 124 -60 124 5 _SReset!
rlabel ndcontact -12 123 -12 123 5 GND!
rlabel pdcontact 12 123 12 123 5 Vdd!
rlabel metal2 -6 97 -6 103 3 x
rlabel metal2 6 97 6 103 7 x
rlabel metal1 0 114 0 114 1 x
rlabel metal1 18 60 18 60 1 x
rlabel m2contact 18 86 18 86 5 Vdd!
rlabel metal1 18 34 18 34 1 Vdd!
rlabel metal1 -12 41 -12 41 1 x
rlabel polysilicon 41 40 41 40 3 _a0
rlabel polysilicon 41 53 41 53 3 _b0
rlabel polysilicon 41 66 41 66 3 _b1
rlabel polysilicon 41 79 41 79 3 _a1
rlabel metal1 -36 78 -36 78 5 x
rlabel metal1 -36 33 -36 33 1 GND!
rlabel polysilicon -49 39 -49 39 3 _SReset!
rlabel polysilicon -49 47 -49 47 3 _a0
rlabel polysilicon -49 71 -49 71 3 _a1
rlabel polysilicon -49 55 -49 55 3 _b0
rlabel polysilicon -49 63 -49 63 3 _b1
rlabel m2contact -12 87 -12 87 5 GND!
rlabel polysilicon -27 79 -27 79 1 _SReset!
rlabel metal2 -55 28 -55 28 1 _SReset!
rlabel metal2 0 37 0 43 1 _a0
rlabel metal2 0 49 0 55 3 _b0
rlabel metal2 0 73 0 79 3 _a1
rlabel space -61 25 -48 91 7 ^n
rlabel space -62 24 -25 92 7 ^n
rlabel space 28 29 53 91 3 ^p
rlabel metal2 0 61 0 67 3 _b1
rlabel metal2 -26 25 -26 31 3 ^n
rlabel metal1 26 123 26 123 5 Vdd!
rlabel metal1 -42 116 -42 116 1 GND!
rlabel metal1 50 112 50 112 6 Vdd!
rlabel polysilicon 59 106 59 106 7 _PReset!
rlabel metal2 66 124 66 124 5 _PReset!
rlabel metal1 52 120 52 120 1 Vdd!
rlabel metal2 48 76 48 76 1 _a1
rlabel metal2 48 64 48 64 1 _b1
rlabel metal2 48 52 48 52 1 _b0
<< end >>
