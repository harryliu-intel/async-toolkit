magic
tech scmos
timestamp 969938097
<< ndiffusion >>
rect -24 305 -8 306
rect -24 297 -8 302
rect -24 293 -8 294
<< pdiffusion >>
rect 8 305 24 307
rect 8 297 24 302
rect 8 293 24 294
<< ntransistor >>
rect -24 302 -8 305
rect -24 294 -8 297
<< ptransistor >>
rect 8 302 24 305
rect 8 294 24 297
<< polysilicon >>
rect -28 302 -24 305
rect -8 302 -4 305
rect 4 302 8 305
rect 24 302 28 305
rect -28 294 -24 297
rect -8 294 -4 297
rect 4 294 8 297
rect 24 294 28 297
<< ndcontact >>
rect -24 306 -8 314
rect -24 285 -8 293
<< pdcontact >>
rect 8 307 24 315
rect 8 285 24 293
<< psubstratepcontact >>
rect -41 293 -33 301
<< nsubstratencontact >>
rect 33 299 41 307
<< polycontact >>
rect -4 302 4 310
rect -4 289 4 297
<< metal1 >>
rect -24 306 -8 314
rect -21 303 -8 306
rect -41 293 -33 301
rect -4 302 4 309
rect 8 309 9 315
rect 21 309 41 315
rect 8 307 41 309
rect 33 299 41 307
rect -41 291 -8 293
rect -41 285 -21 291
rect -9 285 -8 291
rect -4 291 4 297
rect 8 293 21 297
rect 8 285 24 293
<< m2contact >>
rect -21 297 -8 303
rect -4 309 4 315
rect 9 309 21 315
rect 8 297 21 303
rect -21 285 -9 291
rect -4 285 4 291
<< metal2 >>
rect -27 309 4 315
rect -21 297 21 303
rect -4 285 27 291
<< m3contact >>
rect 9 309 21 315
rect -21 285 -9 291
<< metal3 >>
rect -21 282 -3 318
rect 3 282 21 318
<< labels >>
rlabel metal1 -12 310 -12 310 5 x
rlabel m2contact -12 289 -12 289 1 GND!
rlabel metal2 12 300 12 300 1 x
rlabel metal2 -12 300 -12 300 1 x
rlabel m2contact 12 310 12 310 5 Vdd!
rlabel metal1 12 289 12 289 1 x
rlabel polysilicon 25 295 25 295 7 a
rlabel polysilicon 25 303 25 303 7 b
rlabel polysilicon -25 295 -25 295 3 a
rlabel polysilicon -25 303 -25 303 3 b
rlabel metal2 26 288 26 288 7 a
rlabel metal2 25 285 27 291 7 ^p
rlabel metal2 -27 309 -25 315 3 ^n
rlabel metal2 -26 312 -26 312 3 b
rlabel metal1 -37 297 -37 297 3 GND!
rlabel metal1 37 303 37 303 7 Vdd!
rlabel space 23 284 42 316 3 ^p
rlabel space -42 284 -23 316 7 ^n
<< end >>
