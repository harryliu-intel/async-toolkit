//-----------------------------------------------------
// DUT IF signal connection
//-----------------------------------------------------
//assign `DUT_IF.XTAL_IN      = `HVL_TOP.xtal_25M_clk.clk;

//------------------------------------------------------
// FCSIG IF signal connection
//------------------------------------------------------
