magic
tech scmos
timestamp 970031125
<< ndiffusion >>
rect -43 50 -35 51
rect -21 52 -13 53
rect -43 46 -35 47
rect -21 44 -13 49
rect -43 37 -35 38
rect -21 36 -13 41
rect -21 32 -13 33
<< pdiffusion >>
rect 63 65 67 70
rect 55 64 67 65
rect 55 58 67 61
rect 55 49 71 50
rect 8 41 12 44
rect 8 32 12 37
rect 25 36 33 37
rect 55 45 71 46
rect 69 37 71 45
rect 55 36 71 37
rect 25 32 33 33
rect 55 32 71 33
<< ntransistor >>
rect -43 47 -35 50
rect -21 49 -13 52
rect -21 41 -13 44
rect -21 33 -13 36
<< ptransistor >>
rect 55 61 67 64
rect 55 46 71 49
rect 8 37 12 41
rect 25 33 33 36
rect 55 33 71 36
<< polysilicon >>
rect -33 50 -30 63
rect 35 61 55 64
rect 67 61 71 64
rect -11 56 21 57
rect -11 54 53 56
rect -11 52 -8 54
rect 18 53 53 54
rect -47 47 -43 50
rect -35 47 -30 50
rect -25 49 -21 52
rect -13 49 -8 52
rect 50 49 53 53
rect 50 46 55 49
rect 71 46 76 49
rect -25 41 -21 44
rect -13 41 -4 44
rect 4 37 8 41
rect 12 37 16 41
rect -26 33 -21 36
rect -13 33 -9 36
rect -26 27 -23 33
rect -47 24 -23 27
rect 37 36 40 37
rect 21 33 25 36
rect 33 33 40 36
rect 50 36 53 46
rect 73 44 76 46
rect 50 33 55 36
rect 71 33 76 36
<< ndcontact >>
rect -43 51 -35 59
rect -21 53 -13 61
rect -43 38 -35 46
rect -21 24 -13 32
<< pdcontact >>
rect 55 65 63 73
rect 8 44 16 52
rect 55 50 71 58
rect 25 37 33 45
rect 55 37 69 45
rect 8 24 16 32
rect 25 24 33 32
rect 55 24 71 32
<< psubstratepcontact >>
rect -43 29 -35 37
<< nsubstratencontact >>
rect 8 60 16 68
<< polycontact >>
rect -33 63 -25 71
rect 27 61 35 69
rect -55 24 -47 32
rect -4 36 4 44
rect 37 37 45 45
rect 73 36 81 44
<< metal1 >>
rect -33 67 -25 72
rect -33 63 -17 67
rect 8 66 16 68
rect 27 66 35 69
rect -21 61 -17 63
rect -43 55 -35 59
rect -21 56 -13 61
rect 42 65 63 72
rect -43 51 -27 55
rect -21 52 12 56
rect -43 32 -35 46
rect -31 44 -27 51
rect 8 44 16 52
rect 42 45 50 65
rect 55 50 71 58
rect -31 40 4 44
rect 25 40 33 45
rect -4 37 33 40
rect 37 37 69 45
rect 73 42 81 44
rect -4 36 29 37
rect -55 30 -47 32
rect -43 30 -13 32
rect 8 30 71 32
rect -43 24 -21 30
rect 21 24 71 30
<< m2contact >>
rect -33 72 -25 78
rect 42 72 63 78
rect 3 60 21 66
rect 27 60 35 66
rect 73 36 81 42
rect -55 24 -47 30
rect -21 24 -3 30
rect 3 24 21 30
<< metal2 >>
rect -33 72 63 78
rect 27 60 38 66
rect 0 36 81 42
rect -55 24 -27 30
<< m3contact >>
rect 3 60 21 66
rect -21 24 -3 30
rect 3 24 21 30
<< metal3 >>
rect -21 21 -3 81
rect 3 21 21 81
<< labels >>
rlabel pdcontact 29 28 29 28 1 Vdd!
rlabel m2contact 12 28 12 28 1 Vdd!
rlabel m2contact -17 28 -17 28 1 GND!
rlabel polysilicon -12 50 -12 50 1 a
rlabel polysilicon -12 34 -12 34 1 _SReset!
rlabel metal1 59 54 59 54 5 Vdd!
rlabel metal1 59 28 59 28 1 Vdd!
rlabel metal1 59 41 59 41 1 x
rlabel metal1 12 48 12 48 1 x
rlabel polysilicon 72 47 72 47 1 a
rlabel polysilicon 72 34 72 34 1 a
rlabel metal1 59 69 59 69 5 x
rlabel polysilicon 68 62 68 62 7 _PReset!
rlabel metal1 -17 56 -17 56 1 x
rlabel metal2 0 72 0 78 1 x
rlabel nsubstratencontact 12 64 12 64 1 Vdd!
rlabel ndcontact -39 42 -39 42 1 GND!
rlabel metal1 -39 33 -39 33 1 GND!
rlabel metal2 -51 27 -51 27 3 _SReset!
rlabel metal2 0 36 0 42 3 a
rlabel metal2 31 63 31 63 1 _PReset!
rlabel space 70 23 82 59 3 ^p
rlabel metal2 -29 75 -29 75 1 x
rlabel metal2 52 75 52 75 1 x
rlabel metal2 77 39 77 39 7 a
<< end >>
