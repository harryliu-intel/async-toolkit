///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit

//  Original version generated by ngen, but it didn't handle RX PPE interfaces with structs (yet)
//  so hand edits are required



///------------------------------------------------------------------------------
// -- Author       : Scott Greenfield
// -- Project Name : MBY 
// -- Description  : 
// ------------------------------------------------------------------- 

module igr_pre_post_wrap 
import mby_igr_pkg::*, shared_pkg::*;
(
//Input List
 input                             cclk, 
 input                             rst, // synchronized warm reset 
 input [4:0]                       i_free_ptr_valid,                         
 input [4:0][19:0]                 i_free_seg_ptr,                           
 input [4:0][3:0]                  i_free_sema,                              
 input igr_pkt_id_t [1:0]          i_return_id,                              
 input [1:0]                       i_return_id_valid,                        
 input shim_pb_data_t              i_shim_pb_data_p0[3:0],
 input shim_pb_data_t              i_shim_pb_data_p1[3:0],
 input shim_pb_data_t              i_shim_pb_data_p2[3:0],
 input shim_pb_data_t              i_shim_pb_data_p3[3:0],
 input shim_pb_md_t                i_shim_pb_md_p0[3:0],
 input shim_pb_md_t                i_shim_pb_md_p1[3:0],
 input shim_pb_md_t                i_shim_pb_md_p2[3:0],
 input shim_pb_md_t                i_shim_pb_md_p3[3:0],
 input logic [2:0]                 i_shim_pb_v_p0[3:0],  
 input logic [2:0]                 i_shim_pb_v_p1[3:0],  
 input logic [2:0]                 i_shim_pb_v_p2[3:0],  
 input logic [2:0]                 i_shim_pb_v_p3[3:0],

//Interface List
 input logic                       egr_igr_wreq_mim_wreq_valid, // Blasted Interface mim_wr_if.receive egr_igr_wreq
 input logic [20-1:0]              egr_igr_wreq_mim_wr_seg_ptr, 
 input logic [4-1:0]               egr_igr_wreq_mim_wr_sema, 
 input logic [2-1:0]               egr_igr_wreq_mim_wr_wd_sel, 
 input logic [13-1:0]              egr_igr_wreq_mim_wreq_id, 
 input logic [(8*64)-1:0]          egr_igr_wreq_mim_wr_data, 
 output logic [1-1:0]              egr_igr_wreq_mim_wreq_credits, 

 output igr_rx_ppe_tail_t          igr_rx_ppe_intf0_tail, // Blasted Interface igr_rx_ppe_if.igr igr_rx_ppe
 output igr_rx_ppe_head_t          igr_rx_ppe_intf0_head, 
 input logic                       igr_rx_ppe_intf0_ack, 
 output igr_rx_ppe_tail_t          igr_rx_ppe_intf1_tail, 
 output igr_rx_ppe_head_t          igr_rx_ppe_intf1_head, 
 input logic                       igr_rx_ppe_intf1_ack, 

 output logic                      mim_wreq_0_mim_wreq_valid, // Blasted Interface mim_wr_if.request mim_wreq_0
 output logic [20-1:0]             mim_wreq_0_mim_wr_seg_ptr, 
 output logic [4-1:0]              mim_wreq_0_mim_wr_sema, 
 output logic [2-1:0]              mim_wreq_0_mim_wr_wd_sel, 
 output logic [13-1:0]             mim_wreq_0_mim_wreq_id, 
 output logic [(8*64)-1:0]         mim_wreq_0_mim_wr_data, 
 input logic [1-1:0]               mim_wreq_0_mim_wreq_credits, 

 output logic                      mim_wreq_1_mim_wreq_valid, // Blasted Interface mim_wr_if.request mim_wreq_1
 output logic [20-1:0]             mim_wreq_1_mim_wr_seg_ptr, 
 output logic [4-1:0]              mim_wreq_1_mim_wr_sema, 
 output logic [2-1:0]              mim_wreq_1_mim_wr_wd_sel, 
 output logic [13-1:0]             mim_wreq_1_mim_wreq_id, 
 output logic [(8*64)-1:0]         mim_wreq_1_mim_wr_data, 
 input logic [1-1:0]               mim_wreq_1_mim_wreq_credits, 

 output logic                      mim_wreq_2_mim_wreq_valid, // Blasted Interface mim_wr_if.request mim_wreq_2
 output logic [20-1:0]             mim_wreq_2_mim_wr_seg_ptr, 
 output logic [4-1:0]              mim_wreq_2_mim_wr_sema, 
 output logic [2-1:0]              mim_wreq_2_mim_wr_wd_sel, 
 output logic [13-1:0]             mim_wreq_2_mim_wreq_id, 
 output logic [(8*64)-1:0]         mim_wreq_2_mim_wr_data, 
 input logic [1-1:0]               mim_wreq_2_mim_wreq_credits, 

 output logic                      mim_wreq_3_mim_wreq_valid, // Blasted Interface mim_wr_if.request mim_wreq_3
 output logic [20-1:0]             mim_wreq_3_mim_wr_seg_ptr, 
 output logic [4-1:0]              mim_wreq_3_mim_wr_sema, 
 output logic [2-1:0]              mim_wreq_3_mim_wr_wd_sel, 
 output logic [13-1:0]             mim_wreq_3_mim_wreq_id, 
 output logic [(8*64)-1:0]         mim_wreq_3_mim_wr_data, 
 input logic [1-1:0]               mim_wreq_3_mim_wreq_credits, 

 output logic                      mim_wreq_4_mim_wreq_valid, // Blasted Interface mim_wr_if.request mim_wreq_4
 output logic [20-1:0]             mim_wreq_4_mim_wr_seg_ptr, 
 output logic [4-1:0]              mim_wreq_4_mim_wr_sema, 
 output logic [2-1:0]              mim_wreq_4_mim_wr_wd_sel, 
 output logic [13-1:0]             mim_wreq_4_mim_wreq_id, 
 output logic [(8*64)-1:0]         mim_wreq_4_mim_wr_data, 
 input logic [1-1:0]               mim_wreq_4_mim_wreq_credits, 

 output logic                      mim_wreq_5_mim_wreq_valid, // Blasted Interface mim_wr_if.request mim_wreq_5
 output logic [20-1:0]             mim_wreq_5_mim_wr_seg_ptr, 
 output logic [4-1:0]              mim_wreq_5_mim_wr_sema, 
 output logic [2-1:0]              mim_wreq_5_mim_wr_wd_sel, 
 output logic [13-1:0]             mim_wreq_5_mim_wreq_id, 
 output logic [(8*64)-1:0]         mim_wreq_5_mim_wr_data, 
 input logic [1-1:0]               mim_wreq_5_mim_wreq_credits, 

 input rx_ppe_igr_t                rx_ppe_igr_intf0, // Blasted Interface rx_ppe_igr_if.igr rx_ppe_igr
 input rx_ppe_igr_t                rx_ppe_igr_intf1, 

//Output List
 output [W_SEG_PTR-1:0][1:0]       o_drop_seg_ptr, //[19:0] 
 output [1:0]                      o_drop_seg_valid, 
 output [W_SEMA-1:0][1:0]          o_drop_sema, 
 output [4:0]                      o_free_ptr_req,
 output [7:0]                      o_port_id, // FIXME -- what is this for?  ring_tag_t also has src & dst ports 
 output [95:0]                     o_post_ppe_tag_at_rate0, 
 output [95:0]                     o_post_ppe_tag_at_rate1, 
 output [95:0]                     o_post_ppe_tag_set_aside0, 
 output [95:0]                     o_post_ppe_tag_set_aside1                 
);
// collage-pragma translate_off

pre_post_ppe_partial_data_if     pdata_lpp0_fpp();
pre_post_ppe_partial_data_if     pdata_lpp1();
pre_post_ppe_sop_if              sop_mdata_lpp0_fpp();
pre_post_ppe_sop_if              sop_mdata_lpp1();
pre_post_ppe_tag_info_if         tag_info_epl[NUM_EPLS-1:0]();
pre_post_ppe_tag_info_if         tag_info_vp();
pre_post_ppe_wr_data_if          wr_data_0();
pre_post_ppe_wr_data_if          wr_data_1();
pre_post_ppe_wr_data_if          wr_data_2();
mim_wr_if egr_igr_wreq();
// Blasted Wires for mim_wr_if receive egr_igr_wreq;
    assign egr_igr_wreq.mim_wreq_valid = egr_igr_wreq_mim_wreq_valid;
    assign egr_igr_wreq.mim_wr_seg_ptr = egr_igr_wreq_mim_wr_seg_ptr;
    assign egr_igr_wreq.mim_wr_sema = egr_igr_wreq_mim_wr_sema;
    assign egr_igr_wreq.mim_wr_wd_sel = egr_igr_wreq_mim_wr_wd_sel;
    assign egr_igr_wreq.mim_wreq_id = egr_igr_wreq_mim_wreq_id;
    assign egr_igr_wreq.mim_wr_data = egr_igr_wreq_mim_wr_data;
    assign egr_igr_wreq_mim_wreq_credits = egr_igr_wreq.mim_wreq_credits;

igr_rx_ppe_if igr_rx_ppe();
// Blasted Wires for igr_rx_ppe_if igr igr_rx_ppe;
    assign igr_rx_ppe_intf0_tail = igr_rx_ppe.intf0_tail;
    assign igr_rx_ppe_intf0_head = igr_rx_ppe.intf0_head;
    assign igr_rx_ppe.intf0_ack = igr_rx_ppe_intf0_ack;
    assign igr_rx_ppe_intf1_tail = igr_rx_ppe.intf1_tail;
    assign igr_rx_ppe_intf1_head = igr_rx_ppe.intf1_head;
    assign igr_rx_ppe.intf1_ack = igr_rx_ppe_intf1_ack;

mim_wr_if mim_wreq_0();
// Blasted Wires for mim_wr_if request mim_wreq_0;
    assign mim_wreq_0_mim_wreq_valid = mim_wreq_0.mim_wreq_valid;
    assign mim_wreq_0_mim_wr_seg_ptr = mim_wreq_0.mim_wr_seg_ptr;
    assign mim_wreq_0_mim_wr_sema = mim_wreq_0.mim_wr_sema;
    assign mim_wreq_0_mim_wr_wd_sel = mim_wreq_0.mim_wr_wd_sel;
    assign mim_wreq_0_mim_wreq_id = mim_wreq_0.mim_wreq_id;
    assign mim_wreq_0_mim_wr_data = mim_wreq_0.mim_wr_data;
    assign mim_wreq_0.mim_wreq_credits = mim_wreq_0_mim_wreq_credits;

mim_wr_if mim_wreq_1();
// Blasted Wires for mim_wr_if request mim_wreq_1;
    assign mim_wreq_1_mim_wreq_valid = mim_wreq_1.mim_wreq_valid;
    assign mim_wreq_1_mim_wr_seg_ptr = mim_wreq_1.mim_wr_seg_ptr;
    assign mim_wreq_1_mim_wr_sema = mim_wreq_1.mim_wr_sema;
    assign mim_wreq_1_mim_wr_wd_sel = mim_wreq_1.mim_wr_wd_sel;
    assign mim_wreq_1_mim_wreq_id = mim_wreq_1.mim_wreq_id;
    assign mim_wreq_1_mim_wr_data = mim_wreq_1.mim_wr_data;
    assign mim_wreq_1.mim_wreq_credits = mim_wreq_1_mim_wreq_credits;

mim_wr_if mim_wreq_2();
// Blasted Wires for mim_wr_if request mim_wreq_2;
    assign mim_wreq_2_mim_wreq_valid = mim_wreq_2.mim_wreq_valid;
    assign mim_wreq_2_mim_wr_seg_ptr = mim_wreq_2.mim_wr_seg_ptr;
    assign mim_wreq_2_mim_wr_sema = mim_wreq_2.mim_wr_sema;
    assign mim_wreq_2_mim_wr_wd_sel = mim_wreq_2.mim_wr_wd_sel;
    assign mim_wreq_2_mim_wreq_id = mim_wreq_2.mim_wreq_id;
    assign mim_wreq_2_mim_wr_data = mim_wreq_2.mim_wr_data;
    assign mim_wreq_2.mim_wreq_credits = mim_wreq_2_mim_wreq_credits;

mim_wr_if mim_wreq_3();
// Blasted Wires for mim_wr_if request mim_wreq_3;
    assign mim_wreq_3_mim_wreq_valid = mim_wreq_3.mim_wreq_valid;
    assign mim_wreq_3_mim_wr_seg_ptr = mim_wreq_3.mim_wr_seg_ptr;
    assign mim_wreq_3_mim_wr_sema = mim_wreq_3.mim_wr_sema;
    assign mim_wreq_3_mim_wr_wd_sel = mim_wreq_3.mim_wr_wd_sel;
    assign mim_wreq_3_mim_wreq_id = mim_wreq_3.mim_wreq_id;
    assign mim_wreq_3_mim_wr_data = mim_wreq_3.mim_wr_data;
    assign mim_wreq_3.mim_wreq_credits = mim_wreq_3_mim_wreq_credits;

mim_wr_if mim_wreq_4();
// Blasted Wires for mim_wr_if request mim_wreq_4;
    assign mim_wreq_4_mim_wreq_valid = mim_wreq_4.mim_wreq_valid;
    assign mim_wreq_4_mim_wr_seg_ptr = mim_wreq_4.mim_wr_seg_ptr;
    assign mim_wreq_4_mim_wr_sema = mim_wreq_4.mim_wr_sema;
    assign mim_wreq_4_mim_wr_wd_sel = mim_wreq_4.mim_wr_wd_sel;
    assign mim_wreq_4_mim_wreq_id = mim_wreq_4.mim_wreq_id;
    assign mim_wreq_4_mim_wr_data = mim_wreq_4.mim_wr_data;
    assign mim_wreq_4.mim_wreq_credits = mim_wreq_4_mim_wreq_credits;

mim_wr_if mim_wreq_5();
// Blasted Wires for mim_wr_if request mim_wreq_5;
    assign mim_wreq_5_mim_wreq_valid = mim_wreq_5.mim_wreq_valid;
    assign mim_wreq_5_mim_wr_seg_ptr = mim_wreq_5.mim_wr_seg_ptr;
    assign mim_wreq_5_mim_wr_sema = mim_wreq_5.mim_wr_sema;
    assign mim_wreq_5_mim_wr_wd_sel = mim_wreq_5.mim_wr_wd_sel;
    assign mim_wreq_5_mim_wreq_id = mim_wreq_5.mim_wreq_id;
    assign mim_wreq_5_mim_wr_data = mim_wreq_5.mim_wr_data;
    assign mim_wreq_5.mim_wreq_credits = mim_wreq_5_mim_wreq_credits;

rx_ppe_igr_if rx_ppe_igr();
// Blasted Wires for rx_ppe_igr_if igr rx_ppe_igr;
    assign rx_ppe_igr.intf0 = rx_ppe_igr_t'(rx_ppe_igr_intf0);
    assign rx_ppe_igr.intf1 = rx_ppe_igr_t'(rx_ppe_igr_intf1);



// module mby_igr_pre_ppe    from mby_igr_pre_ppe using pre_ppe.map 
mby_igr_pre_ppe    mby_igr_pre_ppe(
/* input  logic                               */ .cclk               (cclk),                            
/* input  logic                               */ .rst                (rst),                             // synchronized warm reset 
/* Interface igr_rx_ppe_if.igr                */ .igr_rx_ppe         (igr_rx_ppe),                      
/* input  logic                         [3:0] */ .i_shim_pb_data_p0  (i_shim_pb_data_p0),               
/* input  logic                         [3:0] */ .i_shim_pb_data_p1  (i_shim_pb_data_p1),               
/* input  logic                         [3:0] */ .i_shim_pb_data_p2  (i_shim_pb_data_p2),               
/* input  logic                         [3:0] */ .i_shim_pb_data_p3  (i_shim_pb_data_p3),               
/* input  logic                  [3:0][173:0] */ .i_shim_pb_md_p0    (i_shim_pb_md_p0),                 
/* input  logic                  [3:0][173:0] */ .i_shim_pb_md_p1    (i_shim_pb_md_p1),                 
/* input  logic                  [3:0][173:0] */ .i_shim_pb_md_p2    (i_shim_pb_md_p2),                 
/* input  logic                  [3:0][173:0] */ .i_shim_pb_md_p3    (i_shim_pb_md_p3),                 
/* input  logic                    [2:0][3:0] */ .i_shim_pb_v_p0     (i_shim_pb_v_p0),                  
/* input  logic                    [2:0][3:0] */ .i_shim_pb_v_p1     (i_shim_pb_v_p1),                  
/* input  logic                    [2:0][3:0] */ .i_shim_pb_v_p2     (i_shim_pb_v_p2),                  
/* input  logic                    [2:0][3:0] */ .i_shim_pb_v_p3     (i_shim_pb_v_p3),                  
/* input  logic                         [4:0] */ .i_free_ptr_valid   (i_free_ptr_valid),              
/* output logic                         [4:0] */ .o_free_ptr_req     (o_free_ptr_req),                
/* input  logic                   [4:0][19:0] */ .i_free_seg_ptr     (i_free_seg_ptr),                
/* input  logic                    [4:0][3:0] */ .i_free_sema        (i_free_sema),                   
/* input  logic                    [1:0][0:0] */ .i_return_id        (i_return_id),                   
/* input  logic                         [1:0] */ .i_return_id_valid  (i_return_id_valid),             
/* Interface pre_post_ppe_partial_data_if.src */ .pdata_lpp0_fpp     (pdata_lpp0_fpp),                
/* Interface pre_post_ppe_partial_data_if.src */ .pdata_lpp1         (pdata_lpp1),                    
/* Interface pre_post_ppe_sop_if.src          */ .sop_mdata_lpp0_fpp (sop_mdata_lpp0_fpp),            
/* Interface pre_post_ppe_sop_if.src          */ .sop_mdata_lpp1     (sop_mdata_lpp1),                
/* Interface pre_post_ppe_tag_info_if.src     */ .tag_info_epl       (tag_info_epl),                 
/* Interface pre_post_ppe_tag_info_if.src     */ .tag_info_vp        (tag_info_vp),                   
/* Interface pre_post_ppe_wr_data_if.src      */ .wr_data_0          (wr_data_0),                     
/* Interface pre_post_ppe_wr_data_if.src      */ .wr_data_1          (wr_data_1),                     
/* Interface pre_post_ppe_wr_data_if.src      */ .wr_data_2          (wr_data_2));                     
// End of module mby_igr_pre_ppe from mby_igr_pre_ppe


// module mby_igr_post_ppe    from mby_igr_post_ppe using post_ppe.map 
mby_igr_post_ppe    mby_igr_post_ppe(
/* input  logic                               */ .cclk                      (cclk),                                   
/* input  logic                               */ .rst                       (rst),                                    // synchronized warm reset 
/* Interface rx_ppe_igr_if.igr                */ .rx_ppe_igr                (rx_ppe_igr),                             
/* Interface mim_wr_if.receive                */ .egr_igr_wreq              (egr_igr_wreq),                           
/* Interface mim_wr_if.request                */ .mim_wreq_0                (mim_wreq_0),                             
/* Interface mim_wr_if.request                */ .mim_wreq_1                (mim_wreq_1),                             
/* Interface mim_wr_if.request                */ .mim_wreq_2                (mim_wreq_2),                             
/* Interface mim_wr_if.request                */ .mim_wreq_3                (mim_wreq_3),                             
/* Interface mim_wr_if.request                */ .mim_wreq_4                (mim_wreq_4),                             
/* Interface mim_wr_if.request                */ .mim_wreq_5                (mim_wreq_5),                             
/* Interface pre_post_ppe_partial_data_if.src */ .pdata_lpp0_fpp            (pdata_lpp0_fpp),                         
/* Interface pre_post_ppe_partial_data_if.src */ .pdata_lpp1                (pdata_lpp1),                             
/* Interface pre_post_ppe_sop_if.src          */ .sop_mdata_lpp0_fpp        (sop_mdata_lpp0_fpp),                     
/* Interface pre_post_ppe_sop_if.src          */ .sop_mdata_lpp1            (sop_mdata_lpp1),                         
/* Interface pre_post_ppe_tag_info_if.src     */ .tag_info_epl              (tag_info_epl),                          
/* Interface pre_post_ppe_tag_info_if.src     */ .tag_info_vp               (tag_info_vp),                            
/* Interface pre_post_ppe_wr_data_if.src      */ .wr_data_0                 (wr_data_0),                              
/* Interface pre_post_ppe_wr_data_if.src      */ .wr_data_1                 (wr_data_1),                              
/* Interface pre_post_ppe_wr_data_if.src      */ .wr_data_2                 (wr_data_2),                              
/* output logic                        [95:0] */ .o_post_ppe_tag_at_rate0   (o_post_ppe_tag_at_rate0),                
/* output logic                        [95:0] */ .o_post_ppe_tag_at_rate1   (o_post_ppe_tag_at_rate1),                
/* output logic                        [95:0] */ .o_post_ppe_tag_set_aside0 (o_post_ppe_tag_set_aside0),              
/* output logic                        [95:0] */ .o_post_ppe_tag_set_aside1 (o_post_ppe_tag_set_aside1),              
/* output logic                         [7:0] */ .o_port_id                 (o_port_id),                              // FIXME -- what is this for?  ring_tag_t also has src & dst ports 
/* output logic                         [1:0] */ .o_drop_seg_valid          (o_drop_seg_valid),                       
/* output logic          [W_SEG_PTR-1:0][1:0] */ .o_drop_seg_ptr            (o_drop_seg_ptr),     //[19:0] 
/* output logic             [W_SEMA-1:0][1:0] */ .o_drop_sema               (o_drop_sema) );           
// End of module mby_igr_post_ppe from mby_igr_post_ppe

// collage-pragma translate_on

endmodule // igr_pre_post_wrap
