// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

//-----------------------------------------------------------------------------
// Title         : Ingress hard reset sequence
// Project       : Madison Bay
//-----------------------------------------------------------------------------
// File          : mby_igr_hard_reset_seq.sv
// Author        : jose.j.godinez.carrillo  <jjgodine@ichips.intel.com>
// Created       : 22.08.2018
// Last modified : 22.08.2018
//-----------------------------------------------------------------------------
// Description :
//
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by Intel Corporation This model is the confidential and
// proprietary property of Intel Corporation and the possession or use of this
// file requires a written license from Intel Corporation.
//-----------------------------------------------------------------------------
// Modification history :
// 22.08.2018 : created
//-----------------------------------------------------------------------------

//-----------------------------------------------------------------------------
// Class: mby_igr_hard_reset_seq
//-----------------------------------------------------------------------------
class mby_igr_hard_reset_seq extends mby_igr_extended_base_seq;

   `uvm_object_utils(mby_igr_hard_reset_seq)

   //--------------------------------------------------------------------------
   // Task: body()
   //--------------------------------------------------------------------------
   task body();
      virtual mby_igr_env_if env_if;
      mby_igr_env ingress_env_ptr;
      uvm_event ingress_fusepull_comp_e;
      uvm_event_pool    ingress_epool;

      uvm_report_warning (get_name(), "INTEG - INGRESS_hard_reset should be IMP ");

      assert($cast(ingress_env_ptr, mby_igr_env::get_igr_env()))
      else begin
         `uvm_error(get_name(), $sformatf("Unable to get handle to mby_igr_env."));
      end

      //Pointer to env IF
      env_if = ingress_env_ptr.ingress_if;
      //pointer to event pool and fuse event
      ingress_epool = ingress_epool.get_global_pool();
      ingress_fusepull_comp_e = ingress_epool.get("INGRESS_DETECT_FUSEPULL_COMP_SB_MSG");

      //Reset and power up flow
      env_if.power_good_reset = 0;
      env_if.reset = 0;

      //power good
      #1;
      env_if.power_good_reset = 1;

      ingress_fusepull_comp_e.wait_trigger();

      //Primary interface
      repeat (10) begin
         @(posedge env_if.clock);
      end
      env_if.reset = 1;

   endtask : body

endclass : mby_igr_hard_reset_seq
