magic
tech scmos
timestamp 988943070
<< nselect >>
rect -59 91 0 146
<< pselect >>
rect 0 89 46 154
<< ndiffusion >>
rect -53 132 -33 133
rect -28 132 -8 133
rect -53 124 -33 129
rect -28 124 -8 129
rect -53 116 -33 121
rect -28 116 -8 121
rect -53 108 -33 113
rect -28 108 -8 113
rect -53 104 -33 105
rect -28 104 -8 105
<< pdiffusion >>
rect 8 142 40 143
rect 8 138 40 139
rect 8 129 40 130
rect 8 125 40 126
rect 28 117 40 125
rect 8 116 40 117
rect 8 112 40 113
rect 8 103 40 104
rect 8 99 40 100
<< ntransistor >>
rect -53 129 -33 132
rect -28 129 -8 132
rect -53 121 -33 124
rect -28 121 -8 124
rect -53 113 -33 116
rect -28 113 -8 116
rect -53 105 -33 108
rect -28 105 -8 108
<< ptransistor >>
rect 8 139 40 142
rect 8 126 40 129
rect 8 113 40 116
rect 8 100 40 103
<< polysilicon >>
rect -5 139 8 142
rect 40 139 44 142
rect -5 132 -2 139
rect -57 129 -53 132
rect -33 129 -28 132
rect -8 129 -2 132
rect 3 126 8 129
rect 40 126 44 129
rect 3 124 6 126
rect -57 121 -53 124
rect -33 121 -28 124
rect -8 121 6 124
rect -57 113 -53 116
rect -33 113 -28 116
rect -8 113 8 116
rect 40 113 44 116
rect -57 105 -53 108
rect -33 105 -28 108
rect -8 105 2 108
rect -1 103 2 105
rect -1 100 8 103
rect 40 100 44 103
<< ndcontact >>
rect -53 133 -33 141
rect -28 133 -8 141
rect -53 96 -33 104
rect -28 96 -8 104
<< pdcontact >>
rect 8 143 40 151
rect 8 130 40 138
rect 8 117 28 125
rect 8 104 40 112
rect 8 91 40 99
<< metal1 >>
rect 8 143 40 151
rect -53 133 -33 141
rect -28 133 -8 141
rect -41 125 -33 133
rect 8 130 40 138
rect -41 117 28 125
rect -16 104 -8 117
rect 32 112 40 130
rect 8 104 40 112
rect -53 96 -33 104
rect -28 96 -8 104
rect 8 91 40 99
<< labels >>
rlabel space -61 91 -28 146 7 ^n
rlabel space -60 91 -53 146 7 ^n
rlabel space 28 89 47 154 3 ^p
rlabel metal1 -41 117 28 125 1 x|pin|s|2
rlabel metal1 -41 117 -33 141 1 x|pin|s|2
rlabel metal1 -53 133 -33 141 1 x|pin|s|2
rlabel metal1 -28 96 -8 104 1 x|pin|s|2
rlabel metal1 -16 96 -8 125 1 x|pin|s|2
rlabel polysilicon 40 100 44 103 1 _a0|pin|w|3|poly
rlabel polysilicon -1 100 3 103 1 _a0|pin|w|3|poly
rlabel polysilicon -57 105 -53 108 1 _a0|pin|w|3|poly
rlabel polysilicon -57 113 -53 116 1 _b0|pin|w|4|poly
rlabel polysilicon 40 113 44 116 1 _b0|pin|w|4|poly
rlabel polysilicon 40 126 44 129 1 _b1|pin|w|5|poly
rlabel polysilicon -57 121 -53 124 1 _b1|pin|w|5|poly
rlabel polysilicon -57 129 -53 132 1 _a1|pin|w|6|poly
rlabel polysilicon -2 139 2 142 1 _a1|pin|w|6|poly
rlabel polysilicon 40 139 44 142 1 _a1|pin|w|6|poly
rlabel metal1 8 143 40 151 1 Vdd!|pin|s|1
rlabel metal1 8 91 40 99 1 Vdd!|pin|s|0
rlabel metal1 -28 133 -8 141 1 GND!|pin|s|1
rlabel metal1 -53 96 -33 104 1 GND!|pin|s|0
<< end >>
