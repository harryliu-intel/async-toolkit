// File: mby_test_pack.sv

package mby_test_pack;
    import sla_pkg::*;
    import ovm_pkg::*;
    import mby_env_pkg::*;
  
    `include "ovm_macros.svh"
    `include "sla_macros.svh"

    `include "mby_base_test.svh"
    `include "mby_alive_test/mby_alive_test.svh"
endpackage
