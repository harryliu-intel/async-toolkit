//-----------------------------------------------------------------------------
// Title         : Ingress config object
// Project       : Madison Bay
//-----------------------------------------------------------------------------
// File          : mby_egr_env_cfg.svh
// Author        : jose.j.godinez.carrillo  <jjgodine@ichips.intel.com>
// Created       : 21.08.2018
// Last modified : 21.08.2018
//-----------------------------------------------------------------------------
// Description :
// This is the configuration object to control the mby_egr env.
// This Class contain all the switches to control the ENV setting.
// 
// By default it contains Saola config object:
// 
// checkers_enabled - default 1
// monitors_enabled - default 1
// trackers_enabled - default 1
// coverage_enabled - default 1
// 
// By default Saola will be build this object unless Upper env 
// or a test override it using set_config ...
//
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by Intel Corporation This model is the confidential and
// proprietary property of Intel Corporation and the possession or use of this
// file requires a written license from Intel Corporation.
//-----------------------------------------------------------------------------
// Modification history :
// 21.08.2018 : created
//-----------------------------------------------------------------------------

//-----------------------------------------------------------------------------
// Class: mby_egr_env_cfg
//-----------------------------------------------------------------------------
class mby_egr_env_cfg extends uvm_object;

    string egress_primary_access  = "primary";
    string egress_sideband_access = "sideband";
    bit    egress_chassis_rst_verbose_dbg;
    bit    egress_has_reset_pkg = 0;
    mby_smm_bfm_cfg smm_bfm_cfg;

   `uvm_object_utils_begin(mby_egr_env_cfg)
      `uvm_field_string(egress_primary_access,          UVM_ALL_ON)
      `uvm_field_string(egress_sideband_access,         UVM_ALL_ON)
      `uvm_field_string(egress_chassis_rst_verbose_dbg, UVM_ALL_ON)
   `uvm_object_utils_end

   //--------------------------------------------------------------------------
   // Function: new
   //--------------------------------------------------------------------------
   function new (string name = "mby_egr_env_cfg");
      super.new(name);
   endfunction : new

   //function void build_phase(uvm_phase phase);
   //   super.build_phase(phase);
   //   smm_bfm_cfg = new("smm_bfm_cfg");
   //endfunction : build_phase

endclass : mby_egr_env_cfg
