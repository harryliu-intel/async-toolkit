///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_entropy_map_pkg.vh                                 
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_ENTROPY_MAP_PKG_VH
`define MBY_PPE_ENTROPY_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_entropy_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_entropy_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_entropy_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_entropy_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [31:0] KEY_MASK8;  // RW
} ENTROPY_HASH_CFG0_t;

localparam ENTROPY_HASH_CFG0_REG_STRIDE = 48'h8;
localparam ENTROPY_HASH_CFG0_REG_ENTRIES = 64;
localparam ENTROPY_HASH_CFG0_REGFILE_STRIDE = 48'h200;
localparam ENTROPY_HASH_CFG0_REGFILE_ENTRIES = 3;
localparam ENTROPY_HASH_CFG0_CR_ADDR = 48'h0;
localparam ENTROPY_HASH_CFG0_SIZE = 64;
localparam ENTROPY_HASH_CFG0_KEY_MASK8_LO = 0;
localparam ENTROPY_HASH_CFG0_KEY_MASK8_HI = 31;
localparam ENTROPY_HASH_CFG0_KEY_MASK8_RESET = 32'h0;
localparam ENTROPY_HASH_CFG0_USEMASK = 64'hFFFFFFFF;
localparam ENTROPY_HASH_CFG0_RO_MASK = 64'h0;
localparam ENTROPY_HASH_CFG0_WO_MASK = 64'h0;
localparam ENTROPY_HASH_CFG0_RESET = 64'h0;

typedef struct packed {
    logic  [8:0] reserved0;  // RSVD
    logic  [0:0] SYMMETRIC;  // RW
    logic  [1:0] SYM_PROFILE;  // RW
    logic  [3:0] KEY_MASK_PROFILE;  // RW
    logic [15:0] KEY_MASK32;  // RW
    logic [31:0] KEY_MASK16;  // RW
} ENTROPY_HASH_CFG1_t;

localparam ENTROPY_HASH_CFG1_REG_STRIDE = 48'h8;
localparam ENTROPY_HASH_CFG1_REG_ENTRIES = 64;
localparam ENTROPY_HASH_CFG1_REGFILE_STRIDE = 48'h200;
localparam ENTROPY_HASH_CFG1_REGFILE_ENTRIES = 3;
localparam ENTROPY_HASH_CFG1_CR_ADDR = 48'h800;
localparam ENTROPY_HASH_CFG1_SIZE = 64;
localparam ENTROPY_HASH_CFG1_SYMMETRIC_LO = 54;
localparam ENTROPY_HASH_CFG1_SYMMETRIC_HI = 54;
localparam ENTROPY_HASH_CFG1_SYMMETRIC_RESET = 1'h0;
localparam ENTROPY_HASH_CFG1_SYM_PROFILE_LO = 52;
localparam ENTROPY_HASH_CFG1_SYM_PROFILE_HI = 53;
localparam ENTROPY_HASH_CFG1_SYM_PROFILE_RESET = 2'h0;
localparam ENTROPY_HASH_CFG1_KEY_MASK_PROFILE_LO = 48;
localparam ENTROPY_HASH_CFG1_KEY_MASK_PROFILE_HI = 51;
localparam ENTROPY_HASH_CFG1_KEY_MASK_PROFILE_RESET = 4'h0;
localparam ENTROPY_HASH_CFG1_KEY_MASK32_LO = 32;
localparam ENTROPY_HASH_CFG1_KEY_MASK32_HI = 47;
localparam ENTROPY_HASH_CFG1_KEY_MASK32_RESET = 16'h0;
localparam ENTROPY_HASH_CFG1_KEY_MASK16_LO = 0;
localparam ENTROPY_HASH_CFG1_KEY_MASK16_HI = 31;
localparam ENTROPY_HASH_CFG1_KEY_MASK16_RESET = 32'h0;
localparam ENTROPY_HASH_CFG1_USEMASK = 64'h7FFFFFFFFFFFFF;
localparam ENTROPY_HASH_CFG1_RO_MASK = 64'h0;
localparam ENTROPY_HASH_CFG1_WO_MASK = 64'h0;
localparam ENTROPY_HASH_CFG1_RESET = 64'h0;

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic [11:0] BYTE_DEFAULTS;  // RW
    logic  [5:0] HASH_START;  // RW
    logic  [5:0] HASH_SIZE;  // RW
} ENTROPY_META_CFG_t;

localparam ENTROPY_META_CFG_REG_STRIDE = 48'h8;
localparam ENTROPY_META_CFG_REG_ENTRIES = 64;
localparam ENTROPY_META_CFG_CR_ADDR = 48'hE00;
localparam ENTROPY_META_CFG_SIZE = 64;
localparam ENTROPY_META_CFG_BYTE_DEFAULTS_LO = 12;
localparam ENTROPY_META_CFG_BYTE_DEFAULTS_HI = 23;
localparam ENTROPY_META_CFG_BYTE_DEFAULTS_RESET = 12'h0;
localparam ENTROPY_META_CFG_HASH_START_LO = 6;
localparam ENTROPY_META_CFG_HASH_START_HI = 11;
localparam ENTROPY_META_CFG_HASH_START_RESET = 6'h0;
localparam ENTROPY_META_CFG_HASH_SIZE_LO = 0;
localparam ENTROPY_META_CFG_HASH_SIZE_HI = 5;
localparam ENTROPY_META_CFG_HASH_SIZE_RESET = 6'h0;
localparam ENTROPY_META_CFG_USEMASK = 64'hFFFFFF;
localparam ENTROPY_META_CFG_RO_MASK = 64'h0;
localparam ENTROPY_META_CFG_WO_MASK = 64'h0;
localparam ENTROPY_META_CFG_RESET = 64'h0;

typedef struct packed {
    logic  [3:0] reserved0;  // RSVD
    logic [59:0] KEY_PAIRS;  // RW
} ENTROPY_HASH_SYM8_t;

localparam ENTROPY_HASH_SYM8_REG_STRIDE = 48'h8;
localparam ENTROPY_HASH_SYM8_REG_ENTRIES = 4;
localparam ENTROPY_HASH_SYM8_REGFILE_STRIDE = 48'h20;
localparam ENTROPY_HASH_SYM8_REGFILE_ENTRIES = 3;
localparam ENTROPY_HASH_SYM8_CR_ADDR = 48'h1000;
localparam ENTROPY_HASH_SYM8_SIZE = 64;
localparam ENTROPY_HASH_SYM8_KEY_PAIRS_LO = 0;
localparam ENTROPY_HASH_SYM8_KEY_PAIRS_HI = 59;
localparam ENTROPY_HASH_SYM8_KEY_PAIRS_RESET = 60'h0;
localparam ENTROPY_HASH_SYM8_USEMASK = 64'hFFFFFFFFFFFFFFF;
localparam ENTROPY_HASH_SYM8_RO_MASK = 64'h0;
localparam ENTROPY_HASH_SYM8_WO_MASK = 64'h0;
localparam ENTROPY_HASH_SYM8_RESET = 64'h0;

typedef struct packed {
    logic  [3:0] reserved0;  // RSVD
    logic [59:0] KEY_PAIRS;  // RW
} ENTROPY_HASH_SYM16_t;

localparam ENTROPY_HASH_SYM16_REG_STRIDE = 48'h8;
localparam ENTROPY_HASH_SYM16_REG_ENTRIES = 4;
localparam ENTROPY_HASH_SYM16_REGFILE_STRIDE = 48'h20;
localparam ENTROPY_HASH_SYM16_REGFILE_ENTRIES = 3;
localparam ENTROPY_HASH_SYM16_CR_ADDR = 48'h1080;
localparam ENTROPY_HASH_SYM16_SIZE = 64;
localparam ENTROPY_HASH_SYM16_KEY_PAIRS_LO = 0;
localparam ENTROPY_HASH_SYM16_KEY_PAIRS_HI = 59;
localparam ENTROPY_HASH_SYM16_KEY_PAIRS_RESET = 60'h0;
localparam ENTROPY_HASH_SYM16_USEMASK = 64'hFFFFFFFFFFFFFFF;
localparam ENTROPY_HASH_SYM16_RO_MASK = 64'h0;
localparam ENTROPY_HASH_SYM16_WO_MASK = 64'h0;
localparam ENTROPY_HASH_SYM16_RESET = 64'h0;

typedef struct packed {
    logic [63:0] KEY_PAIRS;  // RW
} ENTROPY_HASH_SYM32_t;

localparam ENTROPY_HASH_SYM32_REG_STRIDE = 48'h8;
localparam ENTROPY_HASH_SYM32_REG_ENTRIES = 4;
localparam ENTROPY_HASH_SYM32_REGFILE_STRIDE = 48'h20;
localparam ENTROPY_HASH_SYM32_REGFILE_ENTRIES = 3;
localparam ENTROPY_HASH_SYM32_CR_ADDR = 48'h1100;
localparam ENTROPY_HASH_SYM32_SIZE = 64;
localparam ENTROPY_HASH_SYM32_KEY_PAIRS_LO = 0;
localparam ENTROPY_HASH_SYM32_KEY_PAIRS_HI = 63;
localparam ENTROPY_HASH_SYM32_KEY_PAIRS_RESET = 64'h0;
localparam ENTROPY_HASH_SYM32_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam ENTROPY_HASH_SYM32_RO_MASK = 64'h0;
localparam ENTROPY_HASH_SYM32_WO_MASK = 64'h0;
localparam ENTROPY_HASH_SYM32_RESET = 64'h0;

typedef struct packed {
    logic [63:0] MASK;  // RW
} ENTROPY_HASH_KEY_MASK_t;

localparam ENTROPY_HASH_KEY_MASK_REG_STRIDE = 48'h8;
localparam ENTROPY_HASH_KEY_MASK_REG_ENTRIES = 128;
localparam ENTROPY_HASH_KEY_MASK_REGFILE_STRIDE = 48'h400;
localparam ENTROPY_HASH_KEY_MASK_REGFILE_ENTRIES = 3;
localparam ENTROPY_HASH_KEY_MASK_CR_ADDR = 48'h2000;
localparam ENTROPY_HASH_KEY_MASK_SIZE = 64;
localparam ENTROPY_HASH_KEY_MASK_MASK_LO = 0;
localparam ENTROPY_HASH_KEY_MASK_MASK_HI = 63;
localparam ENTROPY_HASH_KEY_MASK_MASK_RESET = 64'h0;
localparam ENTROPY_HASH_KEY_MASK_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam ENTROPY_HASH_KEY_MASK_RO_MASK = 64'h0;
localparam ENTROPY_HASH_KEY_MASK_WO_MASK = 64'h0;
localparam ENTROPY_HASH_KEY_MASK_RESET = 64'h0;

typedef struct packed {
    logic [50:0] reserved0;  // RSVD
    logic  [0:0] ECMP_ROTATION;  // RW
    logic  [1:0] ROTATION_B;  // RW
    logic  [1:0] ROTATION_A;  // RW
    logic  [7:0] reserved1;  // RSVD
} ENTROPY_FWD_HASHING_CFG_t;

localparam ENTROPY_FWD_HASHING_CFG_REG_STRIDE = 48'h8;
localparam ENTROPY_FWD_HASHING_CFG_REG_ENTRIES = 64;
localparam [63:0][47:0] ENTROPY_FWD_HASHING_CFG_CR_ADDR = {48'h2DF8, 48'h2DF0, 48'h2DE8, 48'h2DE0, 48'h2DD8, 48'h2DD0, 48'h2DC8, 48'h2DC0, 48'h2DB8, 48'h2DB0, 48'h2DA8, 48'h2DA0, 48'h2D98, 48'h2D90, 48'h2D88, 48'h2D80, 48'h2D78, 48'h2D70, 48'h2D68, 48'h2D60, 48'h2D58, 48'h2D50, 48'h2D48, 48'h2D40, 48'h2D38, 48'h2D30, 48'h2D28, 48'h2D20, 48'h2D18, 48'h2D10, 48'h2D08, 48'h2D00, 48'h2CF8, 48'h2CF0, 48'h2CE8, 48'h2CE0, 48'h2CD8, 48'h2CD0, 48'h2CC8, 48'h2CC0, 48'h2CB8, 48'h2CB0, 48'h2CA8, 48'h2CA0, 48'h2C98, 48'h2C90, 48'h2C88, 48'h2C80, 48'h2C78, 48'h2C70, 48'h2C68, 48'h2C60, 48'h2C58, 48'h2C50, 48'h2C48, 48'h2C40, 48'h2C38, 48'h2C30, 48'h2C28, 48'h2C20, 48'h2C18, 48'h2C10, 48'h2C08, 48'h2C00};
localparam ENTROPY_FWD_HASHING_CFG_SIZE = 64;
localparam ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION_LO = 12;
localparam ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION_HI = 12;
localparam ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION_RESET = 1'h0;
localparam ENTROPY_FWD_HASHING_CFG_ROTATION_B_LO = 10;
localparam ENTROPY_FWD_HASHING_CFG_ROTATION_B_HI = 11;
localparam ENTROPY_FWD_HASHING_CFG_ROTATION_B_RESET = 2'h1;
localparam ENTROPY_FWD_HASHING_CFG_ROTATION_A_LO = 8;
localparam ENTROPY_FWD_HASHING_CFG_ROTATION_A_HI = 9;
localparam ENTROPY_FWD_HASHING_CFG_ROTATION_A_RESET = 2'h0;
localparam ENTROPY_FWD_HASHING_CFG_USEMASK = 64'h1F00;
localparam ENTROPY_FWD_HASHING_CFG_RO_MASK = 64'h0;
localparam ENTROPY_FWD_HASHING_CFG_WO_MASK = 64'h0;
localparam ENTROPY_FWD_HASHING_CFG_RESET = 64'h400;

typedef struct packed {
    ENTROPY_FWD_HASHING_CFG_t [63:0] ENTROPY_FWD_HASHING_CFG;
} mby_ppe_entropy_map_registers_t;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_ENTROPY_HASH_CFG0_t;

typedef logic [7:0] we_ENTROPY_HASH_CFG1_t;

typedef logic [7:0] we_ENTROPY_META_CFG_t;

typedef logic [7:0] we_ENTROPY_HASH_SYM8_t;

typedef logic [7:0] we_ENTROPY_HASH_SYM16_t;

typedef logic [7:0] we_ENTROPY_HASH_SYM32_t;

typedef logic [7:0] we_ENTROPY_HASH_KEY_MASK_t;

typedef struct packed {
    we_ENTROPY_HASH_CFG0_t ENTROPY_HASH_CFG0;
    we_ENTROPY_HASH_CFG1_t ENTROPY_HASH_CFG1;
    we_ENTROPY_META_CFG_t ENTROPY_META_CFG;
    we_ENTROPY_HASH_SYM8_t ENTROPY_HASH_SYM8;
    we_ENTROPY_HASH_SYM16_t ENTROPY_HASH_SYM16;
    we_ENTROPY_HASH_SYM32_t ENTROPY_HASH_SYM32;
    we_ENTROPY_HASH_KEY_MASK_t ENTROPY_HASH_KEY_MASK;
} mby_ppe_entropy_map_handcoded_t;

typedef logic [7:0] re_ENTROPY_HASH_CFG0_t;

typedef logic [7:0] re_ENTROPY_HASH_CFG1_t;

typedef logic [7:0] re_ENTROPY_META_CFG_t;

typedef logic [7:0] re_ENTROPY_HASH_SYM8_t;

typedef logic [7:0] re_ENTROPY_HASH_SYM16_t;

typedef logic [7:0] re_ENTROPY_HASH_SYM32_t;

typedef logic [7:0] re_ENTROPY_HASH_KEY_MASK_t;

typedef struct packed {
    re_ENTROPY_HASH_CFG0_t ENTROPY_HASH_CFG0;
    re_ENTROPY_HASH_CFG1_t ENTROPY_HASH_CFG1;
    re_ENTROPY_META_CFG_t ENTROPY_META_CFG;
    re_ENTROPY_HASH_SYM8_t ENTROPY_HASH_SYM8;
    re_ENTROPY_HASH_SYM16_t ENTROPY_HASH_SYM16;
    re_ENTROPY_HASH_SYM32_t ENTROPY_HASH_SYM32;
    re_ENTROPY_HASH_KEY_MASK_t ENTROPY_HASH_KEY_MASK;
} mby_ppe_entropy_map_hc_re_t;

typedef logic handcode_rvalid_ENTROPY_HASH_CFG0_t;

typedef logic handcode_rvalid_ENTROPY_HASH_CFG1_t;

typedef logic handcode_rvalid_ENTROPY_META_CFG_t;

typedef logic handcode_rvalid_ENTROPY_HASH_SYM8_t;

typedef logic handcode_rvalid_ENTROPY_HASH_SYM16_t;

typedef logic handcode_rvalid_ENTROPY_HASH_SYM32_t;

typedef logic handcode_rvalid_ENTROPY_HASH_KEY_MASK_t;

typedef struct packed {
    handcode_rvalid_ENTROPY_HASH_CFG0_t ENTROPY_HASH_CFG0;
    handcode_rvalid_ENTROPY_HASH_CFG1_t ENTROPY_HASH_CFG1;
    handcode_rvalid_ENTROPY_META_CFG_t ENTROPY_META_CFG;
    handcode_rvalid_ENTROPY_HASH_SYM8_t ENTROPY_HASH_SYM8;
    handcode_rvalid_ENTROPY_HASH_SYM16_t ENTROPY_HASH_SYM16;
    handcode_rvalid_ENTROPY_HASH_SYM32_t ENTROPY_HASH_SYM32;
    handcode_rvalid_ENTROPY_HASH_KEY_MASK_t ENTROPY_HASH_KEY_MASK;
} mby_ppe_entropy_map_hc_rvalid_t;

typedef logic handcode_wvalid_ENTROPY_HASH_CFG0_t;

typedef logic handcode_wvalid_ENTROPY_HASH_CFG1_t;

typedef logic handcode_wvalid_ENTROPY_META_CFG_t;

typedef logic handcode_wvalid_ENTROPY_HASH_SYM8_t;

typedef logic handcode_wvalid_ENTROPY_HASH_SYM16_t;

typedef logic handcode_wvalid_ENTROPY_HASH_SYM32_t;

typedef logic handcode_wvalid_ENTROPY_HASH_KEY_MASK_t;

typedef struct packed {
    handcode_wvalid_ENTROPY_HASH_CFG0_t ENTROPY_HASH_CFG0;
    handcode_wvalid_ENTROPY_HASH_CFG1_t ENTROPY_HASH_CFG1;
    handcode_wvalid_ENTROPY_META_CFG_t ENTROPY_META_CFG;
    handcode_wvalid_ENTROPY_HASH_SYM8_t ENTROPY_HASH_SYM8;
    handcode_wvalid_ENTROPY_HASH_SYM16_t ENTROPY_HASH_SYM16;
    handcode_wvalid_ENTROPY_HASH_SYM32_t ENTROPY_HASH_SYM32;
    handcode_wvalid_ENTROPY_HASH_KEY_MASK_t ENTROPY_HASH_KEY_MASK;
} mby_ppe_entropy_map_hc_wvalid_t;

typedef logic handcode_error_ENTROPY_HASH_CFG0_t;

typedef logic handcode_error_ENTROPY_HASH_CFG1_t;

typedef logic handcode_error_ENTROPY_META_CFG_t;

typedef logic handcode_error_ENTROPY_HASH_SYM8_t;

typedef logic handcode_error_ENTROPY_HASH_SYM16_t;

typedef logic handcode_error_ENTROPY_HASH_SYM32_t;

typedef logic handcode_error_ENTROPY_HASH_KEY_MASK_t;

typedef struct packed {
    handcode_error_ENTROPY_HASH_CFG0_t ENTROPY_HASH_CFG0;
    handcode_error_ENTROPY_HASH_CFG1_t ENTROPY_HASH_CFG1;
    handcode_error_ENTROPY_META_CFG_t ENTROPY_META_CFG;
    handcode_error_ENTROPY_HASH_SYM8_t ENTROPY_HASH_SYM8;
    handcode_error_ENTROPY_HASH_SYM16_t ENTROPY_HASH_SYM16;
    handcode_error_ENTROPY_HASH_SYM32_t ENTROPY_HASH_SYM32;
    handcode_error_ENTROPY_HASH_KEY_MASK_t ENTROPY_HASH_KEY_MASK;
} mby_ppe_entropy_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    ENTROPY_HASH_CFG0_t ENTROPY_HASH_CFG0;
    ENTROPY_HASH_CFG1_t ENTROPY_HASH_CFG1;
    ENTROPY_META_CFG_t ENTROPY_META_CFG;
    ENTROPY_HASH_SYM8_t ENTROPY_HASH_SYM8;
    ENTROPY_HASH_SYM16_t ENTROPY_HASH_SYM16;
    ENTROPY_HASH_SYM32_t ENTROPY_HASH_SYM32;
    ENTROPY_HASH_KEY_MASK_t ENTROPY_HASH_KEY_MASK;
} mby_ppe_entropy_map_hc_reg_read_t;

typedef struct packed {
    ENTROPY_HASH_CFG0_t ENTROPY_HASH_CFG0;
    ENTROPY_HASH_CFG1_t ENTROPY_HASH_CFG1;
    ENTROPY_META_CFG_t ENTROPY_META_CFG;
    ENTROPY_HASH_SYM8_t ENTROPY_HASH_SYM8;
    ENTROPY_HASH_SYM16_t ENTROPY_HASH_SYM16;
    ENTROPY_HASH_SYM32_t ENTROPY_HASH_SYM32;
    ENTROPY_HASH_KEY_MASK_t ENTROPY_HASH_KEY_MASK;
} mby_ppe_entropy_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_entropy_map_pkg

`endif // MBY_PPE_ENTROPY_MAP_PKG_VH
