///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
// ---------------------------------------------------------------------------------------------------------------------
// -- Author : Luis Alfonso Maeda-Nunez
// -- Project Name : Madison Bay (MBY) 
// -- Description  : Packet Read Controller
//------------------------------------------------------------------------------

module prc 
(
    input logic        clk,
    input logic     arst_n, 

    //EGR Internal Interfaces    
    dp_if.provider  dpb_if, //Dirty Pointer Interface. Connected with the Dirty Pointer Broker
    prc_lcm_if.prc  lcm_if, //Packet Read Controller - Local Congestion Manager Interface
    rrq_if.provider mri_if, //Read Request Interface.  Connected with the Mesh Read Interface

    mtm_prc_if.prc  mtm_if, //Multicast Tag Manager  - Packet Read Controller   Interface
    utm_prc_if.prc  utm_if, //Unicast Tag Manager    - Packet Read Controller   Interface
    pfs_prc_if.prc  pfs_if, //Packet Fetch Scheduler - Packet Read Controller   Interface
    epb_prc_if.prc  epb_if, //Egress Packet Buffer   - Packet Read Controller   Interface
    txc_prc_if.prc  txc_if  //Transmit Controller    - Packet Read Controller   Interface
    
    //EGR External Interfaces

);

endmodule : prc
