magic
tech scmos
timestamp 965071348
<< ndiffusion >>
rect 135 81 139 86
rect 160 85 168 86
rect 127 80 139 81
rect 127 76 139 77
rect 127 68 131 76
rect 160 81 168 82
rect 160 72 168 73
rect 127 67 139 68
rect 127 63 139 64
rect 135 55 139 63
rect 160 68 168 69
rect 160 59 168 60
rect 127 54 139 55
rect 127 46 139 51
rect 160 55 168 56
rect 160 46 168 47
rect 127 42 139 43
rect 160 42 168 43
<< pdiffusion >>
rect 100 91 103 96
rect 100 90 111 91
rect 100 84 111 87
rect 110 76 111 84
rect 184 85 192 86
rect 86 75 111 76
rect 86 67 111 72
rect 184 81 192 82
rect 184 72 192 73
rect 86 63 111 64
rect 94 58 103 63
rect 86 54 94 55
rect 107 52 111 55
rect 184 68 192 69
rect 184 59 192 60
rect 86 46 94 51
rect 86 42 94 43
rect 107 42 111 48
rect 184 55 192 56
rect 184 46 192 47
rect 184 42 192 43
<< ntransistor >>
rect 127 77 139 80
rect 160 82 168 85
rect 160 69 168 72
rect 127 64 139 67
rect 127 51 139 54
rect 160 56 168 59
rect 127 43 139 46
rect 160 43 168 46
<< ptransistor >>
rect 100 87 111 90
rect 86 72 111 75
rect 184 82 192 85
rect 184 69 192 72
rect 86 64 111 67
rect 86 51 94 54
rect 107 48 111 52
rect 184 56 192 59
rect 86 43 94 46
rect 184 43 192 46
<< polysilicon >>
rect 96 87 100 90
rect 111 87 115 90
rect 122 77 127 80
rect 139 77 143 80
rect 122 75 125 77
rect 82 72 86 75
rect 111 72 125 75
rect 156 82 160 85
rect 168 82 184 85
rect 192 82 196 85
rect 156 72 158 82
rect 156 69 160 72
rect 168 69 184 72
rect 192 69 196 72
rect 156 68 158 69
rect 82 64 86 67
rect 111 64 127 67
rect 139 64 143 67
rect 82 51 86 54
rect 94 51 98 54
rect 155 59 158 68
rect 113 52 127 54
rect 103 48 107 52
rect 111 51 127 52
rect 139 51 141 54
rect 155 56 160 59
rect 168 56 184 59
rect 192 56 196 59
rect 111 48 116 51
rect 82 43 86 46
rect 94 43 98 46
rect 155 46 158 56
rect 123 43 127 46
rect 139 43 143 46
rect 155 43 160 46
rect 168 43 184 46
rect 192 43 196 46
<< ndcontact >>
rect 127 81 135 89
rect 160 86 168 94
rect 131 68 139 76
rect 160 73 168 81
rect 127 55 135 63
rect 160 60 168 68
rect 160 47 168 55
rect 127 34 139 42
rect 160 34 168 42
<< pdcontact >>
rect 103 91 111 99
rect 86 76 110 84
rect 184 86 192 94
rect 184 73 192 81
rect 86 55 94 63
rect 103 55 111 63
rect 184 60 192 68
rect 184 47 192 55
rect 86 34 94 42
rect 103 34 111 42
rect 184 34 192 42
<< polycontact >>
rect 148 68 156 85
rect 141 51 149 59
<< metal1 >>
rect 103 98 111 99
rect 103 93 144 98
rect 103 91 119 93
rect 86 76 110 84
rect 114 63 119 91
rect 127 85 135 89
rect 86 58 119 63
rect 123 81 135 85
rect 139 85 144 93
rect 160 86 168 94
rect 184 86 192 94
rect 123 63 127 81
rect 139 76 156 85
rect 131 68 156 76
rect 160 73 192 81
rect 123 59 135 63
rect 160 60 168 68
rect 86 55 94 58
rect 103 55 111 58
rect 127 55 135 59
rect 141 55 149 59
rect 172 55 180 73
rect 184 60 192 68
rect 141 51 192 55
rect 160 47 192 51
rect 86 34 111 42
rect 127 34 168 42
rect 184 34 192 42
<< labels >>
rlabel metal1 107 38 107 38 1 Vdd!
rlabel polysilicon 85 73 85 73 3 b
rlabel polysilicon 85 65 85 65 3 a
rlabel polysilicon 85 52 85 52 3 b
rlabel polysilicon 85 44 85 44 3 a
rlabel metal1 90 80 90 80 1 Vdd!
rlabel metal1 90 38 90 38 1 Vdd!
rlabel metal1 133 38 133 38 1 GND!
rlabel polysilicon 126 52 126 52 1 x
rlabel polysilicon 126 78 126 78 1 b
rlabel polysilicon 126 65 126 65 1 a
rlabel metal1 135 73 135 73 1 _x
rlabel polysilicon 193 83 193 83 1 _x
rlabel pdcontact 188 90 188 90 5 Vdd!
rlabel ndcontact 164 90 164 90 5 GND!
rlabel ndcontact 164 38 164 38 1 GND!
rlabel polysilicon 193 58 193 58 5 _x
rlabel polysilicon 193 45 193 45 5 _x
rlabel pdcontact 188 38 188 38 1 Vdd!
rlabel pdcontact 188 51 188 51 5 x
rlabel ndcontact 164 64 164 64 1 GND!
rlabel polysilicon 193 70 193 70 1 _x
rlabel pdcontact 188 64 188 64 1 Vdd!
rlabel pdcontact 188 77 188 77 1 x
rlabel ndcontact 164 77 164 77 1 x
rlabel ndcontact 164 51 164 51 5 x
rlabel polysilicon 126 44 126 44 1 _SReset!
rlabel polysilicon 112 49 112 49 5 x
rlabel metal1 90 59 90 59 1 _x
rlabel metal1 107 59 107 59 1 _x
rlabel metal1 107 95 107 95 5 _x
rlabel polysilicon 99 88 99 88 1 _PReset!
rlabel space 192 34 197 94 3 ^p2
rlabel space 168 33 198 95 3 ^n2
rlabel space 81 34 86 84 7 ^p1
<< end >>
