magic
tech scmos
timestamp 988943070
<< nselect >>
rect -34 44 0 83
rect -28 37 0 44
rect -34 11 0 37
rect -28 10 0 11
rect -34 -24 0 10
<< pselect >>
rect 0 44 34 80
rect 0 43 28 44
rect 0 11 34 43
rect 0 10 28 11
rect 0 -22 34 10
<< ndiffusion >>
rect -28 71 -8 72
rect -28 67 -8 68
rect -28 58 -8 59
rect -28 52 -8 55
rect -28 28 -8 29
rect -28 20 -8 25
rect -28 14 -8 17
rect -28 3 -8 6
rect -28 -1 -8 0
rect -28 -10 -8 -9
rect -28 -14 -8 -13
<< pdiffusion >>
rect 8 66 28 67
rect 8 58 28 63
rect 8 52 28 55
rect 8 33 28 36
rect 8 29 28 30
rect 8 20 28 21
rect 8 14 28 17
rect 8 3 28 6
rect 8 -5 28 0
rect 8 -9 28 -8
<< ntransistor >>
rect -28 68 -8 71
rect -28 55 -8 58
rect -28 25 -8 28
rect -28 17 -8 20
rect -28 0 -8 3
rect -28 -13 -8 -10
<< ptransistor >>
rect 8 63 28 66
rect 8 55 28 58
rect 8 30 28 33
rect 8 17 28 20
rect 8 0 28 3
rect 8 -8 28 -5
<< polysilicon >>
rect -32 68 -28 71
rect -8 68 0 71
rect -3 66 0 68
rect -3 63 8 66
rect 28 63 32 66
rect -32 55 -28 58
rect -8 55 8 58
rect 28 55 32 58
rect 1 33 4 40
rect 1 30 8 33
rect 28 30 32 33
rect 1 28 4 30
rect -32 25 -28 28
rect -8 25 4 28
rect -32 17 -28 20
rect -8 17 -4 20
rect 4 17 8 20
rect 28 17 32 20
rect -32 0 -28 3
rect -8 0 8 3
rect 28 0 32 3
rect -6 -8 8 -5
rect 28 -8 32 -5
rect -6 -10 -3 -8
rect -32 -13 -28 -10
rect -8 -13 -3 -10
<< ndcontact >>
rect -28 72 -8 80
rect -28 59 -8 67
rect -28 44 -8 52
rect -28 29 -8 37
rect -28 6 -8 14
rect -28 -9 -8 -1
rect -28 -22 -8 -14
<< pdcontact >>
rect 8 67 28 75
rect 8 36 28 52
rect 8 21 28 29
rect 8 6 28 14
rect 8 -17 28 -9
<< polycontact >>
rect -4 40 4 48
rect -4 12 4 20
<< metal1 >>
rect -28 72 -8 80
rect 8 67 28 75
rect -28 63 12 67
rect -28 59 -8 63
rect -28 44 -8 52
rect -2 48 2 63
rect -4 40 4 48
rect -28 30 -8 37
rect 8 36 28 52
rect -28 24 28 30
rect 8 21 28 24
rect -28 6 -8 14
rect -4 12 4 20
rect -28 -5 -8 -1
rect -2 -5 2 12
rect 8 6 28 14
rect -28 -9 12 -5
rect -28 -22 -8 -14
rect 8 -17 28 -9
<< labels >>
rlabel metal1 -28 24 28 30 1 av
rlabel space -35 -24 -28 10 7 ^n01
rlabel space -35 11 -28 37 7 ^n03
rlabel space -35 44 -28 83 7 ^n23
rlabel space 28 -22 35 10 3 ^p01
rlabel space 28 11 35 43 3 ^p03
rlabel space 28 44 35 80 3 ^p23
rlabel polysilicon -32 -13 -28 -10 1 a0|pin|w|2|poly
rlabel polysilicon -7 -13 -3 -10 1 a0|pin|w|2|poly
rlabel polysilicon 28 -8 32 -5 1 a0|pin|w|2|poly
rlabel polysilicon 28 0 32 3 1 a1|pin|w|3|poly
rlabel polysilicon -32 0 -28 3 1 a1|pin|w|3|poly
rlabel polysilicon 28 55 32 58 1 a2|pin|w|4|poly
rlabel polysilicon -32 55 -28 58 1 a2|pin|w|4|poly
rlabel polysilicon -32 68 -28 71 1 a3|pin|w|5|poly
rlabel polysilicon -4 68 0 71 1 a3|pin|w|5|poly
rlabel polysilicon 28 63 32 66 1 a3|pin|w|5|poly
rlabel metal1 -28 -9 -8 -1 1 _a_01|pin|s|6
rlabel metal1 -28 59 -8 67 1 _a_23|pin|s|7
rlabel metal1 8 67 28 75 1 _a_23|pin|s|7
rlabel metal1 8 -17 28 -9 1 _a_01|pin|s|6
rlabel metal1 8 36 28 52 1 Vdd!|pin|s|1
rlabel metal1 8 6 28 14 1 Vdd!|pin|s|0
rlabel metal1 -28 6 -8 14 1 GND!|pin|s|1
rlabel metal1 -28 44 -8 52 1 GND!|pin|s|2
rlabel metal1 -28 72 -8 80 1 GND!|pin|s|3
rlabel metal1 -28 -22 -8 -14 1 GND!|pin|s|0
rlabel metal1 -28 24 -8 37 1 av
rlabel metal1 8 21 28 29 1 av
<< end >>
