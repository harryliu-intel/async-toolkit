module read_ecc
  (
input  logic [34-1:0] i_data,
input  logic [7-1:0] i_chk,

output logic          o_err_detect,
output logic          o_err_multpl,
output logic [34-1:0] o_data
  );
logic  xor0000;
logic  xor0001;
logic  xor0002;
logic  xor0003;
logic  xor0004;
logic  xor0005;
logic  xor0006;
logic  xor0007;
logic  xor0008;
logic  xor0009;
logic  xor0010;
logic  xor0011;
logic  xor0012;
logic  xor0013;
logic  xor0014;
logic  xor0015;
logic  xor0016;
logic  xor0017;
logic  xor0018;
logic  xor0019;
logic  xor0020;
logic  xor0021;
logic  xor0022;
logic  xor0023;
logic  xor0024;
logic  xor0025;
logic  xor0026;
logic  xor0027;
logic  xor0028;
logic  xor0029;
logic  xor0030;
logic  xor0031;
logic  xor0032;
logic  xor0033;
logic  xor0034;
logic  xor0035;
logic  xor0036;
logic  xor0037;
logic  xor0038;
logic  xor0039;
logic  xor0040;
logic  xor0041;
logic  xor0042;
logic  xor0043;
logic[5:-1] ecc_parity;
logic[40:0] input_data;
logic[40:0] corrected;
logic  syn_0000_n;
logic  syn_0000;
logic  syn_0001_n;
logic  syn_0001;
logic  syn_0002_n;
logic  syn_0002;
logic  syn_0003_n;
logic  syn_0003;
logic  syn_0004_n;
logic  syn_0004;
logic  syn_0005_n;
logic  syn_0005;
logic  nand0056;
logic  nand0057;
logic  nand0058;
logic  nand0059;
logic  nand0060;
logic  nand0061;
logic  nand0062;
logic  nand0063;
logic  nand0064;
logic  nand0065;
logic  nand0066;
logic  nand0067;
logic  nand0068;
logic  nand0069;
logic  nand0070;
logic  nand0071;
logic  nor0072;
logic  nor0073;
logic  nor0074;
logic  nor0075;
logic  nor0076;
logic  nor0077;
logic  nor0078;
logic  nor0079;
logic  nor0080;
logic  nor0081;
logic  nor0082;
logic  nor0083;
logic  nor0084;
logic  nor0085;
logic  nor0086;
logic  nor0087;
logic  nor0088;
logic  nor0089;
logic  nor0090;
logic  nor0091;
logic  nor0092;
logic  nor0093;
logic  nor0094;
logic  nor0095;
logic  nor0096;
logic  nor0097;
logic  nor0098;
logic  nor0099;
logic  nor0100;
logic  nor0101;
logic  nor0102;
logic  nor0103;
logic  nor0104;
logic  nor0105;
logic  nor0106;
logic  nor0107;
logic  nor0108;
logic  nor0109;
logic  nor0110;
logic  nor0111;
logic  nor0112;
assign xor0000 = (input_data[0001]^input_data[0000]^input_data[0003]^input_data[0002]); 
assign xor0001 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); 
assign xor0002 = (input_data[0009]^input_data[0008]^input_data[0011]^input_data[0010]); 
assign xor0003 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); 
assign xor0004 = (input_data[0019]^input_data[0018]^input_data[0017]^input_data[0016]); 
assign xor0005 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); 
assign xor0006 = (input_data[0025]^input_data[0024]^input_data[0027]^input_data[0026]); 
assign xor0007 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); 
assign xor0008 = (input_data[0035]^input_data[0034]^input_data[0033]^input_data[0032]); 
assign xor0009 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); 
assign xor0010 = input_data[0040];
assign xor0011 = (input_data[0005]^input_data[0007]^input_data[0001]^input_data[0003]); 
assign xor0012 = (input_data[0009]^input_data[0015]^input_data[0011]^input_data[0013]); 
assign xor0013 = (input_data[0019]^input_data[0017]^input_data[0021]^input_data[0023]); 
assign xor0014 = (input_data[0025]^input_data[0027]^input_data[0031]^input_data[0029]); 
assign xor0015 = (input_data[0035]^input_data[0037]^input_data[0033]^input_data[0039]); 
assign xor0016 = (input_data[0007]^input_data[0006]^input_data[0003]^input_data[0002]); 
assign xor0017 = (input_data[0015]^input_data[0014]^input_data[0011]^input_data[0010]); 
assign xor0018 = (input_data[0019]^input_data[0018]^input_data[0023]^input_data[0022]); 
assign xor0019 = (input_data[0027]^input_data[0031]^input_data[0030]^input_data[0026]); 
assign xor0020 = (input_data[0035]^input_data[0034]^input_data[0039]^input_data[0038]); 
assign xor0021 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); 
assign xor0022 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); 
assign xor0023 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); 
assign xor0024 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); 
assign xor0025 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); 
assign xor0026 = (xor0013^xor0014^xor0011^xor0012); 
assign xor0027 = xor0015;
assign xor0028 = (xor0027^xor0026); 
assign xor0029 = (xor0017^xor0018^xor0016^xor0019); 
assign xor0030 = xor0020;
assign xor0031 = (xor0030^xor0029); 
assign xor0032 = (xor0023^xor0024^xor0021^xor0022); 
assign xor0033 = xor0025;
assign xor0034 = (xor0033^xor0032); 
assign xor0035 = (xor0002^xor0010^xor0006^xor0022); 
assign xor0036 = xor0024;
assign xor0037 = (xor0035^xor0036); 
assign xor0038 = (xor0036^xor0023^xor0006^xor0004); 
assign xor0039 = (xor0010^xor0008^xor0033); 
assign xor0040 = (xor0002^xor0000^xor0021^xor0022); 
assign xor0041 = xor0038;
assign xor0042 = (xor0040^xor0041); 
assign xor0043 = (xor0039^xor0042); 
assign ecc_parity[-1] = xor0043;
assign ecc_parity[0] = xor0028;
assign ecc_parity[1] = xor0031;
assign ecc_parity[2] = xor0034;
assign ecc_parity[3] = xor0037;
assign ecc_parity[4] = xor0038;
assign ecc_parity[5] = xor0039;
assign input_data[0] = i_chk    [0];
assign input_data[1] = i_chk    [1];
assign input_data[2] = i_chk    [2];
assign input_data[3] = i_data   [0];
assign o_data    [0] = corrected[3];
assign input_data[4] = i_chk    [3];
assign input_data[5] = i_data   [1];
assign o_data    [1] = corrected[5];
assign input_data[6] = i_data   [2];
assign o_data    [2] = corrected[6];
assign input_data[7] = i_data   [3];
assign o_data    [3] = corrected[7];
assign input_data[8] = i_chk    [4];
assign input_data[9] = i_data   [4];
assign o_data    [4] = corrected[9];
assign input_data[10] = i_data   [5];
assign o_data    [5] = corrected[10];
assign input_data[11] = i_data   [6];
assign o_data    [6] = corrected[11];
assign input_data[12] = i_data   [7];
assign o_data    [7] = corrected[12];
assign input_data[13] = i_data   [8];
assign o_data    [8] = corrected[13];
assign input_data[14] = i_data   [9];
assign o_data    [9] = corrected[14];
assign input_data[15] = i_data   [10];
assign o_data    [10] = corrected[15];
assign input_data[16] = i_chk    [5];
assign input_data[17] = i_data   [11];
assign o_data    [11] = corrected[17];
assign input_data[18] = i_data   [12];
assign o_data    [12] = corrected[18];
assign input_data[19] = i_data   [13];
assign o_data    [13] = corrected[19];
assign input_data[20] = i_data   [14];
assign o_data    [14] = corrected[20];
assign input_data[21] = i_data   [15];
assign o_data    [15] = corrected[21];
assign input_data[22] = i_data   [16];
assign o_data    [16] = corrected[22];
assign input_data[23] = i_data   [17];
assign o_data    [17] = corrected[23];
assign input_data[24] = i_data   [18];
assign o_data    [18] = corrected[24];
assign input_data[25] = i_data   [19];
assign o_data    [19] = corrected[25];
assign input_data[26] = i_data   [20];
assign o_data    [20] = corrected[26];
assign input_data[27] = i_data   [21];
assign o_data    [21] = corrected[27];
assign input_data[28] = i_data   [22];
assign o_data    [22] = corrected[28];
assign input_data[29] = i_data   [23];
assign o_data    [23] = corrected[29];
assign input_data[30] = i_data   [24];
assign o_data    [24] = corrected[30];
assign input_data[31] = i_data   [25];
assign o_data    [25] = corrected[31];
assign input_data[32] = i_chk    [6];
assign input_data[33] = i_data   [26];
assign o_data    [26] = corrected[33];
assign input_data[34] = i_data   [27];
assign o_data    [27] = corrected[34];
assign input_data[35] = i_data   [28];
assign o_data    [28] = corrected[35];
assign input_data[36] = i_data   [29];
assign o_data    [29] = corrected[36];
assign input_data[37] = i_data   [30];
assign o_data    [30] = corrected[37];
assign input_data[38] = i_data   [31];
assign o_data    [31] = corrected[38];
assign input_data[39] = i_data   [32];
assign o_data    [32] = corrected[39];
assign input_data[40] = i_data   [33];
assign o_data    [33] = corrected[40];
assign syn_0000_n = !(ecc_parity[0]); 
assign syn_0000 = !(syn_0000_n); 
assign syn_0001_n = !(ecc_parity[1]); 
assign syn_0001 = !(syn_0001_n); 
assign syn_0002_n = !(ecc_parity[2]); 
assign syn_0002 = !(syn_0002_n); 
assign syn_0003_n = !(ecc_parity[3]); 
assign syn_0003 = !(syn_0003_n); 
assign syn_0004_n = !(ecc_parity[4]); 
assign syn_0004 = !(syn_0004_n); 
assign syn_0005_n = !(ecc_parity[5]); 
assign syn_0005 = !(syn_0005_n); 
assign nand0056 = !(syn_0002_n&syn_0001_n&syn_0000_n); 
assign nand0057 = !(syn_0002_n&syn_0001_n&syn_0000); 
assign nand0058 = !(syn_0002_n&syn_0001&syn_0000_n); 
assign nand0059 = !(syn_0002_n&syn_0001&syn_0000); 
assign nand0060 = !(syn_0002&syn_0001_n&syn_0000_n); 
assign nand0061 = !(syn_0002&syn_0001_n&syn_0000); 
assign nand0062 = !(syn_0002&syn_0001&syn_0000_n); 
assign nand0063 = !(syn_0002&syn_0001&syn_0000); 
assign nand0064 = !(syn_0003_n&syn_0005_n&syn_0004_n); 
assign nand0065 = !(syn_0003&syn_0005_n&syn_0004_n); 
assign nand0066 = !(syn_0003_n&syn_0004&syn_0005_n); 
assign nand0067 = !(syn_0004&syn_0003&syn_0005_n); 
assign nand0068 = !(syn_0003_n&syn_0005&syn_0004_n); 
assign nand0069 = !(syn_0003&syn_0005&syn_0004_n); 
assign nand0070 = !(syn_0003_n&syn_0004&syn_0005); 
assign nand0071 = !(syn_0004&syn_0003&syn_0005); 
assign nor0072 = !(nand0056|nand0064); 
assign invert0000 = nor0072;
assign nor0073 = !(nand0057|nand0064); 
assign invert0001 = nor0073;
assign nor0074 = !(nand0064|nand0058); 
assign invert0002 = nor0074;
assign nor0075 = !(nand0059|nand0064); 
assign invert0003 = nor0075;
assign nor0076 = !(nand0060|nand0064); 
assign invert0004 = nor0076;
assign nor0077 = !(nand0064|nand0061); 
assign invert0005 = nor0077;
assign nor0078 = !(nand0062|nand0064); 
assign invert0006 = nor0078;
assign nor0079 = !(nand0064|nand0063); 
assign invert0007 = nor0079;
assign nor0080 = !(nand0065|nand0056); 
assign invert0008 = nor0080;
assign nor0081 = !(nand0057|nand0065); 
assign invert0009 = nor0081;
assign nor0082 = !(nand0065|nand0058); 
assign invert0010 = nor0082;
assign nor0083 = !(nand0065|nand0059); 
assign invert0011 = nor0083;
assign nor0084 = !(nand0060|nand0065); 
assign invert0012 = nor0084;
assign nor0085 = !(nand0065|nand0061); 
assign invert0013 = nor0085;
assign nor0086 = !(nand0065|nand0062); 
assign invert0014 = nor0086;
assign nor0087 = !(nand0065|nand0063); 
assign invert0015 = nor0087;
assign nor0088 = !(nand0056|nand0066); 
assign invert0016 = nor0088;
assign nor0089 = !(nand0057|nand0066); 
assign invert0017 = nor0089;
assign nor0090 = !(nand0066|nand0058); 
assign invert0018 = nor0090;
assign nor0091 = !(nand0059|nand0066); 
assign invert0019 = nor0091;
assign nor0092 = !(nand0060|nand0066); 
assign invert0020 = nor0092;
assign nor0093 = !(nand0061|nand0066); 
assign invert0021 = nor0093;
assign nor0094 = !(nand0062|nand0066); 
assign invert0022 = nor0094;
assign nor0095 = !(nand0066|nand0063); 
assign invert0023 = nor0095;
assign nor0096 = !(nand0067|nand0056); 
assign invert0024 = nor0096;
assign nor0097 = !(nand0057|nand0067); 
assign invert0025 = nor0097;
assign nor0098 = !(nand0067|nand0058); 
assign invert0026 = nor0098;
assign nor0099 = !(nand0067|nand0059); 
assign invert0027 = nor0099;
assign nor0100 = !(nand0060|nand0067); 
assign invert0028 = nor0100;
assign nor0101 = !(nand0067|nand0061); 
assign invert0029 = nor0101;
assign nor0102 = !(nand0062|nand0067); 
assign invert0030 = nor0102;
assign nor0103 = !(nand0067|nand0063); 
assign invert0031 = nor0103;
assign nor0104 = !(nand0068|nand0056); 
assign invert0032 = nor0104;
assign nor0105 = !(nand0068|nand0057); 
assign invert0033 = nor0105;
assign nor0106 = !(nand0068|nand0058); 
assign invert0034 = nor0106;
assign nor0107 = !(nand0068|nand0059); 
assign invert0035 = nor0107;
assign nor0108 = !(nand0060|nand0068); 
assign invert0036 = nor0108;
assign nor0109 = !(nand0068|nand0061); 
assign invert0037 = nor0109;
assign nor0110 = !(nand0068|nand0062); 
assign invert0038 = nor0110;
assign nor0111 = !(nand0068|nand0063); 
assign invert0039 = nor0111;
assign nor0112 = !(nand0056|nand0069); 
assign invert0040 = nor0112;
assign corrected[0] = (invert0000^input_data[0]); 
assign corrected[1] = (invert0001^input_data[1]); 
assign corrected[2] = (input_data[2]^invert0002); 
assign corrected[3] = (input_data[3]^invert0003); 
assign corrected[4] = (invert0004^input_data[4]); 
assign corrected[5] = (input_data[5]^invert0005); 
assign corrected[6] = (input_data[6]^invert0006); 
assign corrected[7] = (invert0007^input_data[7]); 
assign corrected[8] = (input_data[8]^invert0008); 
assign corrected[9] = (input_data[9]^invert0009); 
assign corrected[10] = (input_data[10]^invert0010); 
assign corrected[11] = (invert0011^input_data[11]); 
assign corrected[12] = (input_data[12]^invert0012); 
assign corrected[13] = (input_data[13]^invert0013); 
assign corrected[14] = (input_data[14]^invert0014); 
assign corrected[15] = (input_data[15]^invert0015); 
assign corrected[16] = (input_data[16]^invert0016); 
assign corrected[17] = (invert0017^input_data[17]); 
assign corrected[18] = (invert0018^input_data[18]); 
assign corrected[19] = (invert0019^input_data[19]); 
assign corrected[20] = (input_data[20]^invert0020); 
assign corrected[21] = (input_data[21]^invert0021); 
assign corrected[22] = (invert0022^input_data[22]); 
assign corrected[23] = (input_data[23]^invert0023); 
assign corrected[24] = (invert0024^input_data[24]); 
assign corrected[25] = (input_data[25]^invert0025); 
assign corrected[26] = (input_data[26]^invert0026); 
assign corrected[27] = (input_data[27]^invert0027); 
assign corrected[28] = (input_data[28]^invert0028); 
assign corrected[29] = (invert0029^input_data[29]); 
assign corrected[30] = (input_data[30]^invert0030); 
assign corrected[31] = (input_data[31]^invert0031); 
assign corrected[32] = (input_data[32]^invert0032); 
assign corrected[33] = (input_data[33]^invert0033); 
assign corrected[34] = (invert0034^input_data[34]); 
assign corrected[35] = (input_data[35]^invert0035); 
assign corrected[36] = (input_data[36]^invert0036); 
assign corrected[37] = (invert0037^input_data[37]); 
assign corrected[38] = (input_data[38]^invert0038); 
assign corrected[39] = (invert0039^input_data[39]); 
assign corrected[40] = (input_data[40]^invert0040); 
assign o_err_detect = |(ecc_parity[6-1:-1]);
assign o_err_multpl = o_err_detect & !ecc_parity[-1];
endmodule
