///
///  INTEL CONFIDENTIAL
///
///  Copyright 2017 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
// ---------------------------------------------------------------------------------------------------------------------
// -- Author : Jim McCormick <jim.mccormick@intel.com>
// -- Project Name : ??? 
// -- Description  : The DUT interface 
// ---------------------------------------------------------------------------------------------------------------------

// This is a connectivity only interface and thus is just a named bundle of nets that can be passed around as a group 
// to save typing.  Anywhere an interface is defined, individual nets in the interface can be referenced as follows:    
//
//      <interface name>.<net name>
//

interface tmpl_dut_if (
   input clk                                        // clk is passed in a parameter and becomes part of the interface
);


// local paramters
localparam NUM_INPUTS  = tmpl_pkg::NUM_INPUTS;
localparam NUM_OUTPUTS = tmpl_pkg::NUM_OUTPUTS;


// DUT inputs  (direction not specified in this interface)
logic               i_reset;                                // reset
tmpl_pkg::req_in_t  i_reqs          [NUM_INPUTS-1:0];       // incoming request ports


// DUT outputs  (direction not specified in this interface)
tmpl_pkg::req_out_t o_reqs          [NUM_OUTPUTS-1:0];      // outgoing request ports


endinterface // tmpl_dut_if
