///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_trig_apply_map_pkg.vh                              
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_TRIG_APPLY_MAP_PKG_VH
`define MBY_PPE_TRIG_APPLY_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_trig_apply_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_trig_apply_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_trig_apply_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_trig_apply_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic  [1:0] MATCH_TX;  // RW
    logic  [4:0] MATCH_RANDOM_THRESHOLD;  // RW
    logic  [0:0] MATCH_RANDOM_IF_LESS;  // RW
    logic  [0:0] MATCH_RANDOM_NUMBER;  // RW
    logic  [0:0] MATCH_BY_PRECEDENCE;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [1:0] MATCH_EGRESS_DOMAIN;  // RW
    logic  [1:0] MATCH_DEST_GLORT;  // RW
    logic  [1:0] reserved2;  // RSVD
    logic  [1:0] MATCH_TC;  // RW
    logic  [1:0] MATCH_CGRP;  // RW
    logic  [1:0] MATCH_VLAN;  // RW
    logic  [3:0] reserved3;  // RSVD
    logic  [1:0] LEARN;  // RW
    logic  [3:0] reserved4;  // RSVD
} TRIGGER_CONDITION_CFG_t;

localparam TRIGGER_CONDITION_CFG_REG_STRIDE = 48'h8;
localparam TRIGGER_CONDITION_CFG_REG_ENTRIES = 96;
localparam TRIGGER_CONDITION_CFG_CR_ADDR = 48'h0;
localparam TRIGGER_CONDITION_CFG_SIZE = 64;
localparam TRIGGER_CONDITION_CFG_MATCH_TX_LO = 34;
localparam TRIGGER_CONDITION_CFG_MATCH_TX_HI = 35;
localparam TRIGGER_CONDITION_CFG_MATCH_TX_RESET = 2'h0;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_THRESHOLD_LO = 29;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_THRESHOLD_HI = 33;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_THRESHOLD_RESET = 5'h18;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_IF_LESS_LO = 28;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_IF_LESS_HI = 28;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_IF_LESS_RESET = 1'h1;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_NUMBER_LO = 27;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_NUMBER_HI = 27;
localparam TRIGGER_CONDITION_CFG_MATCH_RANDOM_NUMBER_RESET = 1'h0;
localparam TRIGGER_CONDITION_CFG_MATCH_BY_PRECEDENCE_LO = 26;
localparam TRIGGER_CONDITION_CFG_MATCH_BY_PRECEDENCE_HI = 26;
localparam TRIGGER_CONDITION_CFG_MATCH_BY_PRECEDENCE_RESET = 1'h0;
localparam TRIGGER_CONDITION_CFG_MATCH_EGRESS_DOMAIN_LO = 20;
localparam TRIGGER_CONDITION_CFG_MATCH_EGRESS_DOMAIN_HI = 21;
localparam TRIGGER_CONDITION_CFG_MATCH_EGRESS_DOMAIN_RESET = 2'h2;
localparam TRIGGER_CONDITION_CFG_MATCH_DEST_GLORT_LO = 18;
localparam TRIGGER_CONDITION_CFG_MATCH_DEST_GLORT_HI = 19;
localparam TRIGGER_CONDITION_CFG_MATCH_DEST_GLORT_RESET = 2'h2;
localparam TRIGGER_CONDITION_CFG_MATCH_TC_LO = 14;
localparam TRIGGER_CONDITION_CFG_MATCH_TC_HI = 15;
localparam TRIGGER_CONDITION_CFG_MATCH_TC_RESET = 2'h2;
localparam TRIGGER_CONDITION_CFG_MATCH_CGRP_LO = 12;
localparam TRIGGER_CONDITION_CFG_MATCH_CGRP_HI = 13;
localparam TRIGGER_CONDITION_CFG_MATCH_CGRP_RESET = 2'h2;
localparam TRIGGER_CONDITION_CFG_MATCH_VLAN_LO = 10;
localparam TRIGGER_CONDITION_CFG_MATCH_VLAN_HI = 11;
localparam TRIGGER_CONDITION_CFG_MATCH_VLAN_RESET = 2'h2;
localparam TRIGGER_CONDITION_CFG_LEARN_LO = 4;
localparam TRIGGER_CONDITION_CFG_LEARN_HI = 5;
localparam TRIGGER_CONDITION_CFG_LEARN_RESET = 2'h2;
localparam TRIGGER_CONDITION_CFG_USEMASK = 64'hFFC3CFC30;
localparam TRIGGER_CONDITION_CFG_RO_MASK = 64'h0;
localparam TRIGGER_CONDITION_CFG_WO_MASK = 64'h0;
localparam TRIGGER_CONDITION_CFG_RESET = 64'h31028A820;

typedef struct packed {
    logic  [4:0] reserved0;  // RSVD
    logic [13:0] EGRESS_DOMAIN_MASK;  // RW
    logic  [0:0] reserved1;  // RSVD
    logic [13:0] EGRESS_DOMAIN_VALUE;  // RW
    logic  [3:0] reserved2;  // RSVD
    logic  [1:0] ROUTED_MASK;  // RW
    logic  [2:0] FRAME_CLASS_MASK;  // RW
    logic  [2:0] TC;  // RW
    logic  [5:0] VID_ID;  // RW
    logic [11:0] reserved3;  // RSVD
} TRIGGER_CONDITION_PARAM_t;

localparam TRIGGER_CONDITION_PARAM_REG_STRIDE = 48'h8;
localparam TRIGGER_CONDITION_PARAM_REG_ENTRIES = 96;
localparam TRIGGER_CONDITION_PARAM_CR_ADDR = 48'h300;
localparam TRIGGER_CONDITION_PARAM_SIZE = 64;
localparam TRIGGER_CONDITION_PARAM_EGRESS_DOMAIN_MASK_LO = 45;
localparam TRIGGER_CONDITION_PARAM_EGRESS_DOMAIN_MASK_HI = 58;
localparam TRIGGER_CONDITION_PARAM_EGRESS_DOMAIN_MASK_RESET = 14'h0;
localparam TRIGGER_CONDITION_PARAM_EGRESS_DOMAIN_VALUE_LO = 30;
localparam TRIGGER_CONDITION_PARAM_EGRESS_DOMAIN_VALUE_HI = 43;
localparam TRIGGER_CONDITION_PARAM_EGRESS_DOMAIN_VALUE_RESET = 14'h0;
localparam TRIGGER_CONDITION_PARAM_ROUTED_MASK_LO = 24;
localparam TRIGGER_CONDITION_PARAM_ROUTED_MASK_HI = 25;
localparam TRIGGER_CONDITION_PARAM_ROUTED_MASK_RESET = 2'h3;
localparam TRIGGER_CONDITION_PARAM_FRAME_CLASS_MASK_LO = 21;
localparam TRIGGER_CONDITION_PARAM_FRAME_CLASS_MASK_HI = 23;
localparam TRIGGER_CONDITION_PARAM_FRAME_CLASS_MASK_RESET = 3'h7;
localparam TRIGGER_CONDITION_PARAM_TC_LO = 18;
localparam TRIGGER_CONDITION_PARAM_TC_HI = 20;
localparam TRIGGER_CONDITION_PARAM_TC_RESET = 3'h0;
localparam TRIGGER_CONDITION_PARAM_VID_ID_LO = 12;
localparam TRIGGER_CONDITION_PARAM_VID_ID_HI = 17;
localparam TRIGGER_CONDITION_PARAM_VID_ID_RESET = 6'h0;
localparam TRIGGER_CONDITION_PARAM_USEMASK = 64'h7FFEFFFC3FFF000;
localparam TRIGGER_CONDITION_PARAM_RO_MASK = 64'h0;
localparam TRIGGER_CONDITION_PARAM_WO_MASK = 64'h0;
localparam TRIGGER_CONDITION_PARAM_RESET = 64'h3E00000;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic  [7:0] CGRP_MASK;  // RW
    logic  [7:0] CGRP_ID;  // RW
} TRIGGER_CONDITION_CGRP_t;

localparam TRIGGER_CONDITION_CGRP_REG_STRIDE = 48'h8;
localparam TRIGGER_CONDITION_CGRP_REG_ENTRIES = 96;
localparam TRIGGER_CONDITION_CGRP_CR_ADDR = 48'h600;
localparam TRIGGER_CONDITION_CGRP_SIZE = 64;
localparam TRIGGER_CONDITION_CGRP_CGRP_MASK_LO = 8;
localparam TRIGGER_CONDITION_CGRP_CGRP_MASK_HI = 15;
localparam TRIGGER_CONDITION_CGRP_CGRP_MASK_RESET = 8'h0;
localparam TRIGGER_CONDITION_CGRP_CGRP_ID_LO = 0;
localparam TRIGGER_CONDITION_CGRP_CGRP_ID_HI = 7;
localparam TRIGGER_CONDITION_CGRP_CGRP_ID_RESET = 8'h0;
localparam TRIGGER_CONDITION_CGRP_USEMASK = 64'hFFFF;
localparam TRIGGER_CONDITION_CGRP_RO_MASK = 64'h0;
localparam TRIGGER_CONDITION_CGRP_WO_MASK = 64'h0;
localparam TRIGGER_CONDITION_CGRP_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [15:0] GLORT_MASK;  // RW
    logic [15:0] DEST_GLORT;  // RW
} TRIGGER_CONDITION_GLORT_t;

localparam TRIGGER_CONDITION_GLORT_REG_STRIDE = 48'h8;
localparam TRIGGER_CONDITION_GLORT_REG_ENTRIES = 96;
localparam TRIGGER_CONDITION_GLORT_CR_ADDR = 48'h900;
localparam TRIGGER_CONDITION_GLORT_SIZE = 64;
localparam TRIGGER_CONDITION_GLORT_GLORT_MASK_LO = 16;
localparam TRIGGER_CONDITION_GLORT_GLORT_MASK_HI = 31;
localparam TRIGGER_CONDITION_GLORT_GLORT_MASK_RESET = 16'h0;
localparam TRIGGER_CONDITION_GLORT_DEST_GLORT_LO = 0;
localparam TRIGGER_CONDITION_GLORT_DEST_GLORT_HI = 15;
localparam TRIGGER_CONDITION_GLORT_DEST_GLORT_RESET = 16'h0;
localparam TRIGGER_CONDITION_GLORT_USEMASK = 64'hFFFFFFFF;
localparam TRIGGER_CONDITION_GLORT_RO_MASK = 64'h0;
localparam TRIGGER_CONDITION_GLORT_WO_MASK = 64'h0;
localparam TRIGGER_CONDITION_GLORT_RESET = 64'h0;

typedef struct packed {
    logic [45:0] reserved0;  // RSVD
    logic [17:0] SRC_PORT_MASK;  // RW
} TRIGGER_CONDITION_RX_t;

localparam TRIGGER_CONDITION_RX_REG_STRIDE = 48'h8;
localparam TRIGGER_CONDITION_RX_REG_ENTRIES = 96;
localparam TRIGGER_CONDITION_RX_CR_ADDR = 48'hC00;
localparam TRIGGER_CONDITION_RX_SIZE = 64;
localparam TRIGGER_CONDITION_RX_SRC_PORT_MASK_LO = 0;
localparam TRIGGER_CONDITION_RX_SRC_PORT_MASK_HI = 17;
localparam TRIGGER_CONDITION_RX_SRC_PORT_MASK_RESET = 18'h0;
localparam TRIGGER_CONDITION_RX_USEMASK = 64'h3FFFF;
localparam TRIGGER_CONDITION_RX_RO_MASK = 64'h0;
localparam TRIGGER_CONDITION_RX_WO_MASK = 64'h0;
localparam TRIGGER_CONDITION_RX_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [31:0] HANDLER_ACTION_MASK;  // RW
} TRIGGER_CONDITION_AMASK_1_t;

localparam TRIGGER_CONDITION_AMASK_1_REG_STRIDE = 48'h8;
localparam TRIGGER_CONDITION_AMASK_1_REG_ENTRIES = 96;
localparam TRIGGER_CONDITION_AMASK_1_CR_ADDR = 48'hF00;
localparam TRIGGER_CONDITION_AMASK_1_SIZE = 64;
localparam TRIGGER_CONDITION_AMASK_1_HANDLER_ACTION_MASK_LO = 0;
localparam TRIGGER_CONDITION_AMASK_1_HANDLER_ACTION_MASK_HI = 31;
localparam TRIGGER_CONDITION_AMASK_1_HANDLER_ACTION_MASK_RESET = 32'h0;
localparam TRIGGER_CONDITION_AMASK_1_USEMASK = 64'hFFFFFFFF;
localparam TRIGGER_CONDITION_AMASK_1_RO_MASK = 64'h0;
localparam TRIGGER_CONDITION_AMASK_1_WO_MASK = 64'h0;
localparam TRIGGER_CONDITION_AMASK_1_RESET = 64'h0;

typedef struct packed {
    logic [50:0] reserved0;  // RSVD
    logic [12:0] HANDLER_ACTION_MASK;  // RW
} TRIGGER_CONDITION_AMASK_2_t;

localparam TRIGGER_CONDITION_AMASK_2_REG_STRIDE = 48'h8;
localparam TRIGGER_CONDITION_AMASK_2_REG_ENTRIES = 96;
localparam TRIGGER_CONDITION_AMASK_2_CR_ADDR = 48'h1200;
localparam TRIGGER_CONDITION_AMASK_2_SIZE = 64;
localparam TRIGGER_CONDITION_AMASK_2_HANDLER_ACTION_MASK_LO = 0;
localparam TRIGGER_CONDITION_AMASK_2_HANDLER_ACTION_MASK_HI = 12;
localparam TRIGGER_CONDITION_AMASK_2_HANDLER_ACTION_MASK_RESET = 13'h0;
localparam TRIGGER_CONDITION_AMASK_2_USEMASK = 64'h1FFF;
localparam TRIGGER_CONDITION_AMASK_2_RO_MASK = 64'h0;
localparam TRIGGER_CONDITION_AMASK_2_WO_MASK = 64'h0;
localparam TRIGGER_CONDITION_AMASK_2_RESET = 64'h0;

typedef struct packed {
    logic [34:0] reserved0;  // RSVD
    logic  [1:0] MIRRORING_ACTION3;  // RW
    logic  [1:0] MIRRORING_ACTION2;  // RW
    logic  [1:0] MIRRORING_ACTION1;  // RW
    logic  [1:0] MIRRORING_ACTION0;  // RW
    logic  [0:0] NO_MODIFY_ACTION;  // RW
    logic  [0:0] POLICER_ACTION;  // RW
    logic  [0:0] EGRESS_L3_DOMAIN_ACTION;  // RW
    logic  [0:0] EGRESS_L2_DOMAIN_ACTION;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [0:0] RATE_LIMIT_ACTION;  // RW
    logic  [1:0] LEARNING_ACTION;  // RW
    logic  [0:0] VLAN_ACTION;  // RW
    logic  [0:0] TC_ACTION;  // RW
    logic  [3:0] reserved2;  // RSVD
    logic  [1:0] TRAP_ACTION;  // RW
    logic  [1:0] FORWARDING_ACTION;  // RW
} TRIGGER_ACTION_CFG_1_t;

localparam TRIGGER_ACTION_CFG_1_REG_STRIDE = 48'h8;
localparam TRIGGER_ACTION_CFG_1_REG_ENTRIES = 96;
localparam TRIGGER_ACTION_CFG_1_CR_ADDR = 48'h1500;
localparam TRIGGER_ACTION_CFG_1_SIZE = 64;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION3_LO = 27;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION3_HI = 28;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION3_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION2_LO = 25;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION2_HI = 26;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION2_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION1_LO = 23;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION1_HI = 24;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION1_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION0_LO = 21;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION0_HI = 22;
localparam TRIGGER_ACTION_CFG_1_MIRRORING_ACTION0_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_1_NO_MODIFY_ACTION_LO = 20;
localparam TRIGGER_ACTION_CFG_1_NO_MODIFY_ACTION_HI = 20;
localparam TRIGGER_ACTION_CFG_1_NO_MODIFY_ACTION_RESET = 1'h0;
localparam TRIGGER_ACTION_CFG_1_POLICER_ACTION_LO = 19;
localparam TRIGGER_ACTION_CFG_1_POLICER_ACTION_HI = 19;
localparam TRIGGER_ACTION_CFG_1_POLICER_ACTION_RESET = 1'h0;
localparam TRIGGER_ACTION_CFG_1_EGRESS_L3_DOMAIN_ACTION_LO = 18;
localparam TRIGGER_ACTION_CFG_1_EGRESS_L3_DOMAIN_ACTION_HI = 18;
localparam TRIGGER_ACTION_CFG_1_EGRESS_L3_DOMAIN_ACTION_RESET = 1'h0;
localparam TRIGGER_ACTION_CFG_1_EGRESS_L2_DOMAIN_ACTION_LO = 17;
localparam TRIGGER_ACTION_CFG_1_EGRESS_L2_DOMAIN_ACTION_HI = 17;
localparam TRIGGER_ACTION_CFG_1_EGRESS_L2_DOMAIN_ACTION_RESET = 1'h0;
localparam TRIGGER_ACTION_CFG_1_RATE_LIMIT_ACTION_LO = 12;
localparam TRIGGER_ACTION_CFG_1_RATE_LIMIT_ACTION_HI = 12;
localparam TRIGGER_ACTION_CFG_1_RATE_LIMIT_ACTION_RESET = 1'h0;
localparam TRIGGER_ACTION_CFG_1_LEARNING_ACTION_LO = 10;
localparam TRIGGER_ACTION_CFG_1_LEARNING_ACTION_HI = 11;
localparam TRIGGER_ACTION_CFG_1_LEARNING_ACTION_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_1_VLAN_ACTION_LO = 9;
localparam TRIGGER_ACTION_CFG_1_VLAN_ACTION_HI = 9;
localparam TRIGGER_ACTION_CFG_1_VLAN_ACTION_RESET = 1'h0;
localparam TRIGGER_ACTION_CFG_1_TC_ACTION_LO = 8;
localparam TRIGGER_ACTION_CFG_1_TC_ACTION_HI = 8;
localparam TRIGGER_ACTION_CFG_1_TC_ACTION_RESET = 1'h0;
localparam TRIGGER_ACTION_CFG_1_TRAP_ACTION_LO = 2;
localparam TRIGGER_ACTION_CFG_1_TRAP_ACTION_HI = 3;
localparam TRIGGER_ACTION_CFG_1_TRAP_ACTION_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_1_FORWARDING_ACTION_LO = 0;
localparam TRIGGER_ACTION_CFG_1_FORWARDING_ACTION_HI = 1;
localparam TRIGGER_ACTION_CFG_1_FORWARDING_ACTION_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_1_USEMASK = 64'h1FFE1F0F;
localparam TRIGGER_ACTION_CFG_1_RO_MASK = 64'h0;
localparam TRIGGER_ACTION_CFG_1_WO_MASK = 64'h0;
localparam TRIGGER_ACTION_CFG_1_RESET = 64'h0;

typedef struct packed {
    logic [41:0] reserved0;  // RSVD
    logic  [2:0] TRAP_CODE;  // RW
    logic  [3:0] RATE_LIMIT_NUM;  // RW
    logic [11:0] NEW_EVID;  // RW
    logic  [2:0] NEW_TC;  // RW
} TRIGGER_ACTION_CFG_2_t;

localparam TRIGGER_ACTION_CFG_2_REG_STRIDE = 48'h8;
localparam TRIGGER_ACTION_CFG_2_REG_ENTRIES = 96;
localparam TRIGGER_ACTION_CFG_2_CR_ADDR = 48'h1800;
localparam TRIGGER_ACTION_CFG_2_SIZE = 64;
localparam TRIGGER_ACTION_CFG_2_TRAP_CODE_LO = 19;
localparam TRIGGER_ACTION_CFG_2_TRAP_CODE_HI = 21;
localparam TRIGGER_ACTION_CFG_2_TRAP_CODE_RESET = 2'h0;
localparam TRIGGER_ACTION_CFG_2_RATE_LIMIT_NUM_LO = 15;
localparam TRIGGER_ACTION_CFG_2_RATE_LIMIT_NUM_HI = 18;
localparam TRIGGER_ACTION_CFG_2_RATE_LIMIT_NUM_RESET = 4'h0;
localparam TRIGGER_ACTION_CFG_2_NEW_EVID_LO = 3;
localparam TRIGGER_ACTION_CFG_2_NEW_EVID_HI = 14;
localparam TRIGGER_ACTION_CFG_2_NEW_EVID_RESET = 12'h0;
localparam TRIGGER_ACTION_CFG_2_NEW_TC_LO = 0;
localparam TRIGGER_ACTION_CFG_2_NEW_TC_HI = 2;
localparam TRIGGER_ACTION_CFG_2_NEW_TC_RESET = 3'h0;
localparam TRIGGER_ACTION_CFG_2_USEMASK = 64'h3FFFFF;
localparam TRIGGER_ACTION_CFG_2_RO_MASK = 64'h0;
localparam TRIGGER_ACTION_CFG_2_WO_MASK = 64'h0;
localparam TRIGGER_ACTION_CFG_2_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [15:0] NEW_DEST_GLORT_MASK;  // RW
    logic [15:0] NEW_DEST_GLORT;  // RW
} TRIGGER_ACTION_GLORT_t;

localparam TRIGGER_ACTION_GLORT_REG_STRIDE = 48'h8;
localparam TRIGGER_ACTION_GLORT_REG_ENTRIES = 96;
localparam TRIGGER_ACTION_GLORT_CR_ADDR = 48'h1B00;
localparam TRIGGER_ACTION_GLORT_SIZE = 64;
localparam TRIGGER_ACTION_GLORT_NEW_DEST_GLORT_MASK_LO = 16;
localparam TRIGGER_ACTION_GLORT_NEW_DEST_GLORT_MASK_HI = 31;
localparam TRIGGER_ACTION_GLORT_NEW_DEST_GLORT_MASK_RESET = 16'h0;
localparam TRIGGER_ACTION_GLORT_NEW_DEST_GLORT_LO = 0;
localparam TRIGGER_ACTION_GLORT_NEW_DEST_GLORT_HI = 15;
localparam TRIGGER_ACTION_GLORT_NEW_DEST_GLORT_RESET = 16'h0;
localparam TRIGGER_ACTION_GLORT_USEMASK = 64'hFFFFFFFF;
localparam TRIGGER_ACTION_GLORT_RO_MASK = 64'h0;
localparam TRIGGER_ACTION_GLORT_WO_MASK = 64'h0;
localparam TRIGGER_ACTION_GLORT_RESET = 64'h0;

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic  [5:0] MIRROR_PROFILE_INDEX3;  // RW
    logic  [5:0] MIRROR_PROFILE_INDEX2;  // RW
    logic  [5:0] MIRROR_PROFILE_INDEX1;  // RW
    logic  [5:0] MIRROR_PROFILE_INDEX0;  // RW
} TRIGGER_ACTION_MIRROR_t;

localparam TRIGGER_ACTION_MIRROR_REG_STRIDE = 48'h8;
localparam TRIGGER_ACTION_MIRROR_REG_ENTRIES = 96;
localparam TRIGGER_ACTION_MIRROR_CR_ADDR = 48'h1E00;
localparam TRIGGER_ACTION_MIRROR_SIZE = 64;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX3_LO = 18;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX3_HI = 23;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX3_RESET = 6'h0;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX2_LO = 12;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX2_HI = 17;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX2_RESET = 6'h0;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX1_LO = 6;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX1_HI = 11;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX1_RESET = 6'h0;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX0_LO = 0;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX0_HI = 5;
localparam TRIGGER_ACTION_MIRROR_MIRROR_PROFILE_INDEX0_RESET = 6'h0;
localparam TRIGGER_ACTION_MIRROR_USEMASK = 64'hFFFFFF;
localparam TRIGGER_ACTION_MIRROR_RO_MASK = 64'h0;
localparam TRIGGER_ACTION_MIRROR_WO_MASK = 64'h0;
localparam TRIGGER_ACTION_MIRROR_RESET = 64'h0;

typedef struct packed {
    logic [63:0] COUNT;  // RW/V
} TRIGGER_STATS_t;

localparam TRIGGER_STATS_REG_STRIDE = 48'h8;
localparam TRIGGER_STATS_REG_ENTRIES = 96;
localparam TRIGGER_STATS_CR_ADDR = 48'h2100;
localparam TRIGGER_STATS_SIZE = 64;
localparam TRIGGER_STATS_COUNT_LO = 0;
localparam TRIGGER_STATS_COUNT_HI = 63;
localparam TRIGGER_STATS_COUNT_RESET = 64'h0;
localparam TRIGGER_STATS_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_STATS_RO_MASK = 64'h0;
localparam TRIGGER_STATS_WO_MASK = 64'h0;
localparam TRIGGER_STATS_RESET = 64'h0;

typedef struct packed {
    logic  [0:0] GO_COMPL;  // RW/V
    logic  [0:0] STATUS;  // RW/V
    logic  [0:0] OP_TYPE;  // RW
    logic [12:0] reserved0;  // RSVD
    logic  [7:0] REG_ID;  // RW
    logic  [7:0] REG_SUB_ID;  // RW
    logic [31:0] REG_INDX;  // RW
} TRIGGER_DIRECT_MAP_CTRL_t;

localparam TRIGGER_DIRECT_MAP_CTRL_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_CTRL_CR_ADDR = 48'h2400;
localparam TRIGGER_DIRECT_MAP_CTRL_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_CTRL_GO_COMPL_LO = 63;
localparam TRIGGER_DIRECT_MAP_CTRL_GO_COMPL_HI = 63;
localparam TRIGGER_DIRECT_MAP_CTRL_GO_COMPL_RESET = 1'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_STATUS_LO = 62;
localparam TRIGGER_DIRECT_MAP_CTRL_STATUS_HI = 62;
localparam TRIGGER_DIRECT_MAP_CTRL_STATUS_RESET = 1'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_OP_TYPE_LO = 61;
localparam TRIGGER_DIRECT_MAP_CTRL_OP_TYPE_HI = 61;
localparam TRIGGER_DIRECT_MAP_CTRL_OP_TYPE_RESET = 1'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_ID_LO = 40;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_ID_HI = 47;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_ID_RESET = 8'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_SUB_ID_LO = 32;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_SUB_ID_HI = 39;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_SUB_ID_RESET = 8'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_INDX_LO = 0;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_INDX_HI = 31;
localparam TRIGGER_DIRECT_MAP_CTRL_REG_INDX_RESET = 32'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_USEMASK = 64'hE000FFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_CTRL_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTRL_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_PORT_MASK;  // RW
} TRIGGER_DIRECT_MAP_CTX0_t;

localparam TRIGGER_DIRECT_MAP_CTX0_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_CTX0_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_CTX0_CR_ADDR = 48'h2408;
localparam TRIGGER_DIRECT_MAP_CTX0_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_CTX0_DEST_PORT_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_CTX0_DEST_PORT_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_CTX0_DEST_PORT_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX0_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_CTX0_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX0_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX0_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_PORT_MASK;  // RW
} TRIGGER_DIRECT_MAP_CTX1_t;

localparam TRIGGER_DIRECT_MAP_CTX1_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_CTX1_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_CTX1_CR_ADDR = 48'h2410;
localparam TRIGGER_DIRECT_MAP_CTX1_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_CTX1_DEST_PORT_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_CTX1_DEST_PORT_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_CTX1_DEST_PORT_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX1_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_CTX1_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX1_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX1_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_PORT_MASK;  // RW
} TRIGGER_DIRECT_MAP_CTX2_t;

localparam TRIGGER_DIRECT_MAP_CTX2_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_CTX2_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_CTX2_CR_ADDR = 48'h2418;
localparam TRIGGER_DIRECT_MAP_CTX2_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_CTX2_DEST_PORT_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_CTX2_DEST_PORT_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_CTX2_DEST_PORT_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX2_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_CTX2_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX2_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX2_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_PORT_MASK;  // RW
} TRIGGER_DIRECT_MAP_CTX3_t;

localparam TRIGGER_DIRECT_MAP_CTX3_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_CTX3_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_CTX3_CR_ADDR = 48'h2420;
localparam TRIGGER_DIRECT_MAP_CTX3_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_CTX3_DEST_PORT_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_CTX3_DEST_PORT_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_CTX3_DEST_PORT_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX3_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_CTX3_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX3_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX3_RESET = 64'h0;

typedef struct packed {
    logic [61:0] reserved0;  // RSVD
    logic  [1:0] DEST_PORT_MASK;  // RW
} TRIGGER_DIRECT_MAP_CTX4_t;

localparam TRIGGER_DIRECT_MAP_CTX4_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_CTX4_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_CTX4_CR_ADDR = 48'h2428;
localparam TRIGGER_DIRECT_MAP_CTX4_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_CTX4_DEST_PORT_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_CTX4_DEST_PORT_MASK_HI = 1;
localparam TRIGGER_DIRECT_MAP_CTX4_DEST_PORT_MASK_RESET = 2'h0;
localparam TRIGGER_DIRECT_MAP_CTX4_USEMASK = 64'h3;
localparam TRIGGER_DIRECT_MAP_CTX4_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX4_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_CTX4_RESET = 64'h0;

typedef struct packed {
    logic [63:0] NEW_DEST_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADM0_t;

localparam TRIGGER_DIRECT_MAP_ADM0_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADM0_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADM0_CR_ADDR = 48'h2430;
localparam TRIGGER_DIRECT_MAP_ADM0_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADM0_NEW_DEST_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADM0_NEW_DEST_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADM0_NEW_DEST_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM0_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADM0_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM0_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM0_RESET = 64'h0;

typedef struct packed {
    logic [63:0] NEW_DEST_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADM1_t;

localparam TRIGGER_DIRECT_MAP_ADM1_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADM1_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADM1_CR_ADDR = 48'h2438;
localparam TRIGGER_DIRECT_MAP_ADM1_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADM1_NEW_DEST_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADM1_NEW_DEST_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADM1_NEW_DEST_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM1_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADM1_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM1_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM1_RESET = 64'h0;

typedef struct packed {
    logic [63:0] NEW_DEST_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADM2_t;

localparam TRIGGER_DIRECT_MAP_ADM2_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADM2_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADM2_CR_ADDR = 48'h2440;
localparam TRIGGER_DIRECT_MAP_ADM2_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADM2_NEW_DEST_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADM2_NEW_DEST_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADM2_NEW_DEST_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM2_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADM2_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM2_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM2_RESET = 64'h0;

typedef struct packed {
    logic [63:0] NEW_DEST_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADM3_t;

localparam TRIGGER_DIRECT_MAP_ADM3_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADM3_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADM3_CR_ADDR = 48'h2448;
localparam TRIGGER_DIRECT_MAP_ADM3_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADM3_NEW_DEST_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADM3_NEW_DEST_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADM3_NEW_DEST_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM3_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADM3_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM3_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM3_RESET = 64'h0;

typedef struct packed {
    logic [60:0] reserved0;  // RSVD
    logic  [0:0] FILTER_DEST_MASK;  // RW
    logic  [1:0] NEW_DEST_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADM4_t;

localparam TRIGGER_DIRECT_MAP_ADM4_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADM4_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADM4_CR_ADDR = 48'h2450;
localparam TRIGGER_DIRECT_MAP_ADM4_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADM4_FILTER_DEST_MASK_LO = 2;
localparam TRIGGER_DIRECT_MAP_ADM4_FILTER_DEST_MASK_HI = 2;
localparam TRIGGER_DIRECT_MAP_ADM4_FILTER_DEST_MASK_RESET = 1'h1;
localparam TRIGGER_DIRECT_MAP_ADM4_NEW_DEST_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADM4_NEW_DEST_MASK_HI = 1;
localparam TRIGGER_DIRECT_MAP_ADM4_NEW_DEST_MASK_RESET = 2'h0;
localparam TRIGGER_DIRECT_MAP_ADM4_USEMASK = 64'h7;
localparam TRIGGER_DIRECT_MAP_ADM4_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM4_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADM4_RESET = 64'h4;

typedef struct packed {
    logic [63:0] DROP_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADR0_t;

localparam TRIGGER_DIRECT_MAP_ADR0_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADR0_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADR0_CR_ADDR = 48'h2458;
localparam TRIGGER_DIRECT_MAP_ADR0_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADR0_DROP_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADR0_DROP_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADR0_DROP_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR0_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADR0_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR0_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR0_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DROP_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADR1_t;

localparam TRIGGER_DIRECT_MAP_ADR1_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADR1_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADR1_CR_ADDR = 48'h2460;
localparam TRIGGER_DIRECT_MAP_ADR1_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADR1_DROP_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADR1_DROP_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADR1_DROP_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR1_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADR1_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR1_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR1_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DROP_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADR2_t;

localparam TRIGGER_DIRECT_MAP_ADR2_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADR2_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADR2_CR_ADDR = 48'h2468;
localparam TRIGGER_DIRECT_MAP_ADR2_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADR2_DROP_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADR2_DROP_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADR2_DROP_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR2_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADR2_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR2_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR2_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DROP_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADR3_t;

localparam TRIGGER_DIRECT_MAP_ADR3_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADR3_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADR3_CR_ADDR = 48'h2470;
localparam TRIGGER_DIRECT_MAP_ADR3_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADR3_DROP_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADR3_DROP_MASK_HI = 63;
localparam TRIGGER_DIRECT_MAP_ADR3_DROP_MASK_RESET = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR3_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam TRIGGER_DIRECT_MAP_ADR3_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR3_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR3_RESET = 64'h0;

typedef struct packed {
    logic [61:0] reserved0;  // RSVD
    logic  [1:0] DROP_MASK;  // RW
} TRIGGER_DIRECT_MAP_ADR4_t;

localparam TRIGGER_DIRECT_MAP_ADR4_REG_STRIDE = 48'h8;
localparam TRIGGER_DIRECT_MAP_ADR4_REG_ENTRIES = 1;
localparam TRIGGER_DIRECT_MAP_ADR4_CR_ADDR = 48'h2478;
localparam TRIGGER_DIRECT_MAP_ADR4_SIZE = 64;
localparam TRIGGER_DIRECT_MAP_ADR4_DROP_MASK_LO = 0;
localparam TRIGGER_DIRECT_MAP_ADR4_DROP_MASK_HI = 1;
localparam TRIGGER_DIRECT_MAP_ADR4_DROP_MASK_RESET = 2'h0;
localparam TRIGGER_DIRECT_MAP_ADR4_USEMASK = 64'h3;
localparam TRIGGER_DIRECT_MAP_ADR4_RO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR4_WO_MASK = 64'h0;
localparam TRIGGER_DIRECT_MAP_ADR4_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_TRIGGER_CONDITION_CFG_t;

typedef logic [7:0] we_TRIGGER_CONDITION_PARAM_t;

typedef logic [7:0] we_TRIGGER_CONDITION_CGRP_t;

typedef logic [7:0] we_TRIGGER_CONDITION_GLORT_t;

typedef logic [7:0] we_TRIGGER_CONDITION_RX_t;

typedef logic [7:0] we_TRIGGER_CONDITION_AMASK_1_t;

typedef logic [7:0] we_TRIGGER_CONDITION_AMASK_2_t;

typedef logic [7:0] we_TRIGGER_ACTION_CFG_1_t;

typedef logic [7:0] we_TRIGGER_ACTION_CFG_2_t;

typedef logic [7:0] we_TRIGGER_ACTION_GLORT_t;

typedef logic [7:0] we_TRIGGER_ACTION_MIRROR_t;

typedef logic [7:0] we_TRIGGER_STATS_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_CTRL_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_CTX0_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_CTX1_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_CTX2_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_CTX3_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_CTX4_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADM0_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADM1_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADM2_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADM3_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADM4_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADR0_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADR1_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADR2_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADR3_t;

typedef logic [7:0] we_TRIGGER_DIRECT_MAP_ADR4_t;

typedef struct packed {
    we_TRIGGER_CONDITION_CFG_t TRIGGER_CONDITION_CFG;
    we_TRIGGER_CONDITION_PARAM_t TRIGGER_CONDITION_PARAM;
    we_TRIGGER_CONDITION_CGRP_t TRIGGER_CONDITION_CGRP;
    we_TRIGGER_CONDITION_GLORT_t TRIGGER_CONDITION_GLORT;
    we_TRIGGER_CONDITION_RX_t TRIGGER_CONDITION_RX;
    we_TRIGGER_CONDITION_AMASK_1_t TRIGGER_CONDITION_AMASK_1;
    we_TRIGGER_CONDITION_AMASK_2_t TRIGGER_CONDITION_AMASK_2;
    we_TRIGGER_ACTION_CFG_1_t TRIGGER_ACTION_CFG_1;
    we_TRIGGER_ACTION_CFG_2_t TRIGGER_ACTION_CFG_2;
    we_TRIGGER_ACTION_GLORT_t TRIGGER_ACTION_GLORT;
    we_TRIGGER_ACTION_MIRROR_t TRIGGER_ACTION_MIRROR;
    we_TRIGGER_STATS_t TRIGGER_STATS;
    we_TRIGGER_DIRECT_MAP_CTRL_t TRIGGER_DIRECT_MAP_CTRL;
    we_TRIGGER_DIRECT_MAP_CTX0_t TRIGGER_DIRECT_MAP_CTX0;
    we_TRIGGER_DIRECT_MAP_CTX1_t TRIGGER_DIRECT_MAP_CTX1;
    we_TRIGGER_DIRECT_MAP_CTX2_t TRIGGER_DIRECT_MAP_CTX2;
    we_TRIGGER_DIRECT_MAP_CTX3_t TRIGGER_DIRECT_MAP_CTX3;
    we_TRIGGER_DIRECT_MAP_CTX4_t TRIGGER_DIRECT_MAP_CTX4;
    we_TRIGGER_DIRECT_MAP_ADM0_t TRIGGER_DIRECT_MAP_ADM0;
    we_TRIGGER_DIRECT_MAP_ADM1_t TRIGGER_DIRECT_MAP_ADM1;
    we_TRIGGER_DIRECT_MAP_ADM2_t TRIGGER_DIRECT_MAP_ADM2;
    we_TRIGGER_DIRECT_MAP_ADM3_t TRIGGER_DIRECT_MAP_ADM3;
    we_TRIGGER_DIRECT_MAP_ADM4_t TRIGGER_DIRECT_MAP_ADM4;
    we_TRIGGER_DIRECT_MAP_ADR0_t TRIGGER_DIRECT_MAP_ADR0;
    we_TRIGGER_DIRECT_MAP_ADR1_t TRIGGER_DIRECT_MAP_ADR1;
    we_TRIGGER_DIRECT_MAP_ADR2_t TRIGGER_DIRECT_MAP_ADR2;
    we_TRIGGER_DIRECT_MAP_ADR3_t TRIGGER_DIRECT_MAP_ADR3;
    we_TRIGGER_DIRECT_MAP_ADR4_t TRIGGER_DIRECT_MAP_ADR4;
} mby_ppe_trig_apply_map_handcoded_t;

typedef logic [7:0] re_TRIGGER_CONDITION_CFG_t;

typedef logic [7:0] re_TRIGGER_CONDITION_PARAM_t;

typedef logic [7:0] re_TRIGGER_CONDITION_CGRP_t;

typedef logic [7:0] re_TRIGGER_CONDITION_GLORT_t;

typedef logic [7:0] re_TRIGGER_CONDITION_RX_t;

typedef logic [7:0] re_TRIGGER_CONDITION_AMASK_1_t;

typedef logic [7:0] re_TRIGGER_CONDITION_AMASK_2_t;

typedef logic [7:0] re_TRIGGER_ACTION_CFG_1_t;

typedef logic [7:0] re_TRIGGER_ACTION_CFG_2_t;

typedef logic [7:0] re_TRIGGER_ACTION_GLORT_t;

typedef logic [7:0] re_TRIGGER_ACTION_MIRROR_t;

typedef logic [7:0] re_TRIGGER_STATS_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_CTRL_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_CTX0_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_CTX1_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_CTX2_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_CTX3_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_CTX4_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADM0_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADM1_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADM2_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADM3_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADM4_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADR0_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADR1_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADR2_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADR3_t;

typedef logic [7:0] re_TRIGGER_DIRECT_MAP_ADR4_t;

typedef struct packed {
    re_TRIGGER_CONDITION_CFG_t TRIGGER_CONDITION_CFG;
    re_TRIGGER_CONDITION_PARAM_t TRIGGER_CONDITION_PARAM;
    re_TRIGGER_CONDITION_CGRP_t TRIGGER_CONDITION_CGRP;
    re_TRIGGER_CONDITION_GLORT_t TRIGGER_CONDITION_GLORT;
    re_TRIGGER_CONDITION_RX_t TRIGGER_CONDITION_RX;
    re_TRIGGER_CONDITION_AMASK_1_t TRIGGER_CONDITION_AMASK_1;
    re_TRIGGER_CONDITION_AMASK_2_t TRIGGER_CONDITION_AMASK_2;
    re_TRIGGER_ACTION_CFG_1_t TRIGGER_ACTION_CFG_1;
    re_TRIGGER_ACTION_CFG_2_t TRIGGER_ACTION_CFG_2;
    re_TRIGGER_ACTION_GLORT_t TRIGGER_ACTION_GLORT;
    re_TRIGGER_ACTION_MIRROR_t TRIGGER_ACTION_MIRROR;
    re_TRIGGER_STATS_t TRIGGER_STATS;
    re_TRIGGER_DIRECT_MAP_CTRL_t TRIGGER_DIRECT_MAP_CTRL;
    re_TRIGGER_DIRECT_MAP_CTX0_t TRIGGER_DIRECT_MAP_CTX0;
    re_TRIGGER_DIRECT_MAP_CTX1_t TRIGGER_DIRECT_MAP_CTX1;
    re_TRIGGER_DIRECT_MAP_CTX2_t TRIGGER_DIRECT_MAP_CTX2;
    re_TRIGGER_DIRECT_MAP_CTX3_t TRIGGER_DIRECT_MAP_CTX3;
    re_TRIGGER_DIRECT_MAP_CTX4_t TRIGGER_DIRECT_MAP_CTX4;
    re_TRIGGER_DIRECT_MAP_ADM0_t TRIGGER_DIRECT_MAP_ADM0;
    re_TRIGGER_DIRECT_MAP_ADM1_t TRIGGER_DIRECT_MAP_ADM1;
    re_TRIGGER_DIRECT_MAP_ADM2_t TRIGGER_DIRECT_MAP_ADM2;
    re_TRIGGER_DIRECT_MAP_ADM3_t TRIGGER_DIRECT_MAP_ADM3;
    re_TRIGGER_DIRECT_MAP_ADM4_t TRIGGER_DIRECT_MAP_ADM4;
    re_TRIGGER_DIRECT_MAP_ADR0_t TRIGGER_DIRECT_MAP_ADR0;
    re_TRIGGER_DIRECT_MAP_ADR1_t TRIGGER_DIRECT_MAP_ADR1;
    re_TRIGGER_DIRECT_MAP_ADR2_t TRIGGER_DIRECT_MAP_ADR2;
    re_TRIGGER_DIRECT_MAP_ADR3_t TRIGGER_DIRECT_MAP_ADR3;
    re_TRIGGER_DIRECT_MAP_ADR4_t TRIGGER_DIRECT_MAP_ADR4;
} mby_ppe_trig_apply_map_hc_re_t;

typedef logic handcode_rvalid_TRIGGER_CONDITION_CFG_t;

typedef logic handcode_rvalid_TRIGGER_CONDITION_PARAM_t;

typedef logic handcode_rvalid_TRIGGER_CONDITION_CGRP_t;

typedef logic handcode_rvalid_TRIGGER_CONDITION_GLORT_t;

typedef logic handcode_rvalid_TRIGGER_CONDITION_RX_t;

typedef logic handcode_rvalid_TRIGGER_CONDITION_AMASK_1_t;

typedef logic handcode_rvalid_TRIGGER_CONDITION_AMASK_2_t;

typedef logic handcode_rvalid_TRIGGER_ACTION_CFG_1_t;

typedef logic handcode_rvalid_TRIGGER_ACTION_CFG_2_t;

typedef logic handcode_rvalid_TRIGGER_ACTION_GLORT_t;

typedef logic handcode_rvalid_TRIGGER_ACTION_MIRROR_t;

typedef logic handcode_rvalid_TRIGGER_STATS_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_CTRL_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_CTX0_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_CTX1_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_CTX2_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_CTX3_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_CTX4_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADM0_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADM1_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADM2_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADM3_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADM4_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADR0_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADR1_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADR2_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADR3_t;

typedef logic handcode_rvalid_TRIGGER_DIRECT_MAP_ADR4_t;

typedef struct packed {
    handcode_rvalid_TRIGGER_CONDITION_CFG_t TRIGGER_CONDITION_CFG;
    handcode_rvalid_TRIGGER_CONDITION_PARAM_t TRIGGER_CONDITION_PARAM;
    handcode_rvalid_TRIGGER_CONDITION_CGRP_t TRIGGER_CONDITION_CGRP;
    handcode_rvalid_TRIGGER_CONDITION_GLORT_t TRIGGER_CONDITION_GLORT;
    handcode_rvalid_TRIGGER_CONDITION_RX_t TRIGGER_CONDITION_RX;
    handcode_rvalid_TRIGGER_CONDITION_AMASK_1_t TRIGGER_CONDITION_AMASK_1;
    handcode_rvalid_TRIGGER_CONDITION_AMASK_2_t TRIGGER_CONDITION_AMASK_2;
    handcode_rvalid_TRIGGER_ACTION_CFG_1_t TRIGGER_ACTION_CFG_1;
    handcode_rvalid_TRIGGER_ACTION_CFG_2_t TRIGGER_ACTION_CFG_2;
    handcode_rvalid_TRIGGER_ACTION_GLORT_t TRIGGER_ACTION_GLORT;
    handcode_rvalid_TRIGGER_ACTION_MIRROR_t TRIGGER_ACTION_MIRROR;
    handcode_rvalid_TRIGGER_STATS_t TRIGGER_STATS;
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTRL_t TRIGGER_DIRECT_MAP_CTRL;
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX0_t TRIGGER_DIRECT_MAP_CTX0;
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX1_t TRIGGER_DIRECT_MAP_CTX1;
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX2_t TRIGGER_DIRECT_MAP_CTX2;
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX3_t TRIGGER_DIRECT_MAP_CTX3;
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX4_t TRIGGER_DIRECT_MAP_CTX4;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM0_t TRIGGER_DIRECT_MAP_ADM0;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM1_t TRIGGER_DIRECT_MAP_ADM1;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM2_t TRIGGER_DIRECT_MAP_ADM2;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM3_t TRIGGER_DIRECT_MAP_ADM3;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM4_t TRIGGER_DIRECT_MAP_ADM4;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR0_t TRIGGER_DIRECT_MAP_ADR0;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR1_t TRIGGER_DIRECT_MAP_ADR1;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR2_t TRIGGER_DIRECT_MAP_ADR2;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR3_t TRIGGER_DIRECT_MAP_ADR3;
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR4_t TRIGGER_DIRECT_MAP_ADR4;
} mby_ppe_trig_apply_map_hc_rvalid_t;

typedef logic handcode_wvalid_TRIGGER_CONDITION_CFG_t;

typedef logic handcode_wvalid_TRIGGER_CONDITION_PARAM_t;

typedef logic handcode_wvalid_TRIGGER_CONDITION_CGRP_t;

typedef logic handcode_wvalid_TRIGGER_CONDITION_GLORT_t;

typedef logic handcode_wvalid_TRIGGER_CONDITION_RX_t;

typedef logic handcode_wvalid_TRIGGER_CONDITION_AMASK_1_t;

typedef logic handcode_wvalid_TRIGGER_CONDITION_AMASK_2_t;

typedef logic handcode_wvalid_TRIGGER_ACTION_CFG_1_t;

typedef logic handcode_wvalid_TRIGGER_ACTION_CFG_2_t;

typedef logic handcode_wvalid_TRIGGER_ACTION_GLORT_t;

typedef logic handcode_wvalid_TRIGGER_ACTION_MIRROR_t;

typedef logic handcode_wvalid_TRIGGER_STATS_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_CTRL_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_CTX0_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_CTX1_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_CTX2_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_CTX3_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_CTX4_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADM0_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADM1_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADM2_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADM3_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADM4_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADR0_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADR1_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADR2_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADR3_t;

typedef logic handcode_wvalid_TRIGGER_DIRECT_MAP_ADR4_t;

typedef struct packed {
    handcode_wvalid_TRIGGER_CONDITION_CFG_t TRIGGER_CONDITION_CFG;
    handcode_wvalid_TRIGGER_CONDITION_PARAM_t TRIGGER_CONDITION_PARAM;
    handcode_wvalid_TRIGGER_CONDITION_CGRP_t TRIGGER_CONDITION_CGRP;
    handcode_wvalid_TRIGGER_CONDITION_GLORT_t TRIGGER_CONDITION_GLORT;
    handcode_wvalid_TRIGGER_CONDITION_RX_t TRIGGER_CONDITION_RX;
    handcode_wvalid_TRIGGER_CONDITION_AMASK_1_t TRIGGER_CONDITION_AMASK_1;
    handcode_wvalid_TRIGGER_CONDITION_AMASK_2_t TRIGGER_CONDITION_AMASK_2;
    handcode_wvalid_TRIGGER_ACTION_CFG_1_t TRIGGER_ACTION_CFG_1;
    handcode_wvalid_TRIGGER_ACTION_CFG_2_t TRIGGER_ACTION_CFG_2;
    handcode_wvalid_TRIGGER_ACTION_GLORT_t TRIGGER_ACTION_GLORT;
    handcode_wvalid_TRIGGER_ACTION_MIRROR_t TRIGGER_ACTION_MIRROR;
    handcode_wvalid_TRIGGER_STATS_t TRIGGER_STATS;
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTRL_t TRIGGER_DIRECT_MAP_CTRL;
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX0_t TRIGGER_DIRECT_MAP_CTX0;
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX1_t TRIGGER_DIRECT_MAP_CTX1;
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX2_t TRIGGER_DIRECT_MAP_CTX2;
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX3_t TRIGGER_DIRECT_MAP_CTX3;
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX4_t TRIGGER_DIRECT_MAP_CTX4;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM0_t TRIGGER_DIRECT_MAP_ADM0;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM1_t TRIGGER_DIRECT_MAP_ADM1;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM2_t TRIGGER_DIRECT_MAP_ADM2;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM3_t TRIGGER_DIRECT_MAP_ADM3;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM4_t TRIGGER_DIRECT_MAP_ADM4;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR0_t TRIGGER_DIRECT_MAP_ADR0;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR1_t TRIGGER_DIRECT_MAP_ADR1;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR2_t TRIGGER_DIRECT_MAP_ADR2;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR3_t TRIGGER_DIRECT_MAP_ADR3;
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR4_t TRIGGER_DIRECT_MAP_ADR4;
} mby_ppe_trig_apply_map_hc_wvalid_t;

typedef logic handcode_error_TRIGGER_CONDITION_CFG_t;

typedef logic handcode_error_TRIGGER_CONDITION_PARAM_t;

typedef logic handcode_error_TRIGGER_CONDITION_CGRP_t;

typedef logic handcode_error_TRIGGER_CONDITION_GLORT_t;

typedef logic handcode_error_TRIGGER_CONDITION_RX_t;

typedef logic handcode_error_TRIGGER_CONDITION_AMASK_1_t;

typedef logic handcode_error_TRIGGER_CONDITION_AMASK_2_t;

typedef logic handcode_error_TRIGGER_ACTION_CFG_1_t;

typedef logic handcode_error_TRIGGER_ACTION_CFG_2_t;

typedef logic handcode_error_TRIGGER_ACTION_GLORT_t;

typedef logic handcode_error_TRIGGER_ACTION_MIRROR_t;

typedef logic handcode_error_TRIGGER_STATS_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_CTRL_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_CTX0_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_CTX1_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_CTX2_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_CTX3_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_CTX4_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADM0_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADM1_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADM2_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADM3_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADM4_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADR0_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADR1_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADR2_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADR3_t;

typedef logic handcode_error_TRIGGER_DIRECT_MAP_ADR4_t;

typedef struct packed {
    handcode_error_TRIGGER_CONDITION_CFG_t TRIGGER_CONDITION_CFG;
    handcode_error_TRIGGER_CONDITION_PARAM_t TRIGGER_CONDITION_PARAM;
    handcode_error_TRIGGER_CONDITION_CGRP_t TRIGGER_CONDITION_CGRP;
    handcode_error_TRIGGER_CONDITION_GLORT_t TRIGGER_CONDITION_GLORT;
    handcode_error_TRIGGER_CONDITION_RX_t TRIGGER_CONDITION_RX;
    handcode_error_TRIGGER_CONDITION_AMASK_1_t TRIGGER_CONDITION_AMASK_1;
    handcode_error_TRIGGER_CONDITION_AMASK_2_t TRIGGER_CONDITION_AMASK_2;
    handcode_error_TRIGGER_ACTION_CFG_1_t TRIGGER_ACTION_CFG_1;
    handcode_error_TRIGGER_ACTION_CFG_2_t TRIGGER_ACTION_CFG_2;
    handcode_error_TRIGGER_ACTION_GLORT_t TRIGGER_ACTION_GLORT;
    handcode_error_TRIGGER_ACTION_MIRROR_t TRIGGER_ACTION_MIRROR;
    handcode_error_TRIGGER_STATS_t TRIGGER_STATS;
    handcode_error_TRIGGER_DIRECT_MAP_CTRL_t TRIGGER_DIRECT_MAP_CTRL;
    handcode_error_TRIGGER_DIRECT_MAP_CTX0_t TRIGGER_DIRECT_MAP_CTX0;
    handcode_error_TRIGGER_DIRECT_MAP_CTX1_t TRIGGER_DIRECT_MAP_CTX1;
    handcode_error_TRIGGER_DIRECT_MAP_CTX2_t TRIGGER_DIRECT_MAP_CTX2;
    handcode_error_TRIGGER_DIRECT_MAP_CTX3_t TRIGGER_DIRECT_MAP_CTX3;
    handcode_error_TRIGGER_DIRECT_MAP_CTX4_t TRIGGER_DIRECT_MAP_CTX4;
    handcode_error_TRIGGER_DIRECT_MAP_ADM0_t TRIGGER_DIRECT_MAP_ADM0;
    handcode_error_TRIGGER_DIRECT_MAP_ADM1_t TRIGGER_DIRECT_MAP_ADM1;
    handcode_error_TRIGGER_DIRECT_MAP_ADM2_t TRIGGER_DIRECT_MAP_ADM2;
    handcode_error_TRIGGER_DIRECT_MAP_ADM3_t TRIGGER_DIRECT_MAP_ADM3;
    handcode_error_TRIGGER_DIRECT_MAP_ADM4_t TRIGGER_DIRECT_MAP_ADM4;
    handcode_error_TRIGGER_DIRECT_MAP_ADR0_t TRIGGER_DIRECT_MAP_ADR0;
    handcode_error_TRIGGER_DIRECT_MAP_ADR1_t TRIGGER_DIRECT_MAP_ADR1;
    handcode_error_TRIGGER_DIRECT_MAP_ADR2_t TRIGGER_DIRECT_MAP_ADR2;
    handcode_error_TRIGGER_DIRECT_MAP_ADR3_t TRIGGER_DIRECT_MAP_ADR3;
    handcode_error_TRIGGER_DIRECT_MAP_ADR4_t TRIGGER_DIRECT_MAP_ADR4;
} mby_ppe_trig_apply_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    TRIGGER_CONDITION_CFG_t TRIGGER_CONDITION_CFG;
    TRIGGER_CONDITION_PARAM_t TRIGGER_CONDITION_PARAM;
    TRIGGER_CONDITION_CGRP_t TRIGGER_CONDITION_CGRP;
    TRIGGER_CONDITION_GLORT_t TRIGGER_CONDITION_GLORT;
    TRIGGER_CONDITION_RX_t TRIGGER_CONDITION_RX;
    TRIGGER_CONDITION_AMASK_1_t TRIGGER_CONDITION_AMASK_1;
    TRIGGER_CONDITION_AMASK_2_t TRIGGER_CONDITION_AMASK_2;
    TRIGGER_ACTION_CFG_1_t TRIGGER_ACTION_CFG_1;
    TRIGGER_ACTION_CFG_2_t TRIGGER_ACTION_CFG_2;
    TRIGGER_ACTION_GLORT_t TRIGGER_ACTION_GLORT;
    TRIGGER_ACTION_MIRROR_t TRIGGER_ACTION_MIRROR;
    TRIGGER_STATS_t TRIGGER_STATS;
    TRIGGER_DIRECT_MAP_CTRL_t TRIGGER_DIRECT_MAP_CTRL;
    TRIGGER_DIRECT_MAP_CTX0_t TRIGGER_DIRECT_MAP_CTX0;
    TRIGGER_DIRECT_MAP_CTX1_t TRIGGER_DIRECT_MAP_CTX1;
    TRIGGER_DIRECT_MAP_CTX2_t TRIGGER_DIRECT_MAP_CTX2;
    TRIGGER_DIRECT_MAP_CTX3_t TRIGGER_DIRECT_MAP_CTX3;
    TRIGGER_DIRECT_MAP_CTX4_t TRIGGER_DIRECT_MAP_CTX4;
    TRIGGER_DIRECT_MAP_ADM0_t TRIGGER_DIRECT_MAP_ADM0;
    TRIGGER_DIRECT_MAP_ADM1_t TRIGGER_DIRECT_MAP_ADM1;
    TRIGGER_DIRECT_MAP_ADM2_t TRIGGER_DIRECT_MAP_ADM2;
    TRIGGER_DIRECT_MAP_ADM3_t TRIGGER_DIRECT_MAP_ADM3;
    TRIGGER_DIRECT_MAP_ADM4_t TRIGGER_DIRECT_MAP_ADM4;
    TRIGGER_DIRECT_MAP_ADR0_t TRIGGER_DIRECT_MAP_ADR0;
    TRIGGER_DIRECT_MAP_ADR1_t TRIGGER_DIRECT_MAP_ADR1;
    TRIGGER_DIRECT_MAP_ADR2_t TRIGGER_DIRECT_MAP_ADR2;
    TRIGGER_DIRECT_MAP_ADR3_t TRIGGER_DIRECT_MAP_ADR3;
    TRIGGER_DIRECT_MAP_ADR4_t TRIGGER_DIRECT_MAP_ADR4;
} mby_ppe_trig_apply_map_hc_reg_read_t;

typedef struct packed {
    TRIGGER_CONDITION_CFG_t TRIGGER_CONDITION_CFG;
    TRIGGER_CONDITION_PARAM_t TRIGGER_CONDITION_PARAM;
    TRIGGER_CONDITION_CGRP_t TRIGGER_CONDITION_CGRP;
    TRIGGER_CONDITION_GLORT_t TRIGGER_CONDITION_GLORT;
    TRIGGER_CONDITION_RX_t TRIGGER_CONDITION_RX;
    TRIGGER_CONDITION_AMASK_1_t TRIGGER_CONDITION_AMASK_1;
    TRIGGER_CONDITION_AMASK_2_t TRIGGER_CONDITION_AMASK_2;
    TRIGGER_ACTION_CFG_1_t TRIGGER_ACTION_CFG_1;
    TRIGGER_ACTION_CFG_2_t TRIGGER_ACTION_CFG_2;
    TRIGGER_ACTION_GLORT_t TRIGGER_ACTION_GLORT;
    TRIGGER_ACTION_MIRROR_t TRIGGER_ACTION_MIRROR;
    TRIGGER_STATS_t TRIGGER_STATS;
    TRIGGER_DIRECT_MAP_CTRL_t TRIGGER_DIRECT_MAP_CTRL;
    TRIGGER_DIRECT_MAP_CTX0_t TRIGGER_DIRECT_MAP_CTX0;
    TRIGGER_DIRECT_MAP_CTX1_t TRIGGER_DIRECT_MAP_CTX1;
    TRIGGER_DIRECT_MAP_CTX2_t TRIGGER_DIRECT_MAP_CTX2;
    TRIGGER_DIRECT_MAP_CTX3_t TRIGGER_DIRECT_MAP_CTX3;
    TRIGGER_DIRECT_MAP_CTX4_t TRIGGER_DIRECT_MAP_CTX4;
    TRIGGER_DIRECT_MAP_ADM0_t TRIGGER_DIRECT_MAP_ADM0;
    TRIGGER_DIRECT_MAP_ADM1_t TRIGGER_DIRECT_MAP_ADM1;
    TRIGGER_DIRECT_MAP_ADM2_t TRIGGER_DIRECT_MAP_ADM2;
    TRIGGER_DIRECT_MAP_ADM3_t TRIGGER_DIRECT_MAP_ADM3;
    TRIGGER_DIRECT_MAP_ADM4_t TRIGGER_DIRECT_MAP_ADM4;
    TRIGGER_DIRECT_MAP_ADR0_t TRIGGER_DIRECT_MAP_ADR0;
    TRIGGER_DIRECT_MAP_ADR1_t TRIGGER_DIRECT_MAP_ADR1;
    TRIGGER_DIRECT_MAP_ADR2_t TRIGGER_DIRECT_MAP_ADR2;
    TRIGGER_DIRECT_MAP_ADR3_t TRIGGER_DIRECT_MAP_ADR3;
    TRIGGER_DIRECT_MAP_ADR4_t TRIGGER_DIRECT_MAP_ADR4;
} mby_ppe_trig_apply_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_trig_apply_map_pkg

`endif // MBY_PPE_TRIG_APPLY_MAP_PKG_VH
