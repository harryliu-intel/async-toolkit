magic
tech scmos
timestamp 965071231
<< ndiffusion >>
rect 160 141 168 142
rect 160 133 168 138
rect 130 117 146 118
rect 160 125 168 130
rect 160 117 168 122
rect 130 109 146 114
rect 160 109 168 114
rect 130 105 146 106
rect 130 97 138 105
rect 130 96 146 97
rect 160 105 168 106
rect 160 96 168 97
rect 130 88 146 93
rect 160 88 168 93
rect 130 84 146 85
rect 138 79 146 84
rect 160 80 168 85
rect 160 72 168 77
rect 138 65 146 70
rect 130 64 146 65
rect 160 64 168 69
rect 130 56 146 61
rect 160 60 168 61
rect 130 52 146 53
rect 130 44 132 52
rect 130 43 146 44
rect 130 39 146 40
<< pdiffusion >>
rect 198 163 214 164
rect 198 157 214 160
rect 220 149 224 154
rect 198 148 224 149
rect 229 149 233 154
rect 229 148 241 149
rect 198 144 224 145
rect 220 136 224 144
rect 198 135 224 136
rect 229 144 241 145
rect 237 136 241 144
rect 229 135 241 136
rect 198 131 224 132
rect 198 123 206 131
rect 198 122 224 123
rect 229 131 241 132
rect 229 123 233 131
rect 229 122 241 123
rect 198 118 224 119
rect 220 110 224 118
rect 198 109 224 110
rect 229 118 241 119
rect 237 110 241 118
rect 229 109 241 110
rect 198 105 224 106
rect 220 97 224 105
rect 198 96 224 97
rect 229 105 241 106
rect 229 97 233 105
rect 229 96 241 97
rect 198 92 224 93
rect 220 84 224 92
rect 198 83 224 84
rect 229 92 241 93
rect 237 84 241 92
rect 229 83 241 84
rect 198 79 224 80
rect 198 71 206 79
rect 198 70 224 71
rect 229 79 241 80
rect 229 71 233 79
rect 229 70 241 71
rect 198 66 224 67
rect 220 58 224 66
rect 198 57 224 58
rect 229 66 241 67
rect 237 58 241 66
rect 229 57 241 58
rect 198 53 224 54
rect 198 51 208 53
rect 191 46 208 51
rect 191 43 203 46
rect 229 53 241 54
rect 229 45 233 53
rect 229 43 241 45
rect 191 39 203 40
rect 229 39 241 40
<< ntransistor >>
rect 160 138 168 141
rect 160 130 168 133
rect 160 122 168 125
rect 130 114 146 117
rect 160 114 168 117
rect 130 106 146 109
rect 160 106 168 109
rect 130 93 146 96
rect 160 93 168 96
rect 130 85 146 88
rect 160 85 168 88
rect 160 77 168 80
rect 160 69 168 72
rect 130 61 146 64
rect 160 61 168 64
rect 130 53 146 56
rect 130 40 146 43
<< ptransistor >>
rect 198 160 214 163
rect 198 145 224 148
rect 229 145 241 148
rect 198 132 224 135
rect 229 132 241 135
rect 198 119 224 122
rect 229 119 241 122
rect 198 106 224 109
rect 229 106 241 109
rect 198 93 224 96
rect 229 93 241 96
rect 198 80 224 83
rect 229 80 241 83
rect 198 67 224 70
rect 229 67 241 70
rect 198 54 224 57
rect 229 54 241 57
rect 191 40 203 43
rect 229 40 241 43
<< polysilicon >>
rect 194 160 198 163
rect 214 160 218 163
rect 177 145 198 148
rect 224 145 229 148
rect 241 145 245 148
rect 156 138 160 141
rect 168 138 172 141
rect 177 133 180 145
rect 148 130 160 133
rect 168 130 180 133
rect 185 132 198 135
rect 224 132 229 135
rect 241 132 245 135
rect 148 117 151 130
rect 185 125 188 132
rect 156 122 160 125
rect 168 122 188 125
rect 193 119 198 122
rect 224 119 229 122
rect 241 119 245 122
rect 193 117 196 119
rect 126 114 130 117
rect 146 114 151 117
rect 156 114 160 117
rect 168 114 196 117
rect 126 106 130 109
rect 146 106 160 109
rect 168 106 198 109
rect 224 106 229 109
rect 241 106 245 109
rect 126 93 130 96
rect 146 93 160 96
rect 168 93 198 96
rect 224 93 229 96
rect 241 93 245 96
rect 126 85 130 88
rect 146 85 151 88
rect 156 85 160 88
rect 168 85 196 88
rect 148 72 151 85
rect 193 83 196 85
rect 193 80 198 83
rect 224 80 229 83
rect 241 80 245 83
rect 156 77 160 80
rect 168 77 188 80
rect 148 69 160 72
rect 168 69 180 72
rect 126 61 130 64
rect 146 61 160 64
rect 168 61 172 64
rect 128 53 130 56
rect 146 53 152 56
rect 177 57 180 69
rect 185 70 188 77
rect 185 67 198 70
rect 224 67 229 70
rect 241 67 245 70
rect 177 54 198 57
rect 224 54 229 57
rect 241 54 245 57
rect 126 40 130 43
rect 146 40 179 43
rect 187 40 191 43
rect 203 40 207 43
rect 217 41 229 43
rect 220 40 229 41
rect 241 40 245 43
<< ndcontact >>
rect 160 142 168 150
rect 130 118 146 126
rect 138 97 146 105
rect 160 97 168 105
rect 130 65 138 84
rect 160 52 168 60
rect 132 44 146 52
rect 130 31 146 39
<< pdcontact >>
rect 198 164 214 172
rect 198 149 220 157
rect 233 149 241 157
rect 198 136 220 144
rect 229 136 237 144
rect 206 123 224 131
rect 233 123 241 131
rect 198 110 220 118
rect 229 110 237 118
rect 198 97 220 105
rect 233 97 241 105
rect 198 84 220 92
rect 229 84 237 92
rect 206 71 224 79
rect 233 71 241 79
rect 198 58 220 66
rect 229 58 237 66
rect 208 45 224 53
rect 233 45 241 53
rect 191 31 203 39
rect 229 31 241 39
<< polycontact >>
rect 120 48 128 56
rect 179 40 187 48
rect 212 33 220 41
<< metal1 >>
rect 179 164 229 172
rect 160 142 168 150
rect 130 118 146 126
rect 130 84 134 118
rect 179 105 187 164
rect 198 149 220 157
rect 224 144 229 164
rect 233 153 241 157
rect 233 149 245 153
rect 198 136 220 144
rect 224 136 237 144
rect 198 118 202 136
rect 224 131 229 136
rect 241 131 245 149
rect 206 123 229 131
rect 233 123 245 131
rect 224 118 229 123
rect 198 110 220 118
rect 224 110 237 118
rect 138 97 187 105
rect 198 97 220 105
rect 130 65 138 84
rect 120 48 128 56
rect 160 52 168 60
rect 124 39 128 48
rect 132 44 168 52
rect 179 40 187 97
rect 224 92 229 110
rect 241 105 245 123
rect 233 97 245 105
rect 198 84 220 92
rect 224 84 237 92
rect 198 66 202 84
rect 224 79 229 84
rect 241 79 245 97
rect 206 71 229 79
rect 233 71 245 79
rect 224 66 229 71
rect 198 58 220 66
rect 224 62 237 66
rect 229 58 237 62
rect 241 53 245 71
rect 208 45 229 53
rect 233 49 245 53
rect 233 45 241 49
rect 212 39 220 41
rect 124 35 146 39
rect 191 35 220 39
rect 130 34 220 35
rect 130 31 203 34
rect 212 33 220 34
rect 224 39 229 45
rect 224 31 241 39
<< labels >>
rlabel metal1 202 153 202 153 5 Vdd!
rlabel metal1 202 101 202 101 1 Vdd!
rlabel metal1 164 101 164 101 1 x
rlabel metal1 142 101 142 101 1 x
rlabel metal1 164 146 164 146 5 GND!
rlabel polysilicon 159 139 159 139 1 _SReset!
rlabel metal1 164 56 164 56 1 GND!
rlabel metal1 142 48 142 48 1 GND!
rlabel polysilicon 129 62 129 62 1 _SReset!
rlabel metal1 220 127 220 127 1 x
rlabel pdcontact 220 75 220 75 5 x
rlabel metal1 237 35 237 35 1 Vdd!
rlabel polysilicon 242 55 242 55 1 _a0
rlabel polysilicon 242 68 242 68 1 _b0
rlabel polysilicon 242 81 242 81 1 _b1
rlabel polysilicon 242 94 242 94 1 _a1
rlabel polysilicon 242 107 242 107 1 _b0
rlabel polysilicon 242 120 242 120 1 _a0
rlabel polysilicon 242 133 242 133 1 _a1
rlabel polysilicon 242 146 242 146 1 _b1
rlabel metal1 215 49 215 49 1 Vdd!
rlabel metal1 203 168 203 168 5 x
rlabel polysilicon 215 161 215 161 1 _PReset!
rlabel space 125 59 160 150 7 ^n
rlabel space 119 30 153 58 7 ^n
rlabel space 211 30 246 61 3 ^p
rlabel space 219 62 246 170 3 ^p
<< end >>
