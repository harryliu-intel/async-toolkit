///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_mst_glort_map_pkg.vh                               
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_MST_GLORT_MAP_PKG_VH
`define MBY_PPE_MST_GLORT_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_mst_glort_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_mst_glort_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_mst_glort_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_mst_glort_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [63:0] MEMBERSHIP;  // RW
} EGRESS_VID_TABLE_t;

localparam EGRESS_VID_TABLE_REG_STRIDE = 48'h8;
localparam EGRESS_VID_TABLE_REG_ENTRIES = 5;
localparam EGRESS_VID_TABLE_REGFILE_STRIDE = 48'h40;
localparam EGRESS_VID_TABLE_REGFILE_ENTRIES = 4096;
localparam EGRESS_VID_TABLE_CR_ADDR = 48'h0;
localparam EGRESS_VID_TABLE_SIZE = 64;
localparam EGRESS_VID_TABLE_MEMBERSHIP_LO = 0;
localparam EGRESS_VID_TABLE_MEMBERSHIP_HI = 63;
localparam EGRESS_VID_TABLE_MEMBERSHIP_RESET = 64'h0;
localparam EGRESS_VID_TABLE_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam EGRESS_VID_TABLE_RO_MASK = 64'h0;
localparam EGRESS_VID_TABLE_WO_MASK = 64'h0;
localparam EGRESS_VID_TABLE_RESET = 64'h0;

typedef struct packed {
    logic [57:0] reserved0;  // RSVD
    logic  [5:0] TRIG_ID;  // RW
} EGRESS_VID_CFG_t;

localparam EGRESS_VID_CFG_REG_STRIDE = 48'h8;
localparam EGRESS_VID_CFG_REG_ENTRIES = 4096;
localparam EGRESS_VID_CFG_CR_ADDR = 48'h40000;
localparam EGRESS_VID_CFG_SIZE = 64;
localparam EGRESS_VID_CFG_TRIG_ID_LO = 0;
localparam EGRESS_VID_CFG_TRIG_ID_HI = 5;
localparam EGRESS_VID_CFG_TRIG_ID_RESET = 6'h0;
localparam EGRESS_VID_CFG_USEMASK = 64'h3F;
localparam EGRESS_VID_CFG_RO_MASK = 64'h0;
localparam EGRESS_VID_CFG_WO_MASK = 64'h0;
localparam EGRESS_VID_CFG_RESET = 64'h0;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic  [1:0] STP_STATE_17;  // RW
    logic  [1:0] STP_STATE_16;  // RW
    logic  [1:0] STP_STATE_15;  // RW
    logic  [1:0] STP_STATE_14;  // RW
    logic  [1:0] STP_STATE_13;  // RW
    logic  [1:0] STP_STATE_12;  // RW
    logic  [1:0] STP_STATE_11;  // RW
    logic  [1:0] STP_STATE_10;  // RW
    logic  [1:0] STP_STATE_9;  // RW
    logic  [1:0] STP_STATE_8;  // RW
    logic  [1:0] STP_STATE_7;  // RW
    logic  [1:0] STP_STATE_6;  // RW
    logic  [1:0] STP_STATE_5;  // RW
    logic  [1:0] STP_STATE_4;  // RW
    logic  [1:0] STP_STATE_3;  // RW
    logic  [1:0] STP_STATE_2;  // RW
    logic  [1:0] STP_STATE_1;  // RW
    logic  [1:0] STP_STATE_0;  // RW
} INGRESS_MST_TABLE_t;

localparam INGRESS_MST_TABLE_REG_STRIDE = 48'h8;
localparam INGRESS_MST_TABLE_REG_ENTRIES = 4096;
localparam INGRESS_MST_TABLE_CR_ADDR = 48'h48000;
localparam INGRESS_MST_TABLE_SIZE = 64;
localparam INGRESS_MST_TABLE_STP_STATE_17_LO = 34;
localparam INGRESS_MST_TABLE_STP_STATE_17_HI = 35;
localparam INGRESS_MST_TABLE_STP_STATE_17_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_16_LO = 32;
localparam INGRESS_MST_TABLE_STP_STATE_16_HI = 33;
localparam INGRESS_MST_TABLE_STP_STATE_16_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_15_LO = 30;
localparam INGRESS_MST_TABLE_STP_STATE_15_HI = 31;
localparam INGRESS_MST_TABLE_STP_STATE_15_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_14_LO = 28;
localparam INGRESS_MST_TABLE_STP_STATE_14_HI = 29;
localparam INGRESS_MST_TABLE_STP_STATE_14_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_13_LO = 26;
localparam INGRESS_MST_TABLE_STP_STATE_13_HI = 27;
localparam INGRESS_MST_TABLE_STP_STATE_13_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_12_LO = 24;
localparam INGRESS_MST_TABLE_STP_STATE_12_HI = 25;
localparam INGRESS_MST_TABLE_STP_STATE_12_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_11_LO = 22;
localparam INGRESS_MST_TABLE_STP_STATE_11_HI = 23;
localparam INGRESS_MST_TABLE_STP_STATE_11_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_10_LO = 20;
localparam INGRESS_MST_TABLE_STP_STATE_10_HI = 21;
localparam INGRESS_MST_TABLE_STP_STATE_10_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_9_LO = 18;
localparam INGRESS_MST_TABLE_STP_STATE_9_HI = 19;
localparam INGRESS_MST_TABLE_STP_STATE_9_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_8_LO = 16;
localparam INGRESS_MST_TABLE_STP_STATE_8_HI = 17;
localparam INGRESS_MST_TABLE_STP_STATE_8_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_7_LO = 14;
localparam INGRESS_MST_TABLE_STP_STATE_7_HI = 15;
localparam INGRESS_MST_TABLE_STP_STATE_7_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_6_LO = 12;
localparam INGRESS_MST_TABLE_STP_STATE_6_HI = 13;
localparam INGRESS_MST_TABLE_STP_STATE_6_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_5_LO = 10;
localparam INGRESS_MST_TABLE_STP_STATE_5_HI = 11;
localparam INGRESS_MST_TABLE_STP_STATE_5_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_4_LO = 8;
localparam INGRESS_MST_TABLE_STP_STATE_4_HI = 9;
localparam INGRESS_MST_TABLE_STP_STATE_4_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_3_LO = 6;
localparam INGRESS_MST_TABLE_STP_STATE_3_HI = 7;
localparam INGRESS_MST_TABLE_STP_STATE_3_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_2_LO = 4;
localparam INGRESS_MST_TABLE_STP_STATE_2_HI = 5;
localparam INGRESS_MST_TABLE_STP_STATE_2_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_1_LO = 2;
localparam INGRESS_MST_TABLE_STP_STATE_1_HI = 3;
localparam INGRESS_MST_TABLE_STP_STATE_1_RESET = 2'h0;
localparam INGRESS_MST_TABLE_STP_STATE_0_LO = 0;
localparam INGRESS_MST_TABLE_STP_STATE_0_HI = 1;
localparam INGRESS_MST_TABLE_STP_STATE_0_RESET = 2'h0;
localparam INGRESS_MST_TABLE_USEMASK = 64'hFFFFFFFFF;
localparam INGRESS_MST_TABLE_RO_MASK = 64'h0;
localparam INGRESS_MST_TABLE_WO_MASK = 64'h0;
localparam INGRESS_MST_TABLE_RESET = 64'h0;

typedef struct packed {
    logic [63:0] FORWARDING;  // RW
} EGRESS_MST_TABLE_t;

localparam EGRESS_MST_TABLE_REG_STRIDE = 48'h8;
localparam EGRESS_MST_TABLE_REG_ENTRIES = 5;
localparam EGRESS_MST_TABLE_REGFILE_STRIDE = 48'h40;
localparam EGRESS_MST_TABLE_REGFILE_ENTRIES = 4096;
localparam EGRESS_MST_TABLE_CR_ADDR = 48'h80000;
localparam EGRESS_MST_TABLE_SIZE = 64;
localparam EGRESS_MST_TABLE_FORWARDING_LO = 0;
localparam EGRESS_MST_TABLE_FORWARDING_HI = 63;
localparam EGRESS_MST_TABLE_FORWARDING_RESET = 64'h0;
localparam EGRESS_MST_TABLE_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam EGRESS_MST_TABLE_RO_MASK = 64'h0;
localparam EGRESS_MST_TABLE_WO_MASK = 64'h0;
localparam EGRESS_MST_TABLE_RESET = 64'h0;

typedef struct packed {
    logic  [0:0] GO_COMPL;  // RW/V
    logic  [0:0] STATUS;  // RW/V
    logic  [0:0] OP_TYPE;  // RW
    logic [12:0] reserved0;  // RSVD
    logic  [7:0] REG_ID;  // RW
    logic  [7:0] REG_SUB_ID;  // RW
    logic [31:0] REG_INDX;  // RW
} GLORT_DIRECT_MAP_CTRL_t;

localparam GLORT_DIRECT_MAP_CTRL_REG_STRIDE = 48'h8;
localparam GLORT_DIRECT_MAP_CTRL_REG_ENTRIES = 1;
localparam GLORT_DIRECT_MAP_CTRL_CR_ADDR = 48'hC0000;
localparam GLORT_DIRECT_MAP_CTRL_SIZE = 64;
localparam GLORT_DIRECT_MAP_CTRL_GO_COMPL_LO = 63;
localparam GLORT_DIRECT_MAP_CTRL_GO_COMPL_HI = 63;
localparam GLORT_DIRECT_MAP_CTRL_GO_COMPL_RESET = 1'h0;
localparam GLORT_DIRECT_MAP_CTRL_STATUS_LO = 62;
localparam GLORT_DIRECT_MAP_CTRL_STATUS_HI = 62;
localparam GLORT_DIRECT_MAP_CTRL_STATUS_RESET = 1'h0;
localparam GLORT_DIRECT_MAP_CTRL_OP_TYPE_LO = 61;
localparam GLORT_DIRECT_MAP_CTRL_OP_TYPE_HI = 61;
localparam GLORT_DIRECT_MAP_CTRL_OP_TYPE_RESET = 1'h0;
localparam GLORT_DIRECT_MAP_CTRL_REG_ID_LO = 40;
localparam GLORT_DIRECT_MAP_CTRL_REG_ID_HI = 47;
localparam GLORT_DIRECT_MAP_CTRL_REG_ID_RESET = 8'h0;
localparam GLORT_DIRECT_MAP_CTRL_REG_SUB_ID_LO = 32;
localparam GLORT_DIRECT_MAP_CTRL_REG_SUB_ID_HI = 39;
localparam GLORT_DIRECT_MAP_CTRL_REG_SUB_ID_RESET = 8'h0;
localparam GLORT_DIRECT_MAP_CTRL_REG_INDX_LO = 0;
localparam GLORT_DIRECT_MAP_CTRL_REG_INDX_HI = 31;
localparam GLORT_DIRECT_MAP_CTRL_REG_INDX_RESET = 32'h0;
localparam GLORT_DIRECT_MAP_CTRL_USEMASK = 64'hE000FFFFFFFFFFFF;
localparam GLORT_DIRECT_MAP_CTRL_RO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_CTRL_WO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_CTRL_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_MASK;  // RW
} GLORT_DIRECT_MAP_DST0_t;

localparam GLORT_DIRECT_MAP_DST0_REG_STRIDE = 48'h8;
localparam GLORT_DIRECT_MAP_DST0_REG_ENTRIES = 1;
localparam GLORT_DIRECT_MAP_DST0_CR_ADDR = 48'hC0008;
localparam GLORT_DIRECT_MAP_DST0_SIZE = 64;
localparam GLORT_DIRECT_MAP_DST0_DEST_MASK_LO = 0;
localparam GLORT_DIRECT_MAP_DST0_DEST_MASK_HI = 63;
localparam GLORT_DIRECT_MAP_DST0_DEST_MASK_RESET = 64'h0;
localparam GLORT_DIRECT_MAP_DST0_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam GLORT_DIRECT_MAP_DST0_RO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST0_WO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST0_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_MASK;  // RW
} GLORT_DIRECT_MAP_DST1_t;

localparam GLORT_DIRECT_MAP_DST1_REG_STRIDE = 48'h8;
localparam GLORT_DIRECT_MAP_DST1_REG_ENTRIES = 1;
localparam GLORT_DIRECT_MAP_DST1_CR_ADDR = 48'hC0010;
localparam GLORT_DIRECT_MAP_DST1_SIZE = 64;
localparam GLORT_DIRECT_MAP_DST1_DEST_MASK_LO = 0;
localparam GLORT_DIRECT_MAP_DST1_DEST_MASK_HI = 63;
localparam GLORT_DIRECT_MAP_DST1_DEST_MASK_RESET = 64'h0;
localparam GLORT_DIRECT_MAP_DST1_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam GLORT_DIRECT_MAP_DST1_RO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST1_WO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST1_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_MASK;  // RW
} GLORT_DIRECT_MAP_DST2_t;

localparam GLORT_DIRECT_MAP_DST2_REG_STRIDE = 48'h8;
localparam GLORT_DIRECT_MAP_DST2_REG_ENTRIES = 1;
localparam GLORT_DIRECT_MAP_DST2_CR_ADDR = 48'hC0018;
localparam GLORT_DIRECT_MAP_DST2_SIZE = 64;
localparam GLORT_DIRECT_MAP_DST2_DEST_MASK_LO = 0;
localparam GLORT_DIRECT_MAP_DST2_DEST_MASK_HI = 63;
localparam GLORT_DIRECT_MAP_DST2_DEST_MASK_RESET = 64'h0;
localparam GLORT_DIRECT_MAP_DST2_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam GLORT_DIRECT_MAP_DST2_RO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST2_WO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST2_RESET = 64'h0;

typedef struct packed {
    logic [63:0] DEST_MASK;  // RW
} GLORT_DIRECT_MAP_DST3_t;

localparam GLORT_DIRECT_MAP_DST3_REG_STRIDE = 48'h8;
localparam GLORT_DIRECT_MAP_DST3_REG_ENTRIES = 1;
localparam GLORT_DIRECT_MAP_DST3_CR_ADDR = 48'hC0020;
localparam GLORT_DIRECT_MAP_DST3_SIZE = 64;
localparam GLORT_DIRECT_MAP_DST3_DEST_MASK_LO = 0;
localparam GLORT_DIRECT_MAP_DST3_DEST_MASK_HI = 63;
localparam GLORT_DIRECT_MAP_DST3_DEST_MASK_RESET = 64'h0;
localparam GLORT_DIRECT_MAP_DST3_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam GLORT_DIRECT_MAP_DST3_RO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST3_WO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST3_RESET = 64'h0;

typedef struct packed {
    logic [49:0] reserved0;  // RSVD
    logic [11:0] IP_MULTICAST_INDEX;  // RW
    logic  [1:0] DEST_MASK;  // RW
} GLORT_DIRECT_MAP_DST4_t;

localparam GLORT_DIRECT_MAP_DST4_REG_STRIDE = 48'h8;
localparam GLORT_DIRECT_MAP_DST4_REG_ENTRIES = 1;
localparam GLORT_DIRECT_MAP_DST4_CR_ADDR = 48'hC0028;
localparam GLORT_DIRECT_MAP_DST4_SIZE = 64;
localparam GLORT_DIRECT_MAP_DST4_IP_MULTICAST_INDEX_LO = 2;
localparam GLORT_DIRECT_MAP_DST4_IP_MULTICAST_INDEX_HI = 13;
localparam GLORT_DIRECT_MAP_DST4_IP_MULTICAST_INDEX_RESET = 12'h0;
localparam GLORT_DIRECT_MAP_DST4_DEST_MASK_LO = 0;
localparam GLORT_DIRECT_MAP_DST4_DEST_MASK_HI = 1;
localparam GLORT_DIRECT_MAP_DST4_DEST_MASK_RESET = 2'h0;
localparam GLORT_DIRECT_MAP_DST4_USEMASK = 64'h3FFF;
localparam GLORT_DIRECT_MAP_DST4_RO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST4_WO_MASK = 64'h0;
localparam GLORT_DIRECT_MAP_DST4_RESET = 64'h0;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic  [0:0] SKIP_DGLORT_DEC;  // RW
    logic  [0:0] HASH_ROTATION;  // RW
    logic  [3:0] DEST_COUNT;  // RW
    logic  [7:0] RANGE_SUB_INDEX_B;  // RW
    logic  [7:0] RANGE_SUB_INDEX_A;  // RW
    logic [11:0] DEST_INDEX;  // RW
    logic  [1:0] STRICT;  // RW
} GLORT_RAM_t;

localparam GLORT_RAM_REG_STRIDE = 48'h8;
localparam GLORT_RAM_REG_ENTRIES = 64;
localparam GLORT_RAM_CR_ADDR = 48'hC0200;
localparam GLORT_RAM_SIZE = 64;
localparam GLORT_RAM_SKIP_DGLORT_DEC_LO = 35;
localparam GLORT_RAM_SKIP_DGLORT_DEC_HI = 35;
localparam GLORT_RAM_SKIP_DGLORT_DEC_RESET = 1'h0;
localparam GLORT_RAM_HASH_ROTATION_LO = 34;
localparam GLORT_RAM_HASH_ROTATION_HI = 34;
localparam GLORT_RAM_HASH_ROTATION_RESET = 1'h0;
localparam GLORT_RAM_DEST_COUNT_LO = 30;
localparam GLORT_RAM_DEST_COUNT_HI = 33;
localparam GLORT_RAM_DEST_COUNT_RESET = 4'h0;
localparam GLORT_RAM_RANGE_SUB_INDEX_B_LO = 22;
localparam GLORT_RAM_RANGE_SUB_INDEX_B_HI = 29;
localparam GLORT_RAM_RANGE_SUB_INDEX_B_RESET = 8'h0;
localparam GLORT_RAM_RANGE_SUB_INDEX_A_LO = 14;
localparam GLORT_RAM_RANGE_SUB_INDEX_A_HI = 21;
localparam GLORT_RAM_RANGE_SUB_INDEX_A_RESET = 8'h0;
localparam GLORT_RAM_DEST_INDEX_LO = 2;
localparam GLORT_RAM_DEST_INDEX_HI = 13;
localparam GLORT_RAM_DEST_INDEX_RESET = 12'h0;
localparam GLORT_RAM_STRICT_LO = 0;
localparam GLORT_RAM_STRICT_HI = 1;
localparam GLORT_RAM_STRICT_RESET = 2'h0;
localparam GLORT_RAM_USEMASK = 64'hFFFFFFFFF;
localparam GLORT_RAM_RO_MASK = 64'h0;
localparam GLORT_RAM_WO_MASK = 64'h0;
localparam GLORT_RAM_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [15:0] KEY_INVERT;  // RW
    logic [15:0] KEY;  // RW
} GLORT_CAM_t;

localparam GLORT_CAM_REG_STRIDE = 48'h8;
localparam GLORT_CAM_REG_ENTRIES = 64;
localparam GLORT_CAM_CR_ADDR = 48'hC0400;
localparam GLORT_CAM_SIZE = 64;
localparam GLORT_CAM_KEY_INVERT_LO = 16;
localparam GLORT_CAM_KEY_INVERT_HI = 31;
localparam GLORT_CAM_KEY_INVERT_RESET = 16'hffff;
localparam GLORT_CAM_KEY_LO = 0;
localparam GLORT_CAM_KEY_HI = 15;
localparam GLORT_CAM_KEY_RESET = 16'hffff;
localparam GLORT_CAM_USEMASK = 64'hFFFFFFFF;
localparam GLORT_CAM_RO_MASK = 64'h0;
localparam GLORT_CAM_WO_MASK = 64'h0;
localparam GLORT_CAM_RESET = 64'hFFFFFFFF;

typedef struct packed {
    logic [63:0] USED;  // RW/1C/V
} CGRP_USED_TABLE_t;

localparam CGRP_USED_TABLE_REG_STRIDE = 48'h8;
localparam CGRP_USED_TABLE_REG_ENTRIES = 65;
localparam CGRP_USED_TABLE_CR_ADDR = 48'hC0760;
localparam CGRP_USED_TABLE_SIZE = 64;
localparam CGRP_USED_TABLE_USED_LO = 0;
localparam CGRP_USED_TABLE_USED_HI = 63;
localparam CGRP_USED_TABLE_USED_RESET = 64'h0;
localparam CGRP_USED_TABLE_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam CGRP_USED_TABLE_RO_MASK = 64'h0;
localparam CGRP_USED_TABLE_WO_MASK = 64'h0;
localparam CGRP_USED_TABLE_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_EGRESS_VID_TABLE_t;

typedef logic [7:0] we_EGRESS_VID_CFG_t;

typedef logic [7:0] we_INGRESS_MST_TABLE_t;

typedef logic [7:0] we_EGRESS_MST_TABLE_t;

typedef logic [7:0] we_GLORT_DIRECT_MAP_CTRL_t;

typedef logic [7:0] we_GLORT_DIRECT_MAP_DST0_t;

typedef logic [7:0] we_GLORT_DIRECT_MAP_DST1_t;

typedef logic [7:0] we_GLORT_DIRECT_MAP_DST2_t;

typedef logic [7:0] we_GLORT_DIRECT_MAP_DST3_t;

typedef logic [7:0] we_GLORT_DIRECT_MAP_DST4_t;

typedef logic [7:0] we_GLORT_RAM_t;

typedef logic [7:0] we_GLORT_CAM_t;

typedef logic [7:0] we_CGRP_USED_TABLE_t;

typedef struct packed {
    we_EGRESS_VID_TABLE_t EGRESS_VID_TABLE;
    we_EGRESS_VID_CFG_t EGRESS_VID_CFG;
    we_INGRESS_MST_TABLE_t INGRESS_MST_TABLE;
    we_EGRESS_MST_TABLE_t EGRESS_MST_TABLE;
    we_GLORT_DIRECT_MAP_CTRL_t GLORT_DIRECT_MAP_CTRL;
    we_GLORT_DIRECT_MAP_DST0_t GLORT_DIRECT_MAP_DST0;
    we_GLORT_DIRECT_MAP_DST1_t GLORT_DIRECT_MAP_DST1;
    we_GLORT_DIRECT_MAP_DST2_t GLORT_DIRECT_MAP_DST2;
    we_GLORT_DIRECT_MAP_DST3_t GLORT_DIRECT_MAP_DST3;
    we_GLORT_DIRECT_MAP_DST4_t GLORT_DIRECT_MAP_DST4;
    we_GLORT_RAM_t GLORT_RAM;
    we_GLORT_CAM_t GLORT_CAM;
    we_CGRP_USED_TABLE_t CGRP_USED_TABLE;
} mby_ppe_mst_glort_map_handcoded_t;

typedef logic [7:0] re_EGRESS_VID_TABLE_t;

typedef logic [7:0] re_EGRESS_VID_CFG_t;

typedef logic [7:0] re_INGRESS_MST_TABLE_t;

typedef logic [7:0] re_EGRESS_MST_TABLE_t;

typedef logic [7:0] re_GLORT_DIRECT_MAP_CTRL_t;

typedef logic [7:0] re_GLORT_DIRECT_MAP_DST0_t;

typedef logic [7:0] re_GLORT_DIRECT_MAP_DST1_t;

typedef logic [7:0] re_GLORT_DIRECT_MAP_DST2_t;

typedef logic [7:0] re_GLORT_DIRECT_MAP_DST3_t;

typedef logic [7:0] re_GLORT_DIRECT_MAP_DST4_t;

typedef logic [7:0] re_GLORT_RAM_t;

typedef logic [7:0] re_GLORT_CAM_t;

typedef logic [7:0] re_CGRP_USED_TABLE_t;

typedef struct packed {
    re_EGRESS_VID_TABLE_t EGRESS_VID_TABLE;
    re_EGRESS_VID_CFG_t EGRESS_VID_CFG;
    re_INGRESS_MST_TABLE_t INGRESS_MST_TABLE;
    re_EGRESS_MST_TABLE_t EGRESS_MST_TABLE;
    re_GLORT_DIRECT_MAP_CTRL_t GLORT_DIRECT_MAP_CTRL;
    re_GLORT_DIRECT_MAP_DST0_t GLORT_DIRECT_MAP_DST0;
    re_GLORT_DIRECT_MAP_DST1_t GLORT_DIRECT_MAP_DST1;
    re_GLORT_DIRECT_MAP_DST2_t GLORT_DIRECT_MAP_DST2;
    re_GLORT_DIRECT_MAP_DST3_t GLORT_DIRECT_MAP_DST3;
    re_GLORT_DIRECT_MAP_DST4_t GLORT_DIRECT_MAP_DST4;
    re_GLORT_RAM_t GLORT_RAM;
    re_GLORT_CAM_t GLORT_CAM;
    re_CGRP_USED_TABLE_t CGRP_USED_TABLE;
} mby_ppe_mst_glort_map_hc_re_t;

typedef logic handcode_rvalid_EGRESS_VID_TABLE_t;

typedef logic handcode_rvalid_EGRESS_VID_CFG_t;

typedef logic handcode_rvalid_INGRESS_MST_TABLE_t;

typedef logic handcode_rvalid_EGRESS_MST_TABLE_t;

typedef logic handcode_rvalid_GLORT_DIRECT_MAP_CTRL_t;

typedef logic handcode_rvalid_GLORT_DIRECT_MAP_DST0_t;

typedef logic handcode_rvalid_GLORT_DIRECT_MAP_DST1_t;

typedef logic handcode_rvalid_GLORT_DIRECT_MAP_DST2_t;

typedef logic handcode_rvalid_GLORT_DIRECT_MAP_DST3_t;

typedef logic handcode_rvalid_GLORT_DIRECT_MAP_DST4_t;

typedef logic handcode_rvalid_GLORT_RAM_t;

typedef logic handcode_rvalid_GLORT_CAM_t;

typedef logic handcode_rvalid_CGRP_USED_TABLE_t;

typedef struct packed {
    handcode_rvalid_EGRESS_VID_TABLE_t EGRESS_VID_TABLE;
    handcode_rvalid_EGRESS_VID_CFG_t EGRESS_VID_CFG;
    handcode_rvalid_INGRESS_MST_TABLE_t INGRESS_MST_TABLE;
    handcode_rvalid_EGRESS_MST_TABLE_t EGRESS_MST_TABLE;
    handcode_rvalid_GLORT_DIRECT_MAP_CTRL_t GLORT_DIRECT_MAP_CTRL;
    handcode_rvalid_GLORT_DIRECT_MAP_DST0_t GLORT_DIRECT_MAP_DST0;
    handcode_rvalid_GLORT_DIRECT_MAP_DST1_t GLORT_DIRECT_MAP_DST1;
    handcode_rvalid_GLORT_DIRECT_MAP_DST2_t GLORT_DIRECT_MAP_DST2;
    handcode_rvalid_GLORT_DIRECT_MAP_DST3_t GLORT_DIRECT_MAP_DST3;
    handcode_rvalid_GLORT_DIRECT_MAP_DST4_t GLORT_DIRECT_MAP_DST4;
    handcode_rvalid_GLORT_RAM_t GLORT_RAM;
    handcode_rvalid_GLORT_CAM_t GLORT_CAM;
    handcode_rvalid_CGRP_USED_TABLE_t CGRP_USED_TABLE;
} mby_ppe_mst_glort_map_hc_rvalid_t;

typedef logic handcode_wvalid_EGRESS_VID_TABLE_t;

typedef logic handcode_wvalid_EGRESS_VID_CFG_t;

typedef logic handcode_wvalid_INGRESS_MST_TABLE_t;

typedef logic handcode_wvalid_EGRESS_MST_TABLE_t;

typedef logic handcode_wvalid_GLORT_DIRECT_MAP_CTRL_t;

typedef logic handcode_wvalid_GLORT_DIRECT_MAP_DST0_t;

typedef logic handcode_wvalid_GLORT_DIRECT_MAP_DST1_t;

typedef logic handcode_wvalid_GLORT_DIRECT_MAP_DST2_t;

typedef logic handcode_wvalid_GLORT_DIRECT_MAP_DST3_t;

typedef logic handcode_wvalid_GLORT_DIRECT_MAP_DST4_t;

typedef logic handcode_wvalid_GLORT_RAM_t;

typedef logic handcode_wvalid_GLORT_CAM_t;

typedef logic handcode_wvalid_CGRP_USED_TABLE_t;

typedef struct packed {
    handcode_wvalid_EGRESS_VID_TABLE_t EGRESS_VID_TABLE;
    handcode_wvalid_EGRESS_VID_CFG_t EGRESS_VID_CFG;
    handcode_wvalid_INGRESS_MST_TABLE_t INGRESS_MST_TABLE;
    handcode_wvalid_EGRESS_MST_TABLE_t EGRESS_MST_TABLE;
    handcode_wvalid_GLORT_DIRECT_MAP_CTRL_t GLORT_DIRECT_MAP_CTRL;
    handcode_wvalid_GLORT_DIRECT_MAP_DST0_t GLORT_DIRECT_MAP_DST0;
    handcode_wvalid_GLORT_DIRECT_MAP_DST1_t GLORT_DIRECT_MAP_DST1;
    handcode_wvalid_GLORT_DIRECT_MAP_DST2_t GLORT_DIRECT_MAP_DST2;
    handcode_wvalid_GLORT_DIRECT_MAP_DST3_t GLORT_DIRECT_MAP_DST3;
    handcode_wvalid_GLORT_DIRECT_MAP_DST4_t GLORT_DIRECT_MAP_DST4;
    handcode_wvalid_GLORT_RAM_t GLORT_RAM;
    handcode_wvalid_GLORT_CAM_t GLORT_CAM;
    handcode_wvalid_CGRP_USED_TABLE_t CGRP_USED_TABLE;
} mby_ppe_mst_glort_map_hc_wvalid_t;

typedef logic handcode_error_EGRESS_VID_TABLE_t;

typedef logic handcode_error_EGRESS_VID_CFG_t;

typedef logic handcode_error_INGRESS_MST_TABLE_t;

typedef logic handcode_error_EGRESS_MST_TABLE_t;

typedef logic handcode_error_GLORT_DIRECT_MAP_CTRL_t;

typedef logic handcode_error_GLORT_DIRECT_MAP_DST0_t;

typedef logic handcode_error_GLORT_DIRECT_MAP_DST1_t;

typedef logic handcode_error_GLORT_DIRECT_MAP_DST2_t;

typedef logic handcode_error_GLORT_DIRECT_MAP_DST3_t;

typedef logic handcode_error_GLORT_DIRECT_MAP_DST4_t;

typedef logic handcode_error_GLORT_RAM_t;

typedef logic handcode_error_GLORT_CAM_t;

typedef logic handcode_error_CGRP_USED_TABLE_t;

typedef struct packed {
    handcode_error_EGRESS_VID_TABLE_t EGRESS_VID_TABLE;
    handcode_error_EGRESS_VID_CFG_t EGRESS_VID_CFG;
    handcode_error_INGRESS_MST_TABLE_t INGRESS_MST_TABLE;
    handcode_error_EGRESS_MST_TABLE_t EGRESS_MST_TABLE;
    handcode_error_GLORT_DIRECT_MAP_CTRL_t GLORT_DIRECT_MAP_CTRL;
    handcode_error_GLORT_DIRECT_MAP_DST0_t GLORT_DIRECT_MAP_DST0;
    handcode_error_GLORT_DIRECT_MAP_DST1_t GLORT_DIRECT_MAP_DST1;
    handcode_error_GLORT_DIRECT_MAP_DST2_t GLORT_DIRECT_MAP_DST2;
    handcode_error_GLORT_DIRECT_MAP_DST3_t GLORT_DIRECT_MAP_DST3;
    handcode_error_GLORT_DIRECT_MAP_DST4_t GLORT_DIRECT_MAP_DST4;
    handcode_error_GLORT_RAM_t GLORT_RAM;
    handcode_error_GLORT_CAM_t GLORT_CAM;
    handcode_error_CGRP_USED_TABLE_t CGRP_USED_TABLE;
} mby_ppe_mst_glort_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    EGRESS_VID_TABLE_t EGRESS_VID_TABLE;
    EGRESS_VID_CFG_t EGRESS_VID_CFG;
    INGRESS_MST_TABLE_t INGRESS_MST_TABLE;
    EGRESS_MST_TABLE_t EGRESS_MST_TABLE;
    GLORT_DIRECT_MAP_CTRL_t GLORT_DIRECT_MAP_CTRL;
    GLORT_DIRECT_MAP_DST0_t GLORT_DIRECT_MAP_DST0;
    GLORT_DIRECT_MAP_DST1_t GLORT_DIRECT_MAP_DST1;
    GLORT_DIRECT_MAP_DST2_t GLORT_DIRECT_MAP_DST2;
    GLORT_DIRECT_MAP_DST3_t GLORT_DIRECT_MAP_DST3;
    GLORT_DIRECT_MAP_DST4_t GLORT_DIRECT_MAP_DST4;
    GLORT_RAM_t GLORT_RAM;
    GLORT_CAM_t GLORT_CAM;
    CGRP_USED_TABLE_t CGRP_USED_TABLE;
} mby_ppe_mst_glort_map_hc_reg_read_t;

typedef struct packed {
    EGRESS_VID_TABLE_t EGRESS_VID_TABLE;
    EGRESS_VID_CFG_t EGRESS_VID_CFG;
    INGRESS_MST_TABLE_t INGRESS_MST_TABLE;
    EGRESS_MST_TABLE_t EGRESS_MST_TABLE;
    GLORT_DIRECT_MAP_CTRL_t GLORT_DIRECT_MAP_CTRL;
    GLORT_DIRECT_MAP_DST0_t GLORT_DIRECT_MAP_DST0;
    GLORT_DIRECT_MAP_DST1_t GLORT_DIRECT_MAP_DST1;
    GLORT_DIRECT_MAP_DST2_t GLORT_DIRECT_MAP_DST2;
    GLORT_DIRECT_MAP_DST3_t GLORT_DIRECT_MAP_DST3;
    GLORT_DIRECT_MAP_DST4_t GLORT_DIRECT_MAP_DST4;
    GLORT_RAM_t GLORT_RAM;
    GLORT_CAM_t GLORT_CAM;
    CGRP_USED_TABLE_t CGRP_USED_TABLE;
} mby_ppe_mst_glort_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_mst_glort_map_pkg

`endif // MBY_PPE_MST_GLORT_MAP_PKG_VH
