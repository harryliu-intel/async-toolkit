//                                                                             
// File:       MBY_ral_env.svh                                                 
// Creator:    kmoses1                                                         
// Time:       Sunday Feb 2, 2014 [8:21:51 am]                                 
//                                                                             
// Path:       /tmp/kmoses1/nebulon_run/20231                                  
// Arguments:  /p/com/eda/denali/blueprint/3.7.4/Linux/blueprint -fuse -html -I
//             /p/com/eda/intel/nebulon/2.07p2/include/ -ovm                   
//             mby_fusegen_nebulon.rdl                                         
//                                                                             
// Sources:    /nfs/iil/proj/mpg/kmoses1_wa1/ip_template-nhdk-x0_new/source/rdl/mby_fusegen_nebulon.rdl:5b3e806ef7d09a39437507f3cfbd0ecb
//             /p/com/eda/intel/nebulon/2.07p2/generators/generator_common.pm:4973c402c43f97e18c4aba02585df570
//             /p/com/eda/intel/nebulon/2.07p2/generators/html.pm:a408055bdb3ba8a9656d793e9472104f
//             /p/com/eda/intel/nebulon/2.07p2/generators/ovm.pm:e21c7be001887ff41e17c43b43b1fcdc
//             /p/com/eda/intel/nebulon/2.07p2/include/fuse_udp.rdl:c11891ce81c95bc748bf1f2bdbde2f6f
//             /usr/intel/pkgs/perl/5.8.7/lib64/5.8.7/Digest/base.pm:54bebd0439900c1d44d212cba39747b5
//             /usr/intel/pkgs/perl/5.8.7/lib64/site_perl/Devel/StackTrace.pm:3b99e973435e2dea00aa3a8d6f1b9ddd
//                                                                             
// Blueprint:   3.7.4 (Tue Jun 23 00:17:01 PDT 2009)                           
// Machine:    icsl0104                                                        
// OS:         Linux 2.6.16.60-0.58.1.3835.0.PTF.638363-smp                    
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2014 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY DENALI BLUEPRINT, DO NOT EDIT       
//                                                                             


//RAL code compatible with Saola versions: v20131113 and newer 

`ifndef SLA_PATH_TO_STRING
`define SLA_PATH_TO_STRING(SIG_PATH) `"SIG_PATH`"
`endif

`include "mby_fuse_regs.svh"


class MBY_ral_env extends sla_ral_env;

  `ovm_component_utils(MBY_ral_env);

  rand mby_fuse_file mby_fuse;

  // --------------------------
  function new( string n="MBY_ral_env", ovm_component p = null, string hdl_path = "");
    super.new( n, p, hdl_path);
  endfunction : new


  // --------------------------
  virtual function void build();
    super.build();

    mby_fuse = mby_fuse_file::type_id::create("mby_fuse", this);
    add_file("mby_fuse",mby_fuse);

  endfunction : build

  // --------------------------
  function void connect();
    mby_fuse.set_base(4'h0);


    set_bit_blasting(1);
  endfunction : connect


  virtual function string sprint_sv_ral_env();  
     return({"Generated SV RAL Env ---> ", `__FILE__}); 
  endfunction  
endclass : MBY_ral_env
