// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

//-----------------------------------------------------
// DUT IF signal connection
//-----------------------------------------------------
//assign `DUT_IF.XTAL_IN      = `HVL_TOP.xtal_25M_clk.clk;

//------------------------------------------------------
// FCSIG IF signal connection
//------------------------------------------------------
