magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -8 58 -4 59
rect -8 52 -4 56
rect -8 49 -4 50
<< pdiffusion >>
rect 8 61 12 62
rect 8 58 12 59
rect 8 52 12 54
rect 8 49 12 50
<< ntransistor >>
rect -8 56 -4 58
rect -8 50 -4 52
<< ptransistor >>
rect 8 59 12 61
rect 8 50 12 52
<< polysilicon >>
rect 4 59 8 61
rect 12 59 15 61
rect 4 58 6 59
rect -11 56 -8 58
rect -4 56 6 58
rect -11 50 -8 52
rect -4 50 -1 52
rect 5 50 8 52
rect 12 50 15 52
<< ndcontact >>
rect -8 59 -4 63
rect -8 45 -4 49
<< pdcontact >>
rect 8 62 12 66
rect 8 54 12 58
rect 8 45 12 49
<< metal1 >>
rect -8 59 -4 63
rect 8 62 12 66
rect -7 57 -4 59
rect 8 57 12 58
rect -7 54 12 57
rect -8 45 -4 49
rect 8 45 12 49
<< labels >>
rlabel polysilicon -9 51 -9 51 3 _SReset!
rlabel polysilicon -9 57 -9 57 3 a
rlabel polysilicon 13 51 13 51 1 _PReset!
rlabel space -11 45 -8 63 7 ^n
rlabel polysilicon 13 60 13 60 7 a
rlabel space 12 56 15 66 3 ^p
rlabel pdcontact 10 47 10 47 5 Vdd!
rlabel ndcontact -6 61 -6 61 4 x
rlabel ndcontact -6 47 -6 47 5 GND!
rlabel pdcontact 10 64 10 64 5 Vdd!
rlabel pdcontact 10 56 10 56 7 x
<< end >>
