*
* TEST SPICE INPUT FILE FOR
* Subnet test environment generation
* Test of sneak paths between subnet driver networks.
*
*
.SUBCKT TESTCELL a b c d
MXa2s_dout[20]/M+68     GND!    Xa2s_dout[20]/_r:1      
+	Xa2s_dout[20]/58        GND! nmos_2v L=0.18U W=2.4U AD=1.296P
+	 AS=0.36P PD=3.48U PS=0.3U
MXa2s_dout[20]/M+69     odq[20]:1       Xa2s_dout[20]/_R.1:2    
+	Xa2s_dout[20]/58        GND! nmos_2v L=0.18U W=2.4U AD=0.72P
+	 AS=0.36P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+70     Xa2s_dout[20]/57        Xa2s_dout[20]/_r:4
+	odq[20]:1       GND! nmos_2v L=0.18U W=2.4U AD=0.36P AS=0.72P
+	 PD=0.3U PS=0.6U
MXa2s_dout[20]/M+79     Xa2s_dout[20]/Rv:13     Xa2s_dout[20]/_R.1:14
+	Xa2s_dout[20]/72        GND! nmos_2v L=0.18U W=0.96U AD=0.432P
+	 AS=0.144P PD=2.04U PS=0.3U
MXa2s_dout[20]/M+80     Xa2s_dout[20]/72        Xa2s_dout[20]/_R.0:3
+	GND!    GND! nmos_2v L=0.18U W=0.96U AD=0.144P AS=0.518P
+	 PD=0.3U PS=2.04U
MXa2s_dout[20]/M+71     Xa2s_dout[20]/57        Xa2s_dout[20]/_R.1:5
+	GND!    GND! nmos_2v L=0.18U W=2.4U AD=0.36P AS=0.72P PD=0.3U
+	 PS=0.6U
MXa2s_dout[20]/M+64     GND!    Xa2s_dout[20]/_r:10     
+	Xa2s_dout[20]/61        GND! nmos_2v L=0.18U W=2.4U AD=0.72P
+	 AS=0.36P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+65     Xa2s_dout[20]/61        Xa2s_dout[20]/_R.1:8
+	odq[20]:16      GND! nmos_2v L=0.18U W=2.4U AD=0.36P AS=0.72P
+	 PD=0.3U PS=0.6U
MXa2s_dout[20]/M+66     odq[20]:16      Xa2s_dout[20]/_r:7      
+	Xa2s_dout[20]/60        GND! nmos_2v L=0.18U W=2.4U AD=0.72P
+	 AS=0.36P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+67     Xa2s_dout[20]/60        Xa2s_dout[20]/_R.1:11
+	GND!    GND! nmos_2v L=0.18U W=2.4U AD=0.36P AS=1.296P PD=0.3U
+	 PS=3.48U
MXa2s_dout[20]/M+74     Xa2s_dout[20]/_r:16     _SReset!:5205   
+	Xa2s_dout[20]/55        GND! nmos_2v L=0.18U W=4.56U AD=2.462P
+	 AS=0.684P PD=5.64U PS=0.3U
MXa2s_dout[20]/M+75     Xa2s_dout[20]/54        odq[20]:17      
+	Xa2s_dout[20]/55        GND! nmos_2v L=0.18U W=4.56U AD=0.684P
+	 AS=0.684P PD=0.3U PS=0.3U
MXa2s_dout[20]/M+76     Xa2s_dout[20]/54        Xa2s_dout[20]/_R.0:22
+	GND!    GND! nmos_2v L=0.18U W=4.56U AD=0.684P AS=2.462P
+	 PD=0.3U PS=5.64U
MXa2s_dout[20]/M+59     Xa2s_dout[20]/__Le:10   Xa2s_dout[20]/7:6
+	GND!    GND! nmos_2v L=0.48U W=0.24U AD=0.274P AS=0.274P
+	 PD=2.04U PS=2.04U
MXa2s_dout[20]/M+60     Xa2s_dout[20]/_noR:7    Xa2s_dout[20]/6:6
+	GND!    GND! nmos_2v L=0.42U W=0.24U AD=0.302P AS=0.274P
+	 PD=2.28U PS=2.04U
MXa2s_dout[20]/M+77     Xa2s_dout[20]/7:4       Xa2s_dout[20]/__Le:1
+	GND!    GND! nmos_2v L=0.18U W=0.48U AD=0.259P AS=0.259P
+	 PD=1.56U PS=1.56U
MXa2s_dout[20]/M+72     Xa2s_dout[20]/_Le:1     Xa2s_dout[20]/__Le:6
+	Xa2s_dout[20]/56        GND! nmos_2v L=0.18U W=2.82U AD=1.523P
+	 AS=0.423P PD=3.9U PS=0.3U
MXa2s_dout[20]/M+73     GND!    _SReset!:5066   Xa2s_dout[20]/56
+	GND! nmos_2v L=0.18U W=2.82U AD=1.523P AS=0.423P PD=3.9U
+	 PS=0.3U
MXa2s_dout[20]/M+78     GND!    Xa2s_dout[20]/_noR:3    
+	Xa2s_dout[20]/6:4       GND! nmos_2v L=0.18U W=0.48U AD=0.259P
+	 AS=0.259P PD=1.56U PS=1.56U
MXa2s_dout[20]/M+61     Xa2s_dout[20]/71        Xa2s_dout[20]/_noR:11
+	Xa2s_dout[20]/Rc:1      GND! nmos_2v L=0.18U W=1.86U AD=0.279P
+	 AS=1.004P PD=0.3U PS=2.94U
MXa2s_dout[20]/M+62     Xa2s_dout[20]/62        Xa2s_dout[20]/_R.0:19
+	Xa2s_dout[20]/71        GND! nmos_2v L=0.18U W=1.86U AD=0.279P
+	 AS=0.279P PD=0.3U PS=0.3U
MXa2s_dout[20]/M+63     GND!    Xa2s_dout[20]/_R.1:16   
+	Xa2s_dout[20]/62        GND! nmos_2v L=0.18U W=1.86U AD=1.004P
+	 AS=0.279P PD=2.94U PS=0.3U
MXa2s_dout[20]/M+54     Xa2s_dout[20]/53        clk:4342        
+	Xa2s_dout[20]/51:2      GND! nmos_2v L=0.18U W=1.2U AD=0.18P
+	 AS=0.518P PD=0.3U PS=2.28U
MXa2s_dout[20]/M+55     Xa2s_dout[20]/__Le:11   Xa2s_dout[20]/clk0:11
+	Xa2s_dout[20]/53        GND! nmos_2v L=0.18U W=1.2U AD=0.36P
+	 AS=0.18P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+56     Xa2s_dout[20]/__Le:11   Xa2s_dout[20]/_clk0:11
+	Xa2s_dout[20]/52        GND! nmos_2v L=0.18U W=1.2U AD=0.36P
+	 AS=0.18P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+57     Xa2s_dout[20]/52        Xa2s_dout[20]/_clk:7
+	Xa2s_dout[20]/51:1      GND! nmos_2v L=0.18U W=1.2U AD=0.18P
+	 AS=0.36P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+58     Xa2s_dout[20]/51:1      Xa2s_dout[20]/Rv:3
+	GND!    GND! nmos_2v L=0.18U W=1.2U AD=0.36P AS=0.648P PD=0.6U
+	 PS=2.28U
MXa2s_dout[20]/M+29     GND!    Xa2s_dout[20]/8:6       
+	Xa2s_dout[20]/_R.1:41   GND! nmos_2v L=0.48U W=0.24U AD=0.274P
+	 AS=0.274P PD=2.04U PS=2.04U
MXa2s_dout[20]/M+30     Xa2s_dout[20]/Rv:9      Xa2s_dout[20]/9:6
+	GND!    GND! nmos_2v L=0.54U W=0.24U AD=0.288P AS=0.259P
+	 PD=2.16U PS=1.92U
MXa2s_dout[20]/M+31     GND!    Xa2s_dout[20]/Rv:5      
+	Xa2s_dout[20]/9:4       GND! nmos_2v L=0.18U W=0.48U AD=0.259P
+	 AS=0.259P PD=1.56U PS=1.56U
MXa2s_dout[20]/M+32     GND!    Xa2s_dout[20]/_R.1:36   
+	Xa2s_dout[20]/8:4       GND! nmos_2v L=0.18U W=0.48U AD=0.259P
+	 AS=0.259P PD=1.56U PS=1.56U
MXa2s_dout[20]/M+37     dout[22].e:4    Xa2s_dout[20]/_Le:9     GND!
+	GND! nmos_2v L=0.18U W=2.7U AD=0.81P AS=1.458P PD=0.6U
+	 PS=3.78U
MXa2s_dout[20]/M+36     GND!    Xa2s_dout[20]/_Le:17    dout[22].e:4
+	GND! nmos_2v L=0.18U W=2.7U AD=0.81P AS=0.81P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+35     dout[22].e:3    Xa2s_dout[20]/_Le:19    GND!
+	GND! nmos_2v L=0.18U W=2.7U AD=0.81P AS=0.81P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+34     GND!    Xa2s_dout[20]/_Le:20    dout[22].e:3
+	GND! nmos_2v L=0.18U W=2.7U AD=1.458P AS=0.81P PD=3.78U
+	 PS=0.6U
MXa2s_dout[20]/M+33     GND!    _PReset!:6731   Xa2s_dout[20]/PReset:9
+	GND! nmos_2v L=0.18U W=1.2U AD=0.648P AS=0.648P PD=2.28U
+	 PS=2.28U
MXa2s_dout[20]/M+38     Xa2s_dout[20]/33        Xa2s_dout[20]/_clk:18
+	Xa2s_dout[20]/31:2      GND! nmos_2v L=0.18U W=1.44U AD=0.216P
+	 AS=0.605P PD=0.3U PS=2.52U
MXa2s_dout[20]/M+39     GND!    Xa2s_dout[20]/clk0:16   
+	Xa2s_dout[20]/33        GND! nmos_2v L=0.18U W=1.44U AD=0.778P
+	 AS=0.216P PD=2.52U PS=0.3U
MXa2s_dout[20]/M+40     Xa2s_dout[20]/29:1      Xa2s_dout[20]/_grant:4
+	GND!    GND! nmos_2v L=0.18U W=1.44U AD=0.605P AS=0.432P
+	 PD=2.52U PS=0.6U
MXa2s_dout[20]/M+41     GND!    Xa2s_dout[20]/_clk0:13  
+	Xa2s_dout[20]/32        GND! nmos_2v L=0.18U W=1.44U AD=0.432P
+	 AS=0.216P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+42     Xa2s_dout[20]/32        clk:4275        
+	Xa2s_dout[20]/31:1      GND! nmos_2v L=0.18U W=1.44U AD=0.216P
+	 AS=0.432P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+43     Xa2s_dout[20]/_noR:27   Xa2s_dout[20]/_grant:5
+	Xa2s_dout[20]/31:1      GND! nmos_2v L=0.18U W=1.44U AD=0.432P
+	 AS=0.432P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+44     Xa2s_dout[20]/30        Xa2s_dout[20]/clk0:14
+	Xa2s_dout[20]/_noR:27   GND! nmos_2v L=0.18U W=1.44U AD=0.216P
+	 AS=0.432P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+45     Xa2s_dout[20]/30        Xa2s_dout[20]/_clk:17
+	Xa2s_dout[20]/29:2      GND! nmos_2v L=0.18U W=1.44U AD=0.216P
+	 AS=0.432P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+46     Xa2s_dout[20]/29:2      clk:4340        
+	Xa2s_dout[20]/28        GND! nmos_2v L=0.18U W=1.44U AD=0.432P
+	 AS=0.216P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+47     Xa2s_dout[20]/28        Xa2s_dout[20]/_clk0:16
+	Xa2s_dout[20]/_noR:29   GND! nmos_2v L=0.18U W=1.44U AD=0.216P
+	 AS=0.605P PD=0.3U PS=2.52U
MXa2s_dout[20]/M+48     Xa2s_dout[20]/26:2      clk:4343        
+	Xa2s_dout[20]/_clk0:18  GND! nmos_2v L=0.18U W=1.92U AD=0.864P
+	 AS=0.864P PD=3U PS=3U
MXa2s_dout[20]/M+49     Xa2s_dout[20]/27:1      Xa2s_dout[20]/Rc:12
+	Xa2s_dout[20]/_clk0:24  GND! nmos_2v L=0.18U W=1.92U AD=0.864P
+	 AS=0.576P PD=3U PS=0.6U
MXa2s_dout[20]/M+50     Xa2s_dout[20]/27:2      Xa2s_dout[20]/PReset:6
+	Xa2s_dout[20]/_clk0:24  GND! nmos_2v L=0.18U W=1.92U AD=0.576P
+	 AS=0.576P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+51     GND!    clk:4492        Xa2s_dout[20]/27:2
+	GND! nmos_2v L=0.18U W=1.92U AD=0.576P AS=0.576P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+52     GND!    Xa2s_dout[20]/PReset:8  
+	Xa2s_dout[20]/26:1      GND! nmos_2v L=0.18U W=1.92U AD=0.576P
+	 AS=0.576P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+53     Xa2s_dout[20]/26:1      Xa2s_dout[20]/Rc:8
+	GND!    GND! nmos_2v L=0.18U W=1.92U AD=0.576P AS=1.037P
+	 PD=0.6U PS=3U
MXa2s_dout[20]/M+28     Xa2s_dout[20]/15:5      oe:420  GND!    GND!
+	 nmos_2v L=0.18U W=4.08U AD=1.224P AS=2.203P PD=0.6U PS=5.16U
MXa2s_dout[20]/M+18     Xa2s_dout[20]/20        Xa2s_dout[20]/_clk0:41
+	Xa2s_dout[20]/15:5      GND! nmos_2v L=0.18U W=4.08U AD=0.612P
+	 AS=1.224P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+19     Xa2s_dout[20]/17:1      clk:4908        
+	Xa2s_dout[20]/20        GND! nmos_2v L=0.18U W=4.08U AD=1.224P
+	 AS=0.612P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+21     Xa2s_dout[20]/_R.1:46   dout[22].1:6    
+	Xa2s_dout[20]/17:1      GND! nmos_2v L=0.18U W=4.08U AD=1.224P
+	 AS=1.224P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+20     Xa2s_dout[20]/17:5      dout[22].1:7    
+	Xa2s_dout[20]/_R.1:46   GND! nmos_2v L=0.18U W=4.08U AD=1.224P
+	 AS=1.224P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+22     Xa2s_dout[20]/19        Xa2s_dout[20]/_clk:30
+	Xa2s_dout[20]/17:5      GND! nmos_2v L=0.18U W=4.08U AD=0.612P
+	 AS=1.224P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+23     Xa2s_dout[20]/15:7      Xa2s_dout[20]/clk0:28
+	Xa2s_dout[20]/19        GND! nmos_2v L=0.18U W=4.08U AD=1.224P
+	 AS=0.612P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+24     Xa2s_dout[20]/18        clk:4909        
+	Xa2s_dout[20]/15:7      GND! nmos_2v L=0.18U W=4.08U AD=0.612P
+	 AS=1.224P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+25     Xa2s_dout[20]/17:3      Xa2s_dout[20]/_clk0:40
+	Xa2s_dout[20]/18        GND! nmos_2v L=0.18U W=4.08U AD=1.224P
+	 AS=0.612P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+8      Xa2s_dout[20]/_R.0:29   dout[22].0:5    
+	Xa2s_dout[20]/21:1      GND! nmos_2v L=0.18U W=3U AD=0.9P
+	 AS=1.447P PD=0.6U PS=4.08U
MXa2s_dout[20]/M+7      Xa2s_dout[20]/21:2      dout[22].0:3    
+	Xa2s_dout[20]/_R.0:29   GND! nmos_2v L=0.18U W=3U AD=0.9P
+	 AS=0.9P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+9      Xa2s_dout[20]/25        Xa2s_dout[20]/_clk:27
+	Xa2s_dout[20]/21:2      GND! nmos_2v L=0.18U W=3U AD=0.45P
+	 AS=0.9P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+10     Xa2s_dout[20]/15:10     Xa2s_dout[20]/clk0:32
+	Xa2s_dout[20]/25        GND! nmos_2v L=0.18U W=3U AD=0.9P
+	 AS=0.45P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+11     Xa2s_dout[20]/24        Xa2s_dout[20]/_clk:29
+	Xa2s_dout[20]/15:10     GND! nmos_2v L=0.18U W=3U AD=0.45P
+	 AS=0.9P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+26     Xa2s_dout[20]/16        Xa2s_dout[20]/clk0:29
+	Xa2s_dout[20]/17:3      GND! nmos_2v L=0.18U W=4.08U AD=0.612P
+	 AS=1.224P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+27     Xa2s_dout[20]/15:13     Xa2s_dout[20]/_clk:31
+	Xa2s_dout[20]/16        GND! nmos_2v L=0.18U W=4.08U AD=1.224P
+	 AS=0.612P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+17     GND!    oe:452  Xa2s_dout[20]/15:13     GND!
+	 nmos_2v L=0.18U W=4.08U AD=2.203P AS=1.224P PD=5.16U PS=0.6U
MXa2s_dout[20]/M+12     Xa2s_dout[20]/21:4      Xa2s_dout[20]/clk0:33
+	Xa2s_dout[20]/24        GND! nmos_2v L=0.18U W=3U AD=0.9P
+	 AS=0.45P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+0      GND!    Xa2s_dout[20]/clk0:25   
+	Xa2s_dout[20]/_clk0:60  GND! nmos_2v L=0.48U W=0.24U AD=0.288P
+	 AS=0.288P PD=2.16U PS=2.16U
MXa2s_dout[20]/M+1      Xa2s_dout[20]/_R.0:34   Xa2s_dout[20]/10:6
+	GND!    GND! nmos_2v L=0.48U W=0.24U AD=0.274P AS=0.274P
+	 PD=2.04U PS=2.04U
MXa2s_dout[20]/M+2      GND!    oe:175  Xa2s_dout[20]/_grant:7  GND!
+	 nmos_2v L=0.18U W=1.2U AD=0.648P AS=0.648P PD=2.28U PS=2.28U
MXa2s_dout[20]/M+5      Xa2s_dout[20]/_clk:32   clk:4974        GND!
+	GND! nmos_2v L=0.18U W=2.04U AD=1.102P AS=1.102P PD=3.12U
+	 PS=3.12U
MXa2s_dout[20]/M+4      GND!    Xa2s_dout[20]/_clk0:49  
+	Xa2s_dout[20]/clk0:23   GND! nmos_2v L=0.18U W=1.2U AD=0.648P
+	 AS=0.36P PD=2.28U PS=0.6U
MXa2s_dout[20]/M+3      Xa2s_dout[20]/clk0:23   Xa2s_dout[20]/_clk0:51
+	GND!    GND! nmos_2v L=0.18U W=1.2U AD=0.36P AS=0.648P PD=0.6U
+	 PS=2.28U
MXa2s_dout[20]/M+6      Xa2s_dout[20]/10:4      Xa2s_dout[20]/_R.0:30
+	GND!    GND! nmos_2v L=0.18U W=0.48U AD=0.259P AS=0.259P
+	 PD=1.56U PS=1.56U
MXa2s_dout[20]/M+13     Xa2s_dout[20]/23        Xa2s_dout[20]/_clk0:39
+	Xa2s_dout[20]/21:4      GND! nmos_2v L=0.18U W=3U AD=0.45P
+	 AS=0.9P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+14     Xa2s_dout[20]/15:12     clk:4844        
+	Xa2s_dout[20]/23        GND! nmos_2v L=0.18U W=3U AD=0.9P
+	 AS=0.45P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+15     Xa2s_dout[20]/22        Xa2s_dout[20]/_clk0:59
+	Xa2s_dout[20]/15:12     GND! nmos_2v L=0.18U W=3U AD=0.45P
+	 AS=0.9P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+16     Xa2s_dout[20]/21:6      clk:4845        
+	Xa2s_dout[20]/22        GND! nmos_2v L=0.18U W=3U AD=1.447P
+	 AS=0.45P PD=4.08U PS=0.3U
MXa2s_dout[20]/M+138    odq[20]:12      Xa2s_dout[20]/_r:2      Vdd!
+	Vdd! pmos_2v L=0.18U W=2.22U AD=0.666P AS=1.199P PD=0.6U
+	 PS=3.3U
MXa2s_dout[20]/M+139    Vdd!    Xa2s_dout[20]/_R.1:3    odq[20]:12
+	Vdd! pmos_2v L=0.18U W=2.22U AD=0.666P AS=0.666P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+136    odq[20]:1       Xa2s_dout[20]/_r:5      Vdd!
+	Vdd! pmos_2v L=0.18U W=2.22U AD=0.666P AS=0.666P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+137    Vdd!    Xa2s_dout[20]/_R.1:6    odq[20]:1
+	Vdd! pmos_2v L=0.18U W=2.22U AD=0.666P AS=0.666P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+134    odq[20]:16      Xa2s_dout[20]/_r:11     Vdd!
+	Vdd! pmos_2v L=0.18U W=2.22U AD=0.666P AS=0.666P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+135    Vdd!    Xa2s_dout[20]/_R.1:9    odq[20]:16
+	Vdd! pmos_2v L=0.18U W=2.22U AD=0.666P AS=0.666P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+132    odq[20]:11      Xa2s_dout[20]/_r:8      Vdd!
+	Vdd! pmos_2v L=0.18U W=2.22U AD=0.666P AS=0.666P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+133    Vdd!    Xa2s_dout[20]/_R.1:12   odq[20]:11
+	Vdd! pmos_2v L=0.18U W=2.22U AD=1.199P AS=0.666P PD=3.3U
+	 PS=0.6U
MXa2s_dout[20]/M+140    Vdd!    _SReset!:5206   Xa2s_dout[20]/_r:16
+	Vdd! pmos_2v L=0.18U W=3.06U AD=0.918P AS=1.652P PD=0.6U
+	 PS=4.14U
MXa2s_dout[20]/M+99     Vdd!    Xa2s_dout[20]/_r:20     
+	Xa2s_dout[20]/5 Vdd! pmos_2v L=0.18U W=1.2U AD=0.648P AS=0.18P
+	 PD=2.28U PS=0.3U
MXa2s_dout[20]/M+100    Xa2s_dout[20]/5 Xa2s_dout[20]/_R.1:31   
+	Xa2s_dout[20]/Rv:11     Vdd! pmos_2v L=0.18U W=1.2U AD=0.18P
+	 AS=0.36P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+101    Xa2s_dout[20]/Rv:11     Xa2s_dout[20]/_R.0:17
+	Xa2s_dout[20]/4 Vdd! pmos_2v L=0.18U W=1.2U AD=0.36P AS=0.18P
+	 PD=0.6U PS=0.3U
MXa2s_dout[20]/M+102    Vdd!    odq[20]:21      Xa2s_dout[20]/4 Vdd!
+	 pmos_2v L=0.18U W=1.2U AD=0.36P AS=0.18P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+103    Xa2s_dout[20]/3 Xa2s_dout[20]/_R.1:29   Vdd!
+	Vdd! pmos_2v L=0.18U W=1.2U AD=0.18P AS=0.36P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+104    Xa2s_dout[20]/3 Xa2s_dout[20]/_r:19     
+	Xa2s_dout[20]/Rv:14     Vdd! pmos_2v L=0.18U W=1.2U AD=0.18P
+	 AS=0.36P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+105    Xa2s_dout[20]/Rv:14     odq[20]:19      
+	Xa2s_dout[20]/2 Vdd! pmos_2v L=0.18U W=1.2U AD=0.36P AS=0.18P
+	 PD=0.6U PS=0.3U
MXa2s_dout[20]/M+106    Xa2s_dout[20]/2 Xa2s_dout[20]/_R.0:13   Vdd!
+	Vdd! pmos_2v L=0.18U W=1.2U AD=0.18P AS=0.648P PD=0.3U
+	 PS=2.28U
MXa2s_dout[20]/M+107    Xa2s_dout[20]/14        Xa2s_dout[20]/clk0:2
+	Vdd!    Vdd! pmos_2v L=0.18U W=2.16U AD=0.324P AS=1.166P
+	 PD=0.3U PS=3.24U
MXa2s_dout[20]/M+108    Xa2s_dout[20]/14        clk:3718        
+	Xa2s_dout[20]/_noR:21   Vdd! pmos_2v L=0.18U W=2.16U AD=0.324P
+	 AS=0.648P PD=0.3U PS=0.6U
MXa2s_dout[20]/M+109    Xa2s_dout[20]/_noR:21   Xa2s_dout[20]/_clk:5
+	Xa2s_dout[20]/13        Vdd! pmos_2v L=0.18U W=2.16U AD=0.648P
+	 AS=0.324P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+110    Xa2s_dout[20]/13        Xa2s_dout[20]/_clk0:9
+	Vdd!    Vdd! pmos_2v L=0.18U W=2.16U AD=0.324P AS=0.648P
+	 PD=0.3U PS=0.6U
MXa2s_dout[20]/M+111    Vdd!    Xa2s_dout[20]/_clk:3    
+	Xa2s_dout[20]/12        Vdd! pmos_2v L=0.18U W=2.16U AD=0.648P
+	 AS=0.324P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+112    Xa2s_dout[20]/_noR:22   Xa2s_dout[20]/_clk0:10
+	Xa2s_dout[20]/12        Vdd! pmos_2v L=0.18U W=2.16U AD=0.648P
+	 AS=0.324P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+113    Xa2s_dout[20]/_noR:22   Xa2s_dout[20]/clk0:4
+	Xa2s_dout[20]/11        Vdd! pmos_2v L=0.18U W=2.16U AD=0.648P
+	 AS=0.324P PD=0.6U PS=0.3U
MXa2s_dout[20]/M+114    Xa2s_dout[20]/11        clk:3800        Vdd!
+	Vdd! pmos_2v L=0.18U W=2.16U AD=0.324P AS=1.166P PD=0.3U
+	 PS=3.24U
MXa2s_dout[20]/M+115    Vdd!    clk:3797        Xa2s_dout[20]/1:1
+	Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P AS=1.901P PD=0.6U
+	 PS=4.92U
MXa2s_dout[20]/M+98     Vdd!    dout[22].1:3    Xa2s_dout[20]/_R.1:32
+	Vdd! pmos_2v L=0.18U W=4.38U AD=2.365P AS=2.365P PD=5.46U
+	 PS=5.46U
MXa2s_dout[20]/M+89     Xa2s_dout[20]/9:5       Xa2s_dout[20]/Rv:7
+	Vdd!    Vdd! pmos_2v L=0.18U W=0.48U AD=0.259P AS=0.259P
+	 PD=1.56U PS=1.56U
MXa2s_dout[20]/M+90     Xa2s_dout[20]/8:5       Xa2s_dout[20]/_R.1:38
+	Vdd!    Vdd! pmos_2v L=0.18U W=0.48U AD=0.259P AS=0.259P
+	 PD=1.56U PS=1.56U
MXa2s_dout[20]/M+91     Xa2s_dout[20]/PReset:10 _PReset!:6732   Vdd!
+	Vdd! pmos_2v L=0.18U W=1.2U AD=0.648P AS=0.648P PD=2.28U
+	 PS=2.28U
MXa2s_dout[20]/M+92     Xa2s_dout[20]/Rv:10     Xa2s_dout[20]/9:1
+	Vdd!    Vdd! pmos_2v L=0.24U W=0.24U AD=0.302P AS=0.317P
+	 PD=2.28U PS=2.4U
MXa2s_dout[20]/M+93     Xa2s_dout[20]/_R.1:43   Xa2s_dout[20]/8:1
+	Vdd!    Vdd! pmos_2v L=0.24U W=0.24U AD=0.274P AS=0.331P
+	 PD=2.04U PS=2.52U
MXa2s_dout[20]/M+97     dout[22].e:5    Xa2s_dout[20]/_Le:11    Vdd!
+	Vdd! pmos_2v L=0.18U W=2.64U AD=0.792P AS=1.426P PD=0.6U
+	 PS=3.72U
MXa2s_dout[20]/M+96     Vdd!    Xa2s_dout[20]/_Le:16    dout[22].e:5
+	Vdd! pmos_2v L=0.18U W=2.64U AD=0.792P AS=0.792P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+95     Vdd!    Xa2s_dout[20]/_Le:18    dout[22].e:6
+	Vdd! pmos_2v L=0.18U W=2.64U AD=0.792P AS=0.792P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+94     dout[22].e:6    Xa2s_dout[20]/_Le:15    Vdd!
+	Vdd! pmos_2v L=0.18U W=2.64U AD=0.792P AS=1.426P PD=0.6U
+	 PS=3.72U
MXa2s_dout[20]/M+116    Xa2s_dout[20]/0:7       _PReset!:6256   Vdd!
+	Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P AS=1.152P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+117    Xa2s_dout[20]/_clk0:1   clk:3799        
+	Xa2s_dout[20]/0:7       Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P
+	 AS=1.152P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+118    Xa2s_dout[20]/1:2       Xa2s_dout[20]/_R.0:21
+	Xa2s_dout[20]/_clk0:1   Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P
+	 AS=1.152P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+119    Xa2s_dout[20]/_clk0:2   _PReset!:6254   
+	Xa2s_dout[20]/1:2       Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P
+	 AS=1.152P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+127    Vdd!    Xa2s_dout[20]/7:1       
+	Xa2s_dout[20]/__Le:8    Vdd! pmos_2v L=0.24U W=0.24U AD=0.331P
+	 AS=0.274P PD=2.52U PS=2.04U
MXa2s_dout[20]/M+141    Xa2s_dout[20]/_r:13     odq[20]:18      Vdd!
+	Vdd! pmos_2v L=0.18U W=3.06U AD=0.918P AS=0.918P PD=0.6U
+	 PS=0.6U
MXa2s_dout[20]/M+142    Vdd!    Xa2s_dout[20]/_R.0:23   
+	Xa2s_dout[20]/_r:13     Vdd! pmos_2v L=0.18U W=3.06U AD=1.652P
+	 AS=0.918P PD=4.14U PS=0.6U
MXa2s_dout[20]/M+143    Xa2s_dout[20]/__Le:9    Xa2s_dout[20]/Rv:1
+	Vdd!    Vdd! pmos_2v L=0.18U W=2.16U AD=1.166P AS=1.166P
+	 PD=3.24U PS=3.24U
MXa2s_dout[20]/M+125    Vdd!    Xa2s_dout[20]/__Le:3    
+	Xa2s_dout[20]/7:5       Vdd! pmos_2v L=0.18U W=0.48U AD=0.259P
+	 AS=0.259P PD=1.56U PS=1.56U
MXa2s_dout[20]/M+81     Vdd!    oe:176  Xa2s_dout[20]/_grant:6  Vdd!
+	 pmos_2v L=0.18U W=1.2U AD=0.648P AS=0.648P PD=2.28U PS=2.28U
MXa2s_dout[20]/M+120    Xa2s_dout[20]/1:4       Xa2s_dout[20]/_R.1:34
+	Xa2s_dout[20]/_clk0:2   Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P
+	 AS=1.152P PD=0.6U PS=0.6U
MXa2s_dout[20]/M+121    Xa2s_dout[20]/_clk0:4   Xa2s_dout[20]/_noR:25
+	Xa2s_dout[20]/1:4       Vdd! pmos_2v L=0.18U W=3.84U AD=1.901P
+	 AS=1.152P PD=4.92U PS=0.6U
MXa2s_dout[20]/M+122    Vdd!    Xa2s_dout[20]/_noR:26   
+	Xa2s_dout[20]/0:3       Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P
+	 AS=1.901P PD=0.6U PS=4.92U
MXa2s_dout[20]/M+144    Vdd!    Xa2s_dout[20]/__Le:5    
+	Xa2s_dout[20]/_Le:6     Vdd! pmos_2v L=0.18U W=5.52U AD=2.981P
+	 AS=1.656P PD=6.6U PS=0.6U
MXa2s_dout[20]/M+145    Vdd!    _PReset!:6026   Xa2s_dout[20]/_Le:6
+	Vdd! pmos_2v L=0.18U W=5.52U AD=2.981P AS=1.656P PD=6.6U
+	 PS=0.6U
MXa2s_dout[20]/M+123    Xa2s_dout[20]/0:5       Xa2s_dout[20]/_R.1:35
+	Vdd!    Vdd! pmos_2v L=0.18U W=3.84U AD=1.152P AS=1.152P
+	 PD=0.6U PS=0.6U
MXa2s_dout[20]/M+124    Vdd!    Xa2s_dout[20]/_R.0:18   
+	Xa2s_dout[20]/0:5       Vdd! pmos_2v L=0.18U W=3.84U AD=2.074P
+	 AS=1.152P PD=4.92U PS=0.6U
MXa2s_dout[20]/M+126    Xa2s_dout[20]/6:5       Xa2s_dout[20]/_noR:5
+	Vdd!    Vdd! pmos_2v L=0.18U W=0.48U AD=0.259P AS=0.259P
+	 PD=1.56U PS=1.56U
MXa2s_dout[20]/M+128    Xa2s_dout[20]/_noR:10   Xa2s_dout[20]/6:1
+	Vdd!    Vdd! pmos_2v L=0.24U W=0.24U AD=0.302P AS=0.317P
+	 PD=2.28U PS=2.4U
MXa2s_dout[20]/M+129    Xa2s_dout[20]/Rc:5      Xa2s_dout[20]/_noR:13
+	Vdd!    Vdd! pmos_2v L=0.18U W=1.92U AD=1.037P AS=0.576P PD=3U
+	 PS=0.6U
MXa2s_dout[20]/M+130    Xa2s_dout[20]/Rc:6      Xa2s_dout[20]/_R.0:20
+	Vdd!    Vdd! pmos_2v L=0.18U W=1.92U AD=0.576P AS=0.576P
+	 PD=0.6U PS=0.6U
MXa2s_dout[20]/M+131    Vdd!    Xa2s_dout[20]/_R.1:17   
+	Xa2s_dout[20]/Rc:6      Vdd! pmos_2v L=0.18U W=1.92U AD=1.037P
+	 AS=0.576P PD=3U PS=0.6U
MXa2s_dout[20]/M+82     Vdd!    Xa2s_dout[20]/_R.0:32   
+	Xa2s_dout[20]/10:5      Vdd! pmos_2v L=0.18U W=0.48U AD=0.259P
+	 AS=0.259P PD=1.56U PS=1.56U
MXa2s_dout[20]/M+83     Vdd!    Xa2s_dout[20]/10:1      
+	Xa2s_dout[20]/_R.0:35   Vdd! pmos_2v L=0.24U W=0.24U AD=0.331P
+	 AS=0.274P PD=2.52U PS=2.04U
MXa2s_dout[20]/M+85     Xa2s_dout[20]/clk0:24   Xa2s_dout[20]/_clk0:47
+	Vdd!    Vdd! pmos_2v L=0.18U W=1.74U AD=0.522P AS=0.94P
+	 PD=0.6U PS=2.82U
MXa2s_dout[20]/M+84     Vdd!    Xa2s_dout[20]/_clk0:45  
+	Xa2s_dout[20]/clk0:24   Vdd! pmos_2v L=0.18U W=1.74U AD=0.94P
+	 AS=0.522P PD=2.82U PS=0.6U
MXa2s_dout[20]/M+86     Vdd!    clk:4975        Xa2s_dout[20]/_clk:33
+	Vdd! pmos_2v L=0.18U W=3.24U AD=1.75P AS=1.75P PD=4.32U
+	 PS=4.32U
MXa2s_dout[20]/M+87     Xa2s_dout[20]/_clk0:30  Xa2s_dout[20]/clk0:19
+	Vdd!    Vdd! pmos_2v L=0.24U W=0.24U AD=0.274P AS=0.36P
+	 PD=2.04U PS=2.76U
MXa2s_dout[20]/M+88     Vdd!    dout[22].0:2    Xa2s_dout[20]/_R.0:25
+	Vdd! pmos_2v L=0.18U W=3.18U AD=1.717P AS=1.717P PD=4.26U
+	 PS=4.26U
Rg66091 Xa2s_dout[22]/Rv:1      Xa2s_dout[22]/Rv:2 84.3517 $cpoly
Rg66092 Xa2s_dout[21]/Rv:1      Xa2s_dout[21]/Rv:2 84.3517 $cpoly
Rg66093 Xa2s_dout[20]/Rv:1      Xa2s_dout[20]/Rv:2 84.3517 $cpoly
Rg66094 Xa2s_dout[19]/Rv:1      Xa2s_dout[19]/Rv:2 84.3517 $cpoly
Rg66095 Xa2s_dout[18]/Rv:1      Xa2s_dout[18]/Rv:2 84.3517 $cpoly
Rg66140 Xa2s_dout[22]/6:1       Xa2s_dout[22]/6:2 8.7495 $cpoly
Rg66141 Xa2s_dout[21]/6:1       Xa2s_dout[21]/6:2 8.7495 $cpoly
Rg66142 Xa2s_dout[20]/6:1       Xa2s_dout[20]/6:2 8.7495 $cpoly
Rg66143 Xa2s_dout[19]/6:1       Xa2s_dout[19]/6:2 8.7495 $cpoly
Rg66144 Xa2s_dout[18]/6:1       Xa2s_dout[18]/6:2 8.7495 $cpoly
Rg66172 Xa2s_dout[22]/7:1       Xa2s_dout[22]/7:2 11.8495 $cpoly
Rg66173 Xa2s_dout[21]/7:1       Xa2s_dout[21]/7:2 11.8495 $cpoly
Rg66174 Xa2s_dout[20]/7:1       Xa2s_dout[20]/7:2 11.8495 $cpoly
Rg66175 Xa2s_dout[19]/7:1       Xa2s_dout[19]/7:2 11.8495 $cpoly
Rg66176 Xa2s_dout[18]/7:1       Xa2s_dout[18]/7:2 11.8495 $cpoly
Rg66303 Xa2s_dout[21]/_noR:4    Xa2s_dout[21]/_noR:5 23.9733 $cpoly
Rg66304 Xa2s_dout[21]/_noR:4    Xa2s_dout[21]/_noR:8 16.6712 $cpoly
Rg66305 Xa2s_dout[20]/__Le:1    Xa2s_dout[20]/__Le:2 23.9733 $cpoly
Rg66306 Xa2s_dout[20]/__Le:2    Xa2s_dout[20]/__Le:3 23.9733 $cpoly
Rg66307 Xa2s_dout[20]/__Le:2    Xa2s_dout[20]/__Le:4 16.6712 $cpoly
Rg66308 Xa2s_dout[20]/_noR:3    Xa2s_dout[20]/_noR:4 23.9733 $cpoly
Rg66309 Xa2s_dout[20]/_noR:4    Xa2s_dout[20]/_noR:5 23.9733 $cpoly
Rg66310 Xa2s_dout[20]/_noR:4    Xa2s_dout[20]/_noR:8 16.6712 $cpoly
Rg66311 Xa2s_dout[19]/__Le:1    Xa2s_dout[19]/__Le:2 23.9733 $cpoly
Rg66312 Xa2s_dout[19]/__Le:2    Xa2s_dout[19]/__Le:3 23.9733 $cpoly
Rg66444 Xa2s_dout[22]/_R.0:1    Xa2s_dout[22]/_R.0:3 140.1517 $cpoly
Rg66445 Xa2s_dout[21]/_R.0:1    Xa2s_dout[21]/_R.0:3 140.1517 $cpoly
Rg66446 Xa2s_dout[20]/_R.0:1    Xa2s_dout[20]/_R.0:3 140.1517 $cpoly
Rg66447 Xa2s_dout[19]/_R.0:1    Xa2s_dout[19]/_R.0:3 140.1517 $cpoly
Rg66448 Xa2s_dout[18]/_R.0:1    Xa2s_dout[18]/_R.0:3 140.1517 $cpoly
Rg66476 Xa2s_dout[22]/6:3       Xa2s_dout[22]/6:6 3.4068 $cpoly
Rg66477 Xa2s_dout[21]/6:3       Xa2s_dout[21]/6:6 3.4068 $cpoly
Rg66478 Xa2s_dout[20]/6:3       Xa2s_dout[20]/6:6 3.4068 $cpoly
Rg66479 Xa2s_dout[19]/6:3       Xa2s_dout[19]/6:6 3.4068 $cpoly
Rg66480 Xa2s_dout[18]/6:3       Xa2s_dout[18]/6:6 3.4068 $cpoly
Rg66530 Xa2s_dout[21]/_noR:12   Xa2s_dout[21]/_noR:13 48.0869 $cpoly
Rg66531 Xa2s_dout[21]/_noR:12   Xa2s_dout[21]/_noR:1 30.5776 $cpoly
Rg66532 Xa2s_dout[20]/_noR:11   Xa2s_dout[20]/_noR:12 49.1202 $cpoly
Rg66533 Xa2s_dout[20]/_noR:12   Xa2s_dout[20]/_noR:13 48.0869 $cpoly
Rg66534 Xa2s_dout[20]/_noR:12   Xa2s_dout[20]/_noR:1 30.5776 $cpoly
Rg66535 Xa2s_dout[19]/_noR:11   Xa2s_dout[19]/_noR:12 49.1202 $cpoly
Rg66536 Xa2s_dout[19]/_noR:12   Xa2s_dout[19]/_noR:13 48.0869 $cpoly
Rg66604 Xa2s_dout[22]/7:6       Xa2s_dout[22]/7:3 5.8022 $cpoly
Rg66605 Xa2s_dout[21]/7:6       Xa2s_dout[21]/7:3 5.8022 $cpoly
Rg66606 Xa2s_dout[20]/7:6       Xa2s_dout[20]/7:3 5.8022 $cpoly
Rg66607 Xa2s_dout[19]/7:6       Xa2s_dout[19]/7:3 5.8022 $cpoly
Rg66608 Xa2s_dout[18]/7:6       Xa2s_dout[18]/7:3 5.8022 $cpoly
Rg66663 Xa2s_dout[21]/_r:1      Xa2s_dout[21]/_r:2 127.8179 $cpoly
Rg66664 Xa2s_dout[21]/_r:2      Xa2s_dout[21]/_r:3 49.5235 $cpoly
Rg66665 Xa2s_dout[20]/_r:1      Xa2s_dout[20]/_r:2 127.8179 $cpoly
Rg66666 Xa2s_dout[20]/_r:2      Xa2s_dout[20]/_r:3 49.5235 $cpoly
Rg66667 Xa2s_dout[19]/_r:1      Xa2s_dout[19]/_r:2 127.8179 $cpoly
Rg66668 Xa2s_dout[19]/_r:2      Xa2s_dout[19]/_r:3 49.5235 $cpoly
Rg66749 Xa2s_dout[21]/_r:7      Xa2s_dout[21]/_r:8 117.4846 $cpoly
Rg66750 Xa2s_dout[21]/_r:8      Xa2s_dout[21]/_r:9 49.5235 $cpoly
Rg66751 Xa2s_dout[20]/_r:4      Xa2s_dout[20]/_r:5 117.4846 $cpoly
Rg66752 Xa2s_dout[20]/_r:5      Xa2s_dout[20]/_r:6 49.5235 $cpoly
Rg66753 Xa2s_dout[20]/_r:7      Xa2s_dout[20]/_r:8 117.4846 $cpoly
Rg66754 Xa2s_dout[20]/_r:8      Xa2s_dout[20]/_r:9 49.5235 $cpoly
Rg66755 Xa2s_dout[19]/_r:4      Xa2s_dout[19]/_r:5 117.4846 $cpoly
Rg66756 Xa2s_dout[19]/_r:5      Xa2s_dout[19]/_r:6 49.5235 $cpoly
Rg66855 Xa2s_dout[21]/_r:10     Xa2s_dout[21]/_r:11 112.6230 $cpoly
Rg66856 Xa2s_dout[21]/_r:11     Xa2s_dout[21]/_r:12 49.5235 $cpoly
Rg66857 Xa2s_dout[20]/_r:10     Xa2s_dout[20]/_r:11 112.6230 $cpoly
Rg66858 Xa2s_dout[20]/_r:11     Xa2s_dout[20]/_r:12 49.5235 $cpoly
Rg66859 Xa2s_dout[19]/_r:10     Xa2s_dout[19]/_r:11 112.6230 $cpoly
Rg66860 Xa2s_dout[19]/_r:11     Xa2s_dout[19]/_r:12 49.5235 $cpoly
Rg67059 Xa2s_dout[21]/_R.1:10   Xa2s_dout[21]/_R.1:11 52.6235 $cpoly
Rg67060 Xa2s_dout[21]/_R.1:11   Xa2s_dout[21]/_R.1:12 127.8179 $cpoly
Rg67061 Xa2s_dout[20]/_R.1:1    Xa2s_dout[20]/_R.1:2 52.6235 $cpoly
Rg67062 Xa2s_dout[20]/_R.1:2    Xa2s_dout[20]/_R.1:3 117.4846 $cpoly
Rg67063 Xa2s_dout[20]/_R.1:4    Xa2s_dout[20]/_R.1:5 52.6235 $cpoly
Rg67064 Xa2s_dout[20]/_R.1:5    Xa2s_dout[20]/_R.1:6 112.6230 $cpoly
Rg67065 Xa2s_dout[20]/_R.1:7    Xa2s_dout[20]/_R.1:8 52.6235 $cpoly
Rg67066 Xa2s_dout[20]/_R.1:8    Xa2s_dout[20]/_R.1:9 117.4846 $cpoly
Rg67067 Xa2s_dout[20]/_R.1:10   Xa2s_dout[20]/_R.1:11 52.6235 $cpoly
Rg67068 Xa2s_dout[20]/_R.1:11   Xa2s_dout[20]/_R.1:12 127.8179 $cpoly
Rg67069 Xa2s_dout[19]/_R.1:1    Xa2s_dout[19]/_R.1:2 52.6235 $cpoly
Rg67070 Xa2s_dout[19]/_R.1:2    Xa2s_dout[19]/_R.1:3 117.4846 $cpoly
Rg67238 Xa2s_dout[22]/_R.1:13   Xa2s_dout[22]/_R.1:14 114.5237 $cpoly
Rg67239 Xa2s_dout[21]/_R.1:13   Xa2s_dout[21]/_R.1:14 114.5237 $cpoly
Rg67240 Xa2s_dout[20]/_R.1:13   Xa2s_dout[20]/_R.1:14 114.5237 $cpoly
Rg67241 Xa2s_dout[19]/_R.1:13   Xa2s_dout[19]/_R.1:14 114.5237 $cpoly
Rg67242 Xa2s_dout[18]/_R.1:13   Xa2s_dout[18]/_R.1:14 114.5237 $cpoly
Rg67281 Xa2s_dout[21]/_R.1:15   Xa2s_dout[21]/_R.1:16 68.8826 $cpoly
Rg67282 Xa2s_dout[21]/_R.1:16   Xa2s_dout[21]/_R.1:17 113.3512 $cpoly
Rg67283 Xa2s_dout[20]/_R.1:15   Xa2s_dout[20]/_R.1:16 68.8826 $cpoly
Rg67284 Xa2s_dout[20]/_R.1:16   Xa2s_dout[20]/_R.1:17 113.3512 $cpoly
Rg67285 Xa2s_dout[19]/_R.1:15   Xa2s_dout[19]/_R.1:16 68.8826 $cpoly
Rg67286 Xa2s_dout[19]/_R.1:16   Xa2s_dout[19]/_R.1:17 113.3512 $cpoly
Rg67381 Xa2s_dout[21]/__Le:5    Xa2s_dout[21]/__Le:6 181.5512 $cpoly
Rg67382 Xa2s_dout[21]/__Le:6    Xa2s_dout[21]/__Le:7 94.0159 $cpoly
Rg67383 Xa2s_dout[20]/__Le:5    Xa2s_dout[20]/__Le:6 181.5512 $cpoly
Rg67384 Xa2s_dout[20]/__Le:6    Xa2s_dout[20]/__Le:7 94.0159 $cpoly
Rg67385 Xa2s_dout[19]/__Le:5    Xa2s_dout[19]/__Le:6 181.5512 $cpoly
Rg67386 Xa2s_dout[19]/__Le:6    Xa2s_dout[19]/__Le:7 94.0159 $cpoly
Rg68373 Xa2s_dout[22]/_R.1:18   Xa2s_dout[22]/_R.1:29 77.1492 $cpoly
Rg68374 Xa2s_dout[21]/_R.1:18   Xa2s_dout[21]/_R.1:29 77.1492 $cpoly
Rg68375 Xa2s_dout[20]/_R.1:18   Xa2s_dout[20]/_R.1:29 77.1492 $cpoly
Rg68376 Xa2s_dout[19]/_R.1:18   Xa2s_dout[19]/_R.1:29 77.1492 $cpoly
Rg68377 Xa2s_dout[18]/_R.1:18   Xa2s_dout[18]/_R.1:29 77.1492 $cpoly
Rg68405 Xa2s_dout[22]/_r:19     Xa2s_dout[22]/_r:17 54.6902 $cpoly
Rg68406 Xa2s_dout[21]/_r:19     Xa2s_dout[21]/_r:17 54.6902 $cpoly
Rg68407 Xa2s_dout[20]/_r:19     Xa2s_dout[20]/_r:17 54.6902 $cpoly
Rg68408 Xa2s_dout[19]/_r:19     Xa2s_dout[19]/_r:17 54.6902 $cpoly
Rg68409 Xa2s_dout[18]/_r:19     Xa2s_dout[18]/_r:17 54.6902 $cpoly
Rg68437 Xa2s_dout[22]/_r:20     Xa2s_dout[22]/_r:18 100.5210 $cpoly
Rg68438 Xa2s_dout[21]/_r:20     Xa2s_dout[21]/_r:18 100.5210 $cpoly
Rg68439 Xa2s_dout[20]/_r:20     Xa2s_dout[20]/_r:18 100.5210 $cpoly
Rg68440 Xa2s_dout[19]/_r:20     Xa2s_dout[19]/_r:18 100.5210 $cpoly
Rg68441 Xa2s_dout[18]/_r:20     Xa2s_dout[18]/_r:18 100.5210 $cpoly
Rg68469 Xa2s_dout[22]/_R.0:13   Xa2s_dout[22]/_R.0:9 80.4418 $cpoly
Rg68470 Xa2s_dout[21]/_R.0:13   Xa2s_dout[21]/_R.0:9 80.4418 $cpoly
Rg68471 Xa2s_dout[20]/_R.0:13   Xa2s_dout[20]/_R.0:9 80.4418 $cpoly
Rg68472 Xa2s_dout[19]/_R.0:13   Xa2s_dout[19]/_R.0:9 80.4418 $cpoly
Rg68473 Xa2s_dout[18]/_R.0:13   Xa2s_dout[18]/_R.0:9 80.4418 $cpoly
Rg68651 Xa2s_dout[21]/_clk:4    Xa2s_dout[21]/_clk:1 53.3798 $cpoly
Rg68652 Xa2s_dout[21]/_clk:4    Xa2s_dout[21]/_clk:5 60.6793 $cpoly
Rg68653 Xa2s_dout[20]/_clk:3    Xa2s_dout[20]/_clk:4 95.1847 $cpoly
Rg68654 Xa2s_dout[20]/_clk:4    Xa2s_dout[20]/_clk:1 53.3798 $cpoly
Rg68655 Xa2s_dout[20]/_clk:4    Xa2s_dout[20]/_clk:5 60.6793 $cpoly
Rg68656 Xa2s_dout[19]/_clk:3    Xa2s_dout[19]/_clk:4 95.1847 $cpoly
Rg68657 Xa2s_dout[19]/_clk:4    Xa2s_dout[19]/_clk:1 53.3798 $cpoly
Rg69166 Xa2s_dout[22]/_R.0:14   Xa2s_dout[22]/_R.0:17 154.2543 $cpoly
Rg69167 Xa2s_dout[21]/_R.0:14   Xa2s_dout[21]/_R.0:17 154.2543 $cpoly
Rg69168 Xa2s_dout[20]/_R.0:14   Xa2s_dout[20]/_R.0:17 154.2543 $cpoly
Rg69169 Xa2s_dout[19]/_R.0:14   Xa2s_dout[19]/_R.0:17 154.2543 $cpoly
Rg69170 Xa2s_dout[18]/_R.0:14   Xa2s_dout[18]/_R.0:17 154.2543 $cpoly
Rg69510 Xa2s_dout[21]/clk0:1    Xa2s_dout[21]/clk0:2 92.6184 $cpoly
Rg69511 Xa2s_dout[21]/clk0:3    Xa2s_dout[21]/clk0:4 81.5568 $cpoly
Rg69512 Xa2s_dout[20]/_R.1:30   Xa2s_dout[20]/_R.1:31 96.0235 $cpoly
Rg69513 Xa2s_dout[20]/clk0:1    Xa2s_dout[20]/clk0:2 92.6184 $cpoly
Rg69514 Xa2s_dout[20]/clk0:3    Xa2s_dout[20]/clk0:4 81.5568 $cpoly
Rg69515 Xa2s_dout[19]/_R.1:30   Xa2s_dout[19]/_R.1:31 96.0235 $cpoly
Rg69516 Xa2s_dout[19]/clk0:1    Xa2s_dout[19]/clk0:2 92.6184 $cpoly
Rg69740 Xa2s_dout[21]/_R.1:34   Xa2s_dout[21]/_R.1:22 185.2543 $cpoly
Rg69741 Xa2s_dout[21]/_R.1:22   Xa2s_dout[21]/_R.1:35 121.1876 $cpoly
Rg69742 Xa2s_dout[20]/_R.1:34   Xa2s_dout[20]/_R.1:22 185.2543 $cpoly
Rg69743 Xa2s_dout[20]/_R.1:22   Xa2s_dout[20]/_R.1:35 121.1876 $cpoly
Rg69744 Xa2s_dout[19]/_R.1:34   Xa2s_dout[19]/_R.1:22 185.2543 $cpoly
Rg69745 Xa2s_dout[19]/_R.1:22   Xa2s_dout[19]/_R.1:35 121.1876 $cpoly
Rg69826 Xa2s_dout[21]/_R.0:4    Xa2s_dout[21]/_R.0:19 109.8210 $cpoly
Rg69827 Xa2s_dout[21]/_R.0:19   Xa2s_dout[21]/_R.0:20 103.0179 $cpoly
Rg69828 Xa2s_dout[20]/_R.0:18   Xa2s_dout[20]/_R.0:12 132.8524 $cpoly
Rg69829 Xa2s_dout[20]/_R.0:12   Xa2s_dout[20]/_R.0:4 123.0742 $cpoly
Rg69830 Xa2s_dout[20]/_R.0:4    Xa2s_dout[20]/_R.0:19 109.8210 $cpoly
Rg69831 Xa2s_dout[20]/_R.0:19   Xa2s_dout[20]/_R.0:20 103.0179 $cpoly
Rg69832 Xa2s_dout[19]/_R.0:18   Xa2s_dout[19]/_R.0:12 132.8524 $cpoly
Rg69833 Xa2s_dout[19]/_R.0:12   Xa2s_dout[19]/_R.0:4 123.0742 $cpoly
Rg69943 Xa2s_dout[21]/_R.0:11   Xa2s_dout[21]/_R.0:22 144.6492 $cpoly
Rg69944 Xa2s_dout[21]/_R.0:22   Xa2s_dout[21]/_R.0:23 179.4846 $cpoly
Rg69945 Xa2s_dout[20]/_R.0:21   Xa2s_dout[20]/_R.0:11 120.8235 $cpoly
Rg69946 Xa2s_dout[20]/_R.0:11   Xa2s_dout[20]/_R.0:22 144.6492 $cpoly
Rg69947 Xa2s_dout[20]/_R.0:22   Xa2s_dout[20]/_R.0:23 179.4846 $cpoly
Rg69948 Xa2s_dout[19]/_R.0:21   Xa2s_dout[19]/_R.0:11 120.8235 $cpoly
Rg69949 Xa2s_dout[19]/_R.0:11   Xa2s_dout[19]/_R.0:22 144.6492 $cpoly
Rg70228 Xa2s_dout[21]/_clk0:8   Xa2s_dout[21]/_clk0:9 78.4176 $cpoly
Rg70229 Xa2s_dout[21]/_clk0:8   Xa2s_dout[21]/_clk0:10 78.4176 $cpoly
Rg70230 Xa2s_dout[20]/_clk0:7   Xa2s_dout[20]/_clk0:8 87.7751 $cpoly
Rg70231 Xa2s_dout[20]/_clk0:8   Xa2s_dout[20]/_clk0:9 78.4176 $cpoly
Rg70232 Xa2s_dout[20]/_clk0:8   Xa2s_dout[20]/_clk0:10 78.4176 $cpoly
Rg70233 Xa2s_dout[19]/_clk0:7   Xa2s_dout[19]/_clk0:8 87.7751 $cpoly
Rg70234 Xa2s_dout[19]/_clk0:8   Xa2s_dout[19]/_clk0:9 78.4176 $cpoly
Rg70381 Xa2s_dout[21]/_noR:23   Xa2s_dout[21]/_noR:17 14.0443 $cpoly
Rg70382 Xa2s_dout[21]/_noR:24   Xa2s_dout[21]/_noR:26 88.4306 $cpoly
Rg70383 Xa2s_dout[20]/_noR:17   Xa2s_dout[20]/_noR:23 84.1874 $cpoly
Rg70384 Xa2s_dout[20]/_noR:23   Xa2s_dout[20]/_noR:24 42.1900 $cpoly
Rg70385 Xa2s_dout[20]/_noR:24   Xa2s_dout[20]/_noR:25 116.4746 $cpoly
Rg70386 Xa2s_dout[20]/_noR:23   Xa2s_dout[20]/_noR:17 14.0443 $cpoly
Rg70387 Xa2s_dout[20]/_noR:24   Xa2s_dout[20]/_noR:26 88.4306 $cpoly
Rg70388 Xa2s_dout[19]/_noR:17   Xa2s_dout[19]/_noR:23 84.1874 $cpoly
Rg70389 Xa2s_dout[19]/_noR:23   Xa2s_dout[19]/_noR:24 42.1900 $cpoly
Rg70741 Xa2s_dout[22]/Rv:3      Xa2s_dout[22]/Rv:4 72.9851 $cpoly
Rg70742 Xa2s_dout[21]/Rv:3      Xa2s_dout[21]/Rv:4 72.9851 $cpoly
Rg70743 Xa2s_dout[20]/Rv:3      Xa2s_dout[20]/Rv:4 72.9851 $cpoly
Rg70744 Xa2s_dout[19]/Rv:3      Xa2s_dout[19]/Rv:4 72.9851 $cpoly
Rg70745 Xa2s_dout[18]/Rv:3      Xa2s_dout[18]/Rv:4 72.9851 $cpoly
Rg70773 Xa2s_dout[22]/_clk0:11  Xa2s_dout[22]/_clk0:12 103.5211 $cpoly
Rg70774 Xa2s_dout[21]/_clk0:11  Xa2s_dout[21]/_clk0:12 103.5211 $cpoly
Rg70775 Xa2s_dout[20]/_clk0:11  Xa2s_dout[20]/_clk0:12 103.5211 $cpoly
Rg70776 Xa2s_dout[19]/_clk0:11  Xa2s_dout[19]/_clk0:12 103.5211 $cpoly
Rg70777 Xa2s_dout[18]/_clk0:11  Xa2s_dout[18]/_clk0:12 103.5211 $cpoly
Rg71007 Xa2s_dout[22]/clk0:9    Xa2s_dout[22]/clk0:11 46.4235 $cpoly
Rg71008 Xa2s_dout[21]/clk0:9    Xa2s_dout[21]/clk0:11 46.4235 $cpoly
Rg71009 Xa2s_dout[20]/clk0:9    Xa2s_dout[20]/clk0:11 46.4235 $cpoly
Rg71010 Xa2s_dout[19]/clk0:9    Xa2s_dout[19]/clk0:11 46.4235 $cpoly
Rg71011 Xa2s_dout[18]/clk0:9    Xa2s_dout[18]/clk0:11 46.4235 $cpoly
Rg71041 Xa2s_dout[22]/_clk:14   Xa2s_dout[22]/_clk:7 48.4902 $cpoly
Rg71042 Xa2s_dout[21]/_clk:14   Xa2s_dout[21]/_clk:7 48.4902 $cpoly
Rg71043 Xa2s_dout[20]/_clk:14   Xa2s_dout[20]/_clk:7 48.4902 $cpoly
Rg71044 Xa2s_dout[19]/_clk:14   Xa2s_dout[19]/_clk:7 48.4902 $cpoly
Rg71045 Xa2s_dout[18]/_clk:14   Xa2s_dout[18]/_clk:7 48.4902 $cpoly
Rg71310 Xa2s_dout[22]/9:1       Xa2s_dout[22]/9:2 8.7495 $cpoly
Rg71311 Xa2s_dout[21]/9:1       Xa2s_dout[21]/9:2 8.7495 $cpoly
Rg71312 Xa2s_dout[20]/9:1       Xa2s_dout[20]/9:2 8.7495 $cpoly
Rg71313 Xa2s_dout[19]/9:1       Xa2s_dout[19]/9:2 8.7495 $cpoly
Rg71314 Xa2s_dout[18]/9:1       Xa2s_dout[18]/9:2 8.7495 $cpoly
Rg71342 Xa2s_dout[22]/8:1       Xa2s_dout[22]/8:2 11.8495 $cpoly
Rg71343 Xa2s_dout[21]/8:1       Xa2s_dout[21]/8:2 11.8495 $cpoly
Rg71344 Xa2s_dout[20]/8:1       Xa2s_dout[20]/8:2 11.8495 $cpoly
Rg71345 Xa2s_dout[19]/8:1       Xa2s_dout[19]/8:2 11.8495 $cpoly
Rg71346 Xa2s_dout[18]/8:1       Xa2s_dout[18]/8:2 11.8495 $cpoly

Rg71918 Xa2s_dout[22]/_clk:17   Xa2s_dout[22]/_clk:11 113.9543 $cpoly
Rg71919 Xa2s_dout[21]/_clk:17   Xa2s_dout[21]/_clk:11 113.9543 $cpoly
Rg71920 Xa2s_dout[20]/_clk:17   Xa2s_dout[20]/_clk:11 113.9543 $cpoly
Rg71921 Xa2s_dout[19]/_clk:17   Xa2s_dout[19]/_clk:11 113.9543 $cpoly
Rg71922 Xa2s_dout[18]/_clk:17   Xa2s_dout[18]/_clk:11 113.9543 $cpoly

Rg71950 Xa2s_dout[22]/_clk0:13  Xa2s_dout[22]/_clk0:14 112.5568 $cpoly
Rg71951 Xa2s_dout[21]/_clk0:13  Xa2s_dout[21]/_clk0:14 112.5568 $cpoly
Rg71952 Xa2s_dout[20]/_clk0:13  Xa2s_dout[20]/_clk0:14 112.5568 $cpoly
Rg71953 Xa2s_dout[19]/_clk0:13  Xa2s_dout[19]/_clk0:14 112.5568 $cpoly
Rg71954 Xa2s_dout[18]/_clk0:13  Xa2s_dout[18]/_clk0:14 112.5568 $cpoly

Rg72208 Xa2s_dout[21]/PReset:7  Xa2s_dout[21]/PReset:1 13.8209 $cpoly
Rg72209 Xa2s_dout[21]/PReset:7  Xa2s_dout[21]/PReset:8 53.3771 $cpoly
Rg72210 Xa2s_dout[20]/PReset:6  Xa2s_dout[20]/PReset:7 106.3176 $cpoly
Rg72211 Xa2s_dout[20]/PReset:7  Xa2s_dout[20]/PReset:1 13.8209 $cpoly
Rg72212 Xa2s_dout[20]/PReset:7  Xa2s_dout[20]/PReset:8 53.3771 $cpoly
Rg72213 Xa2s_dout[19]/PReset:6  Xa2s_dout[19]/PReset:7 106.3176 $cpoly
Rg72214 Xa2s_dout[19]/PReset:7  Xa2s_dout[19]/PReset:1 13.8209 $cpoly

Rg72337 Xa2s_dout[21]/_R.1:37   Xa2s_dout[21]/_R.1:38 23.9733 $cpoly
Rg72338 Xa2s_dout[21]/_R.1:37   Xa2s_dout[21]/_R.1:39 16.6712 $cpoly
Rg72339 Xa2s_dout[20]/Rv:5      Xa2s_dout[20]/Rv:6 23.9733 $cpoly
Rg72340 Xa2s_dout[20]/Rv:6      Xa2s_dout[20]/Rv:7 23.9733 $cpoly
Rg72341 Xa2s_dout[20]/Rv:6      Xa2s_dout[20]/Rv:8 16.6712 $cpoly
Rg72342 Xa2s_dout[20]/_R.1:36   Xa2s_dout[20]/_R.1:37 23.9733 $cpoly
Rg72343 Xa2s_dout[20]/_R.1:37   Xa2s_dout[20]/_R.1:38 23.9733 $cpoly
Rg72344 Xa2s_dout[20]/_R.1:37   Xa2s_dout[20]/_R.1:39 16.6712 $cpoly
Rg72345 Xa2s_dout[19]/Rv:5      Xa2s_dout[19]/Rv:6 23.9733 $cpoly
Rg72346 Xa2s_dout[19]/Rv:6      Xa2s_dout[19]/Rv:7 23.9733 $cpoly

Rg72474 Xa2s_dout[22]/Rc:7      Xa2s_dout[22]/Rc:8 72.6210 $cpoly
Rg72475 Xa2s_dout[21]/Rc:7      Xa2s_dout[21]/Rc:8 72.6210 $cpoly
Rg72476 Xa2s_dout[20]/Rc:7      Xa2s_dout[20]/Rc:8 72.6210 $cpoly
Rg72477 Xa2s_dout[19]/Rc:7      Xa2s_dout[19]/Rc:8 72.6210 $cpoly
Rg72478 Xa2s_dout[18]/Rc:7      Xa2s_dout[18]/Rc:8 72.6210 $cpoly

Rg72516 Xa2s_dout[22]/_clk:18   Xa2s_dout[22]/_clk:9 114.6235 $cpoly
Rg72517 Xa2s_dout[21]/_clk:18   Xa2s_dout[21]/_clk:9 114.6235 $cpoly
Rg72518 Xa2s_dout[20]/_clk:18   Xa2s_dout[20]/_clk:9 114.6235 $cpoly
Rg72519 Xa2s_dout[19]/_clk:18   Xa2s_dout[19]/_clk:9 114.6235 $cpoly
Rg72520 Xa2s_dout[18]/_clk:18   Xa2s_dout[18]/_clk:9 114.6235 $cpoly

Rg72548 Xa2s_dout[22]/_clk0:15  Xa2s_dout[22]/_clk0:16 47.4568 $cpoly
Rg72549 Xa2s_dout[21]/_clk0:15  Xa2s_dout[21]/_clk0:16 47.4568 $cpoly
Rg72550 Xa2s_dout[20]/_clk0:15  Xa2s_dout[20]/_clk0:16 47.4568 $cpoly
Rg72551 Xa2s_dout[19]/_clk0:15  Xa2s_dout[19]/_clk0:16 47.4568 $cpoly
Rg72552 Xa2s_dout[18]/_clk0:15  Xa2s_dout[18]/_clk0:16 47.4568 $cpoly

Rg72580 Xa2s_dout[22]/clk0:12   Xa2s_dout[22]/clk0:14 71.5876 $cpoly
Rg72581 Xa2s_dout[21]/clk0:12   Xa2s_dout[21]/clk0:14 71.5876 $cpoly
Rg72582 Xa2s_dout[20]/clk0:12   Xa2s_dout[20]/clk0:14 71.5876 $cpoly
Rg72583 Xa2s_dout[19]/clk0:12   Xa2s_dout[19]/clk0:14 71.5876 $cpoly
Rg72584 Xa2s_dout[18]/clk0:12   Xa2s_dout[18]/clk0:14 71.5876 $cpoly

Rg72682 Xa2s_dout[22]/Rc:9      Xa2s_dout[22]/Rc:12 73.2902 $cpoly
Rg72683 Xa2s_dout[21]/Rc:9      Xa2s_dout[21]/Rc:12 73.2902 $cpoly
Rg72684 Xa2s_dout[20]/Rc:9      Xa2s_dout[20]/Rc:12 73.2902 $cpoly
Rg72685 Xa2s_dout[19]/Rc:9      Xa2s_dout[19]/Rc:12 73.2902 $cpoly
Rg72686 Xa2s_dout[18]/Rc:9      Xa2s_dout[18]/Rc:12 73.2902 $cpoly

Rg72743 Xa2s_dout[22]/9:3       Xa2s_dout[22]/9:6 3.0428 $cpoly
Rg72744 Xa2s_dout[21]/9:3       Xa2s_dout[21]/9:6 3.0428 $cpoly
Rg72745 Xa2s_dout[20]/9:3       Xa2s_dout[20]/9:6 3.0428 $cpoly
Rg72746 Xa2s_dout[19]/9:3       Xa2s_dout[19]/9:6 3.0428 $cpoly
Rg72747 Xa2s_dout[18]/9:3       Xa2s_dout[18]/9:6 3.0428 $cpoly

Rg72819 Xa2s_dout[22]/8:6       Xa2s_dout[22]/8:3 5.8022 $cpoly
Rg72820 Xa2s_dout[21]/8:6       Xa2s_dout[21]/8:3 5.8022 $cpoly
Rg72821 Xa2s_dout[20]/8:6       Xa2s_dout[20]/8:3 5.8022 $cpoly
Rg72822 Xa2s_dout[19]/8:6       Xa2s_dout[19]/8:3 5.8022 $cpoly
Rg72823 Xa2s_dout[18]/8:6       Xa2s_dout[18]/8:3 5.8022 $cpoly

Rg72888 Xa2s_dout[21]/_grant:3  Xa2s_dout[21]/_grant:4 112.6412 $cpoly
Rg72889 Xa2s_dout[21]/_grant:3  Xa2s_dout[21]/_grant:5 47.0535 $cpoly
Rg72890 Xa2s_dout[20]/_grant:1  Xa2s_dout[20]/_grant:3 58.3540 $cpoly
Rg72891 Xa2s_dout[20]/_grant:3  Xa2s_dout[20]/_grant:4 112.6412 $cpoly
Rg72892 Xa2s_dout[20]/_grant:3  Xa2s_dout[20]/_grant:5 47.0535 $cpoly
Rg72893 Xa2s_dout[19]/_grant:1  Xa2s_dout[19]/_grant:3 58.3540 $cpoly
Rg72894 Xa2s_dout[19]/_grant:3  Xa2s_dout[19]/_grant:4 112.6412 $cpoly

Rg73108 Xa2s_dout[21]/_Le:13    Xa2s_dout[21]/_Le:19 58.7151 $cpoly
Rg73109 Xa2s_dout[21]/_Le:14    Xa2s_dout[21]/_Le:20 60.1643 $cpoly
Rg73110 Xa2s_dout[20]/_Le:9     Xa2s_dout[20]/_Le:10 60.1643 $cpoly
Rg73111 Xa2s_dout[20]/_Le:10    Xa2s_dout[20]/_Le:11 59.1310 $cpoly
Rg73112 Xa2s_dout[20]/_Le:10    Xa2s_dout[20]/_Le:12 7.8538 $cpoly
Rg73113 Xa2s_dout[20]/_Le:12    Xa2s_dout[20]/_Le:7 6.1036 $cpoly
Rg73114 Xa2s_dout[20]/_Le:7     Xa2s_dout[20]/_Le:13 1.3544 $cpoly
Rg73115 Xa2s_dout[20]/_Le:13    Xa2s_dout[20]/_Le:7 5.2294 $cpoly
Rg73116 Xa2s_dout[20]/_Le:7     Xa2s_dout[20]/_Le:14 0.2788 $cpoly
Rg73117 Xa2s_dout[20]/_Le:14    Xa2s_dout[20]/_Le:15 59.1310 $cpoly
Rg73118 Xa2s_dout[20]/_Le:12    Xa2s_dout[20]/_Le:16 57.6818 $cpoly
Rg73119 Xa2s_dout[20]/_Le:12    Xa2s_dout[20]/_Le:17 58.7151 $cpoly
Rg73120 Xa2s_dout[20]/_Le:13    Xa2s_dout[20]/_Le:18 57.6818 $cpoly
Rg73121 Xa2s_dout[20]/_Le:13    Xa2s_dout[20]/_Le:19 58.7151 $cpoly
Rg73122 Xa2s_dout[20]/_Le:14    Xa2s_dout[20]/_Le:20 60.1643 $cpoly
Rg73123 Xa2s_dout[19]/_Le:9     Xa2s_dout[19]/_Le:10 60.1643 $cpoly
Rg73124 Xa2s_dout[19]/_Le:10    Xa2s_dout[19]/_Le:11 59.1310 $cpoly

Rg73530 Xa2s_dout[22]/clk0:15   Xa2s_dout[22]/clk0:16 118.4517 $cpoly
Rg73531 Xa2s_dout[21]/clk0:15   Xa2s_dout[21]/clk0:16 118.4517 $cpoly
Rg73532 Xa2s_dout[20]/clk0:15   Xa2s_dout[20]/clk0:16 118.4517 $cpoly
Rg73533 Xa2s_dout[19]/clk0:15   Xa2s_dout[19]/clk0:16 118.4517 $cpoly
Rg73534 Xa2s_dout[18]/clk0:15   Xa2s_dout[18]/clk0:16 118.4517 $cpoly

Rg73665 Xa2s_dout[22]/clk0:18   Xa2s_dout[22]/clk0:19 9.6290 $cpoly
Rg73666 Xa2s_dout[21]/clk0:18   Xa2s_dout[21]/clk0:19 9.6290 $cpoly
Rg73667 Xa2s_dout[20]/clk0:18   Xa2s_dout[20]/clk0:19 9.6290 $cpoly
Rg73668 Xa2s_dout[19]/clk0:18   Xa2s_dout[19]/clk0:19 9.6290 $cpoly
Rg73669 Xa2s_dout[18]/clk0:18   Xa2s_dout[18]/clk0:19 9.6290 $cpoly

Rg73698 Xa2s_dout[22]/_clk:25   Xa2s_dout[22]/_clk:22 126.2881 $cpoly
Rg73699 Xa2s_dout[21]/_clk:25   Xa2s_dout[21]/_clk:22 126.2881 $cpoly
Rg73700 Xa2s_dout[20]/_clk:25   Xa2s_dout[20]/_clk:22 126.2881 $cpoly
Rg73701 Xa2s_dout[19]/_clk:25   Xa2s_dout[19]/_clk:22 126.2881 $cpoly
Rg73702 Xa2s_dout[18]/_clk:25   Xa2s_dout[18]/_clk:22 126.2881 $cpoly

Rg73746 Xa2s_dout[22]/10:1      Xa2s_dout[22]/10:2 11.8495 $cpoly
Rg73747 Xa2s_dout[21]/10:1      Xa2s_dout[21]/10:2 11.8495 $cpoly
Rg73748 Xa2s_dout[20]/10:1      Xa2s_dout[20]/10:2 11.8495 $cpoly
Rg73749 Xa2s_dout[19]/10:1      Xa2s_dout[19]/10:2 11.8495 $cpoly
Rg73750 Xa2s_dout[18]/10:1      Xa2s_dout[18]/10:2 11.8495 $cpoly

Rg73836 Xa2s_dout[21]/_R.0:31   Xa2s_dout[21]/_R.0:32 23.9733 $cpoly
Rg73837 Xa2s_dout[21]/_R.0:31   Xa2s_dout[21]/_R.0:33 16.6712 $cpoly
Rg73838 Xa2s_dout[20]/_R.0:30   Xa2s_dout[20]/_R.0:31 23.9733 $cpoly
Rg73839 Xa2s_dout[20]/_R.0:31   Xa2s_dout[20]/_R.0:32 23.9733 $cpoly
Rg73840 Xa2s_dout[20]/_R.0:31   Xa2s_dout[20]/_R.0:33 16.6712 $cpoly
Rg73841 Xa2s_dout[19]/_R.0:30   Xa2s_dout[19]/_R.0:31 23.9733 $cpoly
Rg73842 Xa2s_dout[19]/_R.0:31   Xa2s_dout[19]/_R.0:32 23.9733 $cpoly

Rg73932 Xa2s_dout[21]/_clk:28   Xa2s_dout[21]/_clk:24 25.4110 $cpoly
Rg73933 Xa2s_dout[21]/_clk:28   Xa2s_dout[21]/_clk:29 98.0510 $cpoly
Rg73934 Xa2s_dout[20]/_clk:27   Xa2s_dout[20]/_clk:28 87.7177 $cpoly
Rg73935 Xa2s_dout[20]/_clk:28   Xa2s_dout[20]/_clk:24 25.4110 $cpoly
Rg73936 Xa2s_dout[20]/_clk:28   Xa2s_dout[20]/_clk:29 98.0510 $cpoly
Rg73937 Xa2s_dout[19]/_clk:27   Xa2s_dout[19]/_clk:28 87.7177 $cpoly
Rg73938 Xa2s_dout[19]/_clk:28   Xa2s_dout[19]/_clk:24 25.4110 $cpoly

Rg74070 Xa2s_dout[22]/_clk0:39  Xa2s_dout[22]/_clk0:27 102.2235 $cpoly
Rg74071 Xa2s_dout[21]/_clk0:39  Xa2s_dout[21]/_clk0:27 102.2235 $cpoly
Rg74072 Xa2s_dout[20]/_clk0:39  Xa2s_dout[20]/_clk0:27 102.2235 $cpoly
Rg74073 Xa2s_dout[19]/_clk0:39  Xa2s_dout[19]/_clk0:27 102.2235 $cpoly
Rg74074 Xa2s_dout[18]/_clk0:39  Xa2s_dout[18]/_clk0:27 102.2235 $cpoly

Rg74103 Xa2s_dout[22]/_clk0:40  Xa2s_dout[22]/_clk0:25 114.3184 $cpoly
Rg74104 Xa2s_dout[21]/_clk0:40  Xa2s_dout[21]/_clk0:25 114.3184 $cpoly
Rg74105 Xa2s_dout[20]/_clk0:40  Xa2s_dout[20]/_clk0:25 114.3184 $cpoly
Rg74106 Xa2s_dout[19]/_clk0:40  Xa2s_dout[19]/_clk0:25 114.3184 $cpoly
Rg74107 Xa2s_dout[18]/_clk0:40  Xa2s_dout[18]/_clk0:25 114.3184 $cpoly

Rg74221 Xa2s_dout[21]/_clk0:42  Xa2s_dout[21]/_clk0:43 46.9874 $cpoly
Rg74222 Xa2s_dout[21]/_clk0:42  Xa2s_dout[21]/_clk0:26 37.8110 $cpoly
Rg74223 Xa2s_dout[20]/_clk0:41  Xa2s_dout[20]/_clk0:42 100.1176 $cpoly
Rg74224 Xa2s_dout[20]/_clk0:42  Xa2s_dout[20]/_clk0:43 46.9874 $cpoly
Rg74225 Xa2s_dout[20]/_clk0:42  Xa2s_dout[20]/_clk0:26 37.8110 $cpoly
Rg74226 Xa2s_dout[19]/_clk0:41  Xa2s_dout[19]/_clk0:42 100.1176 $cpoly
Rg74227 Xa2s_dout[19]/_clk0:42  Xa2s_dout[19]/_clk0:43 46.9874 $cpoly

Rg74370 Xa2s_dout[21]/_clk:30   Xa2s_dout[21]/_clk:23 262.0851 $cpoly
Rg74371 Xa2s_dout[21]/_clk:23   Xa2s_dout[21]/_clk:31 102.2235 $cpoly
Rg74372 Xa2s_dout[20]/_clk:30   Xa2s_dout[20]/_clk:23 262.0851 $cpoly
Rg74373 Xa2s_dout[20]/_clk:23   Xa2s_dout[20]/_clk:31 102.2235 $cpoly
Rg74374 Xa2s_dout[19]/_clk:30   Xa2s_dout[19]/_clk:23 262.0851 $cpoly
Rg74375 Xa2s_dout[19]/_clk:23   Xa2s_dout[19]/_clk:31 102.2235 $cpoly

Rg74631 Xa2s_dout[21]/_clk0:52  Xa2s_dout[21]/_clk0:44 9.5629 $cpoly
Rg74632 Xa2s_dout[21]/_clk0:54  Xa2s_dout[21]/_clk0:44 19.2322 $cpoly
Rg74633 Xa2s_dout[20]/_clk0:31  Xa2s_dout[20]/_clk0:44 15.1749 $cpoly
Rg74634 Xa2s_dout[20]/_clk0:44  Xa2s_dout[20]/_clk0:45 45.0629 $cpoly
Rg74635 Xa2s_dout[20]/_clk0:45  Xa2s_dout[20]/_clk0:46 37.6190 $cpoly
Rg74636 Xa2s_dout[20]/_clk0:46  Xa2s_dout[20]/_clk0:29 1.3357 $cpoly
Rg74637 Xa2s_dout[20]/_clk0:46  Xa2s_dout[20]/_clk0:47 42.0065 $cpoly
Rg74638 Xa2s_dout[20]/_clk0:47  Xa2s_dout[20]/_clk0:48 45.6733 $cpoly
Rg74639 Xa2s_dout[20]/_clk0:48  Xa2s_dout[20]/_clk0:49 36.3733 $cpoly
Rg74640 Xa2s_dout[20]/_clk0:49  Xa2s_dout[20]/_clk0:50 32.7065 $cpoly
Rg74641 Xa2s_dout[20]/_clk0:50  Xa2s_dout[20]/_clk0:51 28.3190 $cpoly
Rg74642 Xa2s_dout[20]/_clk0:48  Xa2s_dout[20]/_clk0:52 7.9178 $cpoly
Rg74643 Xa2s_dout[20]/_clk0:50  Xa2s_dout[20]/_clk0:53 1.3357 $cpoly
Rg74644 Xa2s_dout[20]/_clk0:51  Xa2s_dout[20]/_clk0:54 16.5308 $cpoly
Rg74645 Xa2s_dout[20]/_clk0:52  Xa2s_dout[20]/_clk0:44 9.5629 $cpoly
Rg74646 Xa2s_dout[20]/_clk0:54  Xa2s_dout[20]/_clk0:44 19.2322 $cpoly
Rg74647 Xa2s_dout[19]/_clk0:31  Xa2s_dout[19]/_clk0:44 15.1749 $cpoly
Rg74648 Xa2s_dout[19]/_clk0:44  Xa2s_dout[19]/_clk0:45 45.0629 $cpoly

Rg74939 Xa2s_dout[22]/_clk0:58  Xa2s_dout[22]/_clk0:59 77.4235 $cpoly
Rg74940 Xa2s_dout[21]/_clk0:58  Xa2s_dout[21]/_clk0:59 77.4235 $cpoly
Rg74941 Xa2s_dout[20]/_clk0:58  Xa2s_dout[20]/_clk0:59 77.4235 $cpoly
Rg74942 Xa2s_dout[19]/_clk0:58  Xa2s_dout[19]/_clk0:59 77.4235 $cpoly
Rg74943 Xa2s_dout[18]/_clk0:58  Xa2s_dout[18]/_clk0:59 77.4235 $cpoly

Rg74971 Xa2s_dout[22]/10:6      Xa2s_dout[22]/10:3 5.8022 $cpoly
Rg74972 Xa2s_dout[21]/10:6      Xa2s_dout[21]/10:3 5.8022 $cpoly
Rg74973 Xa2s_dout[20]/10:6      Xa2s_dout[20]/10:3 5.8022 $cpoly
Rg74974 Xa2s_dout[19]/10:6      Xa2s_dout[19]/10:3 5.8022 $cpoly
Rg74975 Xa2s_dout[18]/10:6      Xa2s_dout[18]/10:3 5.8022 $cpoly

Rg75078 Xa2s_dout[22]/clk0:25   Xa2s_dout[22]/clk0:21 3.4772 $cpoly
Rg75079 Xa2s_dout[21]/clk0:25   Xa2s_dout[21]/clk0:21 3.4772 $cpoly
Rg75080 Xa2s_dout[20]/clk0:25   Xa2s_dout[20]/clk0:21 3.4772 $cpoly
Rg75081 Xa2s_dout[19]/clk0:25   Xa2s_dout[19]/clk0:21 3.4772 $cpoly
Rg75082 Xa2s_dout[18]/clk0:25   Xa2s_dout[18]/clk0:21 3.4772 $cpoly

Rg75165 Xa2s_dout[21]/clk0:31   Xa2s_dout[21]/clk0:32 120.9079 $cpoly
Rg75166 Xa2s_dout[21]/clk0:31   Xa2s_dout[21]/clk0:33 82.1869 $cpoly
Rg75167 Xa2s_dout[20]/clk0:26   Xa2s_dout[20]/clk0:27 29.4207 $cpoly
Rg75168 Xa2s_dout[20]/clk0:27   Xa2s_dout[20]/clk0:28 158.1079 $cpoly
Rg75169 Xa2s_dout[20]/clk0:27   Xa2s_dout[20]/clk0:29 92.5202 $cpoly
Rg75170 Xa2s_dout[20]/clk0:30   Xa2s_dout[20]/clk0:31 39.7540 $cpoly
Rg75171 Xa2s_dout[20]/clk0:31   Xa2s_dout[20]/clk0:32 120.9079 $cpoly
Rg75172 Xa2s_dout[20]/clk0:31   Xa2s_dout[20]/clk0:33 82.1869 $cpoly
Rg75173 Xa2s_dout[19]/clk0:26   Xa2s_dout[19]/clk0:27 29.4207 $cpoly
Rg75174 Xa2s_dout[19]/clk0:27   Xa2s_dout[19]/clk0:28 158.1079 $cpoly

Rg75308 Xa2s_dout[22]/_clk0:62  Xa2s_dout[22]/_clk0:56 57.7240 $cpoly
Rg75309 Xa2s_dout[21]/_clk0:62  Xa2s_dout[21]/_clk0:56 57.7240 $cpoly
Rg75310 Xa2s_dout[20]/_clk0:62  Xa2s_dout[20]/_clk0:56 57.7240 $cpoly
Rg75311 Xa2s_dout[19]/_clk0:62  Xa2s_dout[19]/_clk0:56 57.7240 $cpoly
Rg75312 Xa2s_dout[18]/_clk0:62  Xa2s_dout[18]/_clk0:56 57.7240 $cpoly

Rf69311 Xa2s_dout[21]/_noR:7    Xa2s_dout[21]/_noR:8 0.4340 $mt1
Rf69313 Xa2s_dout[21]/_noR:8    Xa2s_dout[21]/_noR:10 0.4314 $mt1
Rf69315 Xa2s_dout[20]/_noR:7    Xa2s_dout[20]/_noR:8 0.4340 $mt1
Rf69317 Xa2s_dout[20]/_noR:8    Xa2s_dout[20]/_noR:10 0.4314 $mt1
Rf69319 Xa2s_dout[19]/_noR:7    Xa2s_dout[19]/_noR:8 0.4340 $mt1
Rf69321 Xa2s_dout[19]/_noR:8    Xa2s_dout[19]/_noR:10 0.4314 $mt1

Rf69442 Xa2s_dout[21]/7:4       Xa2s_dout[21]/7:5 0.3762 $mt1
Rf69443 Xa2s_dout[21]/7:5       Xa2s_dout[21]/7:2 0.4737 $mt1
Rf69444 Xa2s_dout[20]/7:3       Xa2s_dout[20]/7:4 0.2085 $mt1
Rf69445 Xa2s_dout[20]/7:4       Xa2s_dout[20]/7:5 0.3762 $mt1
Rf69446 Xa2s_dout[20]/7:5       Xa2s_dout[20]/7:2 0.4737 $mt1
Rf69447 Xa2s_dout[19]/7:3       Xa2s_dout[19]/7:4 0.2085 $mt1
Rf69448 Xa2s_dout[19]/7:4       Xa2s_dout[19]/7:5 0.3762 $mt1

Rf70192 Xa2s_dout[21]/Rc:4      Xa2s_dout[21]/Rc:5 0.1076 $mt1
Rf70193 Xa2s_dout[21]/Rc:4      Xa2s_dout[21]/Rc:6 0.2965 $mt1
Rf70196 Xa2s_dout[20]/Rc:1      Xa2s_dout[20]/Rc:4 0.1022 $mt1
Rf70197 Xa2s_dout[20]/Rc:4      Xa2s_dout[20]/Rc:5 0.1076 $mt1
Rf70198 Xa2s_dout[20]/Rc:4      Xa2s_dout[20]/Rc:6 0.2965 $mt1
Rf70201 Xa2s_dout[19]/Rc:1      Xa2s_dout[19]/Rc:4 0.1022 $mt1
Rf70202 Xa2s_dout[19]/Rc:4      Xa2s_dout[19]/Rc:5 0.1076 $mt1

Rf70331 Xa2s_dout[21]/6:4       Xa2s_dout[21]/6:5 0.3762 $mt1
Rf70332 Xa2s_dout[21]/6:5       Xa2s_dout[21]/6:2 0.4347 $mt1
Rf70333 Xa2s_dout[20]/6:3       Xa2s_dout[20]/6:4 0.4347 $mt1
Rf70334 Xa2s_dout[20]/6:4       Xa2s_dout[20]/6:5 0.3762 $mt1
Rf70335 Xa2s_dout[20]/6:5       Xa2s_dout[20]/6:2 0.4347 $mt1
Rf70336 Xa2s_dout[19]/6:3       Xa2s_dout[19]/6:4 0.4347 $mt1
Rf70337 Xa2s_dout[19]/6:4       Xa2s_dout[19]/6:5 0.3762 $mt1

Rf70458 Xa2s_dout[22]/_Le:1     Xa2s_dout[22]/_Le:6 0.2607 $mt1
Rf70461 Xa2s_dout[21]/_Le:1     Xa2s_dout[21]/_Le:6 0.2607 $mt1
Rf70464 Xa2s_dout[20]/_Le:1     Xa2s_dout[20]/_Le:6 0.2607 $mt1
Rf70467 Xa2s_dout[19]/_Le:1     Xa2s_dout[19]/_Le:6 0.2607 $mt1
Rf70470 Xa2s_dout[18]/_Le:1     Xa2s_dout[18]/_Le:6 0.2607 $mt1

Rf70753 Xa2s_dout[21]/_R.0:9    Xa2s_dout[21]/_R.0:11 2.2244 $mt1
Rf70754 Xa2s_dout[21]/_R.0:11   Xa2s_dout[21]/_R.0:12 1.3074 $mt1
Rf70757 Xa2s_dout[20]/_R.0:9    Xa2s_dout[20]/_R.0:11 2.2244 $mt1
Rf70758 Xa2s_dout[20]/_R.0:11   Xa2s_dout[20]/_R.0:12 1.3074 $mt1
Rf70761 Xa2s_dout[19]/_R.0:9    Xa2s_dout[19]/_R.0:11 2.2244 $mt1
Rf70762 Xa2s_dout[19]/_R.0:11   Xa2s_dout[19]/_R.0:12 1.3074 $mt1

Rf70925 Xa2s_dout[21]/_R.1:7    Xa2s_dout[21]/_R.1:10 0.1690 $mt1
Rf70926 Xa2s_dout[21]/_R.1:21   Xa2s_dout[21]/_R.1:13 0.1635 $mt1
Rf70928 Xa2s_dout[20]/_R.1:18   Xa2s_dout[20]/_R.1:19 0.2307 $mt1
Rf70929 Xa2s_dout[20]/_R.1:19   Xa2s_dout[20]/_R.1:21 0.1478 $mt1
Rf70930 Xa2s_dout[20]/_R.1:21   Xa2s_dout[20]/_R.1:1 0.7417 $mt1
Rf70931 Xa2s_dout[20]/_R.1:1    Xa2s_dout[20]/_R.1:4 0.1690 $mt1
Rf70932 Xa2s_dout[20]/_R.1:4    Xa2s_dout[20]/_R.1:7 0.1690 $mt1
Rf70933 Xa2s_dout[20]/_R.1:7    Xa2s_dout[20]/_R.1:10 0.1690 $mt1
Rf70934 Xa2s_dout[20]/_R.1:21   Xa2s_dout[20]/_R.1:13 0.1635 $mt1
Rf70936 Xa2s_dout[19]/_R.1:18   Xa2s_dout[19]/_R.1:19 0.2307 $mt1
Rf70937 Xa2s_dout[19]/_R.1:19   Xa2s_dout[19]/_R.1:21 0.1478 $mt1

Rf71668 Xa2s_dout[22]/_R.1:24   Xa2s_dout[22]/_R.1:15 0.5492 $mt1
Rf71671 Xa2s_dout[21]/_R.1:24   Xa2s_dout[21]/_R.1:15 0.5492 $mt1
Rf71674 Xa2s_dout[20]/_R.1:24   Xa2s_dout[20]/_R.1:15 0.5492 $mt1
Rf71677 Xa2s_dout[19]/_R.1:24   Xa2s_dout[19]/_R.1:15 0.5492 $mt1
Rf71680 Xa2s_dout[18]/_R.1:24   Xa2s_dout[18]/_R.1:15 0.5492 $mt1

Rf71832 Xa2s_dout[21]/_r:12     Xa2s_dout[21]/_r:6 0.1690 $mt1
Rf71833 Xa2s_dout[21]/_r:6      Xa2s_dout[21]/_r:3 0.2177 $mt1
Rf71834 Xa2s_dout[20]/_r:13     Xa2s_dout[20]/_r:16 0.2973 $mt1
Rf71837 Xa2s_dout[20]/_r:16     Xa2s_dout[20]/_r:17 2.1775 $mt1
Rf71838 Xa2s_dout[20]/_r:17     Xa2s_dout[20]/_r:18 0.3132 $mt1
Rf71839 Xa2s_dout[20]/_r:16     Xa2s_dout[20]/_r:9 0.4241 $mt1
Rf71840 Xa2s_dout[20]/_r:9      Xa2s_dout[20]/_r:12 0.2177 $mt1
Rf71841 Xa2s_dout[20]/_r:12     Xa2s_dout[20]/_r:6 0.1690 $mt1
Rf71842 Xa2s_dout[20]/_r:6      Xa2s_dout[20]/_r:3 0.2177 $mt1
Rf71843 Xa2s_dout[19]/_r:13     Xa2s_dout[19]/_r:16 0.2973 $mt1
Rf71846 Xa2s_dout[19]/_r:16     Xa2s_dout[19]/_r:17 2.1775 $mt1

Rf73534 Xa2s_dout[21]/_noR:20   Xa2s_dout[21]/_noR:21 0.7188 $mt1
Rf73535 Xa2s_dout[21]/_noR:20   Xa2s_dout[21]/_noR:22 0.1939 $mt1
Rf73539 Xa2s_dout[20]/_noR:17   Xa2s_dout[20]/_noR:17 0.6368 $mt1
Rf73540 Xa2s_dout[20]/_noR:17   Xa2s_dout[20]/_noR:14 1.3013 $mt1
Rf73541 Xa2s_dout[20]/_noR:14   Xa2s_dout[20]/_noR:20 2.3675 $mt1
Rf73542 Xa2s_dout[20]/_noR:20   Xa2s_dout[20]/_noR:21 0.7188 $mt1
Rf73543 Xa2s_dout[20]/_noR:20   Xa2s_dout[20]/_noR:22 0.1939 $mt1
Rf73547 Xa2s_dout[19]/_noR:17   Xa2s_dout[19]/_noR:17 0.6368 $mt1
Rf73548 Xa2s_dout[19]/_noR:17   Xa2s_dout[19]/_noR:14 1.3013 $mt1

Rf73840 Xa2s_dout[21]/__Le:10   Xa2s_dout[21]/__Le:7 0.5883 $mt1
Rf73841 Xa2s_dout[21]/__Le:7    Xa2s_dout[21]/__Le:11 3.6046 $mt1
Rf73842 Xa2s_dout[20]/__Le:4    Xa2s_dout[20]/__Le:8 0.3848 $mt1
Rf73843 Xa2s_dout[20]/__Le:8    Xa2s_dout[20]/__Le:9 0.4545 $mt1
Rf73844 Xa2s_dout[20]/__Le:4    Xa2s_dout[20]/__Le:10 0.5752 $mt1
Rf73845 Xa2s_dout[20]/__Le:10   Xa2s_dout[20]/__Le:7 0.5883 $mt1
Rf73846 Xa2s_dout[20]/__Le:7    Xa2s_dout[20]/__Le:11 3.6046 $mt1
Rf73847 Xa2s_dout[19]/__Le:4    Xa2s_dout[19]/__Le:8 0.3848 $mt1
Rf73848 Xa2s_dout[19]/__Le:8    Xa2s_dout[19]/__Le:9 0.4545 $mt1

Rf74028 Xa2s_dout[22]/51:1      Xa2s_dout[22]/51:2 0.6861 $mt1
Rf74029 Xa2s_dout[21]/51:1      Xa2s_dout[21]/51:2 0.6861 $mt1
Rf74030 Xa2s_dout[20]/51:1      Xa2s_dout[20]/51:2 0.6861 $mt1
Rf74031 Xa2s_dout[19]/51:1      Xa2s_dout[19]/51:2 0.6861 $mt1
Rf74032 Xa2s_dout[18]/51:1      Xa2s_dout[18]/51:2 0.6861 $mt1

Rf74100 Xa2s_dout[21]/clk0:6    Xa2s_dout[21]/clk0:3 0.2870 $mt1
Rf74101 Xa2s_dout[21]/clk0:6    Xa2s_dout[21]/clk0:1 0.5730 $mt1
Rf74102 Xa2s_dout[20]/clk0:5    Xa2s_dout[20]/clk0:6 0.7848 $mt1
Rf74103 Xa2s_dout[20]/clk0:6    Xa2s_dout[20]/clk0:3 0.2870 $mt1
Rf74104 Xa2s_dout[20]/clk0:6    Xa2s_dout[20]/clk0:1 0.5730 $mt1
Rf74105 Xa2s_dout[19]/clk0:5    Xa2s_dout[19]/clk0:6 0.7848 $mt1
Rf74106 Xa2s_dout[19]/clk0:6    Xa2s_dout[19]/clk0:3 0.2870 $mt1

Rf74313 Xa2s_dout[22]/clk0:9    Xa2s_dout[22]/clk0:10 0.3978 $mt1
Rf74314 Xa2s_dout[21]/clk0:9    Xa2s_dout[21]/clk0:10 0.3978 $mt1
Rf74315 Xa2s_dout[20]/clk0:9    Xa2s_dout[20]/clk0:10 0.3978 $mt1
Rf74316 Xa2s_dout[19]/clk0:9    Xa2s_dout[19]/clk0:10 0.3978 $mt1
Rf74317 Xa2s_dout[18]/clk0:9    Xa2s_dout[18]/clk0:10 0.3978 $mt1

Rf74387 Xa2s_dout[22]/_clk:9    Xa2s_dout[22]/_clk:11 0.9508 $mt1
Rf74392 Xa2s_dout[21]/_clk:9    Xa2s_dout[21]/_clk:11 0.9508 $mt1
Rf74397 Xa2s_dout[20]/_clk:9    Xa2s_dout[20]/_clk:11 0.9508 $mt1
Rf74402 Xa2s_dout[19]/_clk:9    Xa2s_dout[19]/_clk:11 0.9508 $mt1
Rf74407 Xa2s_dout[18]/_clk:9    Xa2s_dout[18]/_clk:11 0.9508 $mt1

Rf75207 Xa2s_dout[22]/29:1      Xa2s_dout[22]/29:2 1.2321 $mt1
Rf75210 Xa2s_dout[21]/29:1      Xa2s_dout[21]/29:2 1.2321 $mt1
Rf75213 Xa2s_dout[20]/29:1      Xa2s_dout[20]/29:2 1.2321 $mt1
Rf75216 Xa2s_dout[19]/29:1      Xa2s_dout[19]/29:2 1.2321 $mt1
Rf75219 Xa2s_dout[18]/29:1      Xa2s_dout[18]/29:2 1.2321 $mt1

Rf75675 Xa2s_dout[22]/26:1      Xa2s_dout[22]/26:2 1.3169 $mt1
Rf75676 Xa2s_dout[21]/26:1      Xa2s_dout[21]/26:2 1.3169 $mt1
Rf75677 Xa2s_dout[20]/26:1      Xa2s_dout[20]/26:2 1.3169 $mt1
Rf75678 Xa2s_dout[19]/26:1      Xa2s_dout[19]/26:2 1.3169 $mt1
Rf75679 Xa2s_dout[18]/26:1      Xa2s_dout[18]/26:2 1.3169 $mt1

Rf75750 Xa2s_dout[21]/PReset:9  Xa2s_dout[21]/PReset:10 0.2095 $mt1
Rf75751 Xa2s_dout[21]/PReset:10 Xa2s_dout[21]/PReset:4 0.1061 $mt1
Rf75752 Xa2s_dout[20]/PReset:9  Xa2s_dout[20]/PReset:10 0.2095 $mt1
Rf75753 Xa2s_dout[20]/PReset:10 Xa2s_dout[20]/PReset:4 0.1061 $mt1
Rf75754 Xa2s_dout[19]/PReset:9  Xa2s_dout[19]/PReset:10 0.2095 $mt1
Rf75755 Xa2s_dout[19]/PReset:10 Xa2s_dout[19]/PReset:4 0.1061 $mt1

Rf75806 Xa2s_dout[22]/31:1      Xa2s_dout[22]/31:2 1.4141 $mt1
Rf75807 Xa2s_dout[21]/31:1      Xa2s_dout[21]/31:2 1.4141 $mt1
Rf75808 Xa2s_dout[20]/31:1      Xa2s_dout[20]/31:2 1.4141 $mt1
Rf75809 Xa2s_dout[19]/31:1      Xa2s_dout[19]/31:2 1.4141 $mt1
Rf75810 Xa2s_dout[18]/31:1      Xa2s_dout[18]/31:2 1.4141 $mt1

Rf75916 Xa2s_dout[21]/Rv:12     Xa2s_dout[21]/Rv:14 0.6672 $mt1
Rf75917 Xa2s_dout[21]/Rv:2      Xa2s_dout[21]/Rv:4 6.2065 $mt1
Rf75918 Xa2s_dout[20]/Rv:9      Xa2s_dout[20]/Rv:8 0.4347 $mt1
Rf75919 Xa2s_dout[20]/Rv:8      Xa2s_dout[20]/Rv:10 0.4347 $mt1
Rf75920 Xa2s_dout[20]/Rv:10     Xa2s_dout[20]/Rv:11 2.9365 $mt1
Rf75921 Xa2s_dout[20]/Rv:11     Xa2s_dout[20]/Rv:12 0.1873 $mt1
Rf75922 Xa2s_dout[20]/Rv:12     Xa2s_dout[20]/Rv:13 1.5003 $mt1
Rf75923 Xa2s_dout[20]/Rv:13     Xa2s_dout[20]/Rv:2 4.6075 $mt1
Rf75924 Xa2s_dout[20]/Rv:12     Xa2s_dout[20]/Rv:14 0.6672 $mt1
Rf75925 Xa2s_dout[20]/Rv:2      Xa2s_dout[20]/Rv:4 6.2065 $mt1
Rf75926 Xa2s_dout[19]/Rv:9      Xa2s_dout[19]/Rv:8 0.4347 $mt1
Rf75927 Xa2s_dout[19]/Rv:8      Xa2s_dout[19]/Rv:10 0.4347 $mt1

Rf76131 Xa2s_dout[21]/8:4       Xa2s_dout[21]/8:5 0.3762 $mt1
Rf76132 Xa2s_dout[21]/8:5       Xa2s_dout[21]/8:2 0.4737 $mt1
Rf76133 Xa2s_dout[20]/8:3       Xa2s_dout[20]/8:4 0.2085 $mt1
Rf76134 Xa2s_dout[20]/8:4       Xa2s_dout[20]/8:5 0.3762 $mt1
Rf76135 Xa2s_dout[20]/8:5       Xa2s_dout[20]/8:2 0.4737 $mt1
Rf76136 Xa2s_dout[19]/8:3       Xa2s_dout[19]/8:4 0.2085 $mt1
Rf76137 Xa2s_dout[19]/8:4       Xa2s_dout[19]/8:5 0.3762 $mt1

Rf76322 Xa2s_dout[21]/Rc:9      Xa2s_dout[21]/Rc:10 0.5492 $mt1
Rf76323 Xa2s_dout[21]/Rc:10     Xa2s_dout[21]/Rc:7 0.4498 $mt1
Rf76325 Xa2s_dout[20]/Rc:9      Xa2s_dout[20]/Rc:10 0.5492 $mt1
Rf76326 Xa2s_dout[20]/Rc:10     Xa2s_dout[20]/Rc:7 0.4498 $mt1
Rf76328 Xa2s_dout[19]/Rc:9      Xa2s_dout[19]/Rc:10 0.5492 $mt1
Rf76329 Xa2s_dout[19]/Rc:10     Xa2s_dout[19]/Rc:7 0.4498 $mt1

Rf76603 Xa2s_dout[21]/_clk0:20  Xa2s_dout[21]/_clk0:12 0.8961 $mt1
Rf76604 Xa2s_dout[21]/_clk0:21  Xa2s_dout[21]/_clk0:7 1.1677 $mt1
Rf76606 Xa2s_dout[20]/_clk0:17  Xa2s_dout[20]/_clk0:15 0.5473 $mt1
Rf76607 Xa2s_dout[20]/_clk0:15  Xa2s_dout[20]/_clk0:18 0.4570 $mt1
Rf76608 Xa2s_dout[20]/_clk0:18  Xa2s_dout[20]/_clk0:19 0.1077 $mt1
Rf76609 Xa2s_dout[20]/_clk0:19  Xa2s_dout[20]/_clk0:20 0.5341 $mt1
Rf76610 Xa2s_dout[20]/_clk0:20  Xa2s_dout[20]/_clk0:14 1.0550 $mt1
Rf76611 Xa2s_dout[20]/_clk0:14  Xa2s_dout[20]/_clk0:21 0.7027 $mt1
Rf76612 Xa2s_dout[20]/_clk0:21  Xa2s_dout[20]/_clk0:1 0.4022 $mt1
Rf76614 Xa2s_dout[20]/_clk0:19  Xa2s_dout[20]/_clk0:24 0.5565 $mt1
Rf76615 Xa2s_dout[20]/_clk0:20  Xa2s_dout[20]/_clk0:12 0.8961 $mt1
Rf76616 Xa2s_dout[20]/_clk0:21  Xa2s_dout[20]/_clk0:7 1.1677 $mt1
Rf76618 Xa2s_dout[19]/_clk0:17  Xa2s_dout[19]/_clk0:15 0.5473 $mt1
Rf76619 Xa2s_dout[19]/_clk0:15  Xa2s_dout[19]/_clk0:18 0.4570 $mt1

Rf76915 Xa2s_dout[21]/9:4       Xa2s_dout[21]/9:5 0.3762 $mt1
Rf76916 Xa2s_dout[21]/9:5       Xa2s_dout[21]/9:2 0.4347 $mt1
Rf76917 Xa2s_dout[20]/9:3       Xa2s_dout[20]/9:4 0.4347 $mt1
Rf76918 Xa2s_dout[20]/9:4       Xa2s_dout[20]/9:5 0.3762 $mt1
Rf76919 Xa2s_dout[20]/9:5       Xa2s_dout[20]/9:2 0.4347 $mt1
Rf76920 Xa2s_dout[19]/9:3       Xa2s_dout[19]/9:4 0.4347 $mt1
Rf76921 Xa2s_dout[19]/9:4       Xa2s_dout[19]/9:5 0.3762 $mt1

Rf77063 Xa2s_dout[21]/_R.1:43   Xa2s_dout[21]/_R.1:32 0.4496 $mt1
Rf77065 Xa2s_dout[21]/_R.1:32   Xa2s_dout[21]/_R.1:30 0.1462 $mt1
Rf77069 Xa2s_dout[20]/_R.1:41   Xa2s_dout[20]/_R.1:39 0.5785 $mt1
Rf77070 Xa2s_dout[20]/_R.1:39   Xa2s_dout[20]/_R.1:43 0.3848 $mt1
Rf77071 Xa2s_dout[20]/_R.1:43   Xa2s_dout[20]/_R.1:32 0.4496 $mt1
Rf77073 Xa2s_dout[20]/_R.1:32   Xa2s_dout[20]/_R.1:30 0.1462 $mt1
Rf77077 Xa2s_dout[19]/_R.1:41   Xa2s_dout[19]/_R.1:39 0.5785 $mt1
Rf77078 Xa2s_dout[19]/_R.1:39   Xa2s_dout[19]/_R.1:43 0.3848 $mt1

Rf77484 Xa2s_dout[22]/_grant:1  Xa2s_dout[22]/_grant:2 0.4582 $mt1
Rf77485 Xa2s_dout[21]/_grant:1  Xa2s_dout[21]/_grant:2 0.4582 $mt1
Rf77486 Xa2s_dout[20]/_grant:1  Xa2s_dout[20]/_grant:2 0.4582 $mt1
Rf77487 Xa2s_dout[19]/_grant:1  Xa2s_dout[19]/_grant:2 0.4582 $mt1
Rf77488 Xa2s_dout[18]/_grant:1  Xa2s_dout[18]/_grant:2 0.4582 $mt1

Rf77547 Xa2s_dout[22]/clk0:15   Xa2s_dout[22]/clk0:17 0.9847 $mt1
Rf77548 Xa2s_dout[21]/clk0:15   Xa2s_dout[21]/clk0:17 0.9847 $mt1
Rf77549 Xa2s_dout[20]/clk0:15   Xa2s_dout[20]/clk0:17 0.9847 $mt1
Rf77550 Xa2s_dout[19]/clk0:15   Xa2s_dout[19]/clk0:17 0.9847 $mt1
Rf77551 Xa2s_dout[18]/clk0:15   Xa2s_dout[18]/clk0:17 0.9847 $mt1

Rf77777 Xa2s_dout[22]/_clk0:25  Xa2s_dout[22]/_clk0:26 1.1820 $mt1
Rf77778 Xa2s_dout[21]/_clk0:25  Xa2s_dout[21]/_clk0:26 1.1820 $mt1
Rf77779 Xa2s_dout[20]/_clk0:25  Xa2s_dout[20]/_clk0:26 1.1820 $mt1
Rf77780 Xa2s_dout[19]/_clk0:25  Xa2s_dout[19]/_clk0:26 1.1820 $mt1
Rf77781 Xa2s_dout[18]/_clk0:25  Xa2s_dout[18]/_clk0:26 1.1820 $mt1

Rf77831 Xa2s_dout[21]/_clk:24   Xa2s_dout[21]/_clk:25 0.1182 $mt1
Rf77832 Xa2s_dout[21]/_clk:25   Xa2s_dout[21]/_clk:19 0.1778 $mt1
Rf77833 Xa2s_dout[20]/_clk:23   Xa2s_dout[20]/_clk:24 0.9499 $mt1
Rf77834 Xa2s_dout[20]/_clk:24   Xa2s_dout[20]/_clk:25 0.1182 $mt1
Rf77835 Xa2s_dout[20]/_clk:25   Xa2s_dout[20]/_clk:19 0.1778 $mt1
Rf77836 Xa2s_dout[19]/_clk:23   Xa2s_dout[19]/_clk:24 0.9499 $mt1
Rf77837 Xa2s_dout[19]/_clk:24   Xa2s_dout[19]/_clk:25 0.1182 $mt1

Rf77974 Xa2s_dout[22]/_clk0:29  Xa2s_dout[22]/_clk0:30 0.1171 $mt1
Rf77975 Xa2s_dout[21]/_clk0:29  Xa2s_dout[21]/_clk0:30 0.1171 $mt1
Rf77976 Xa2s_dout[20]/_clk0:29  Xa2s_dout[20]/_clk0:30 0.1171 $mt1
Rf77977 Xa2s_dout[19]/_clk0:29  Xa2s_dout[19]/_clk0:30 0.1171 $mt1
Rf77978 Xa2s_dout[18]/_clk0:29  Xa2s_dout[18]/_clk0:30 0.1171 $mt1

Rf78366 Xa2s_dout[22]/_R.0:29   Xa2s_dout[22]/_R.0:28 0.1311 $mt1
Rf78373 Xa2s_dout[21]/_R.0:29   Xa2s_dout[21]/_R.0:28 0.1311 $mt1
Rf78380 Xa2s_dout[20]/_R.0:29   Xa2s_dout[20]/_R.0:28 0.1311 $mt1
Rf78387 Xa2s_dout[19]/_R.0:29   Xa2s_dout[19]/_R.0:28 0.1311 $mt1
Rf78394 Xa2s_dout[18]/_R.0:29   Xa2s_dout[18]/_R.0:28 0.1311 $mt1

Rf78789 Xa2s_dout[22]/_grant:7  Xa2s_dout[22]/_grant:6 0.2126 $mt1
Rf78792 Xa2s_dout[21]/_grant:7  Xa2s_dout[21]/_grant:6 0.2126 $mt1
Rf78795 Xa2s_dout[20]/_grant:7  Xa2s_dout[20]/_grant:6 0.2126 $mt1
Rf78798 Xa2s_dout[19]/_grant:7  Xa2s_dout[19]/_grant:6 0.2126 $mt1
Rf78801 Xa2s_dout[18]/_grant:7  Xa2s_dout[18]/_grant:6 0.2126 $mt1

Rf78896 Xa2s_dout[21]/10:4      Xa2s_dout[21]/10:5 0.3762 $mt1
Rf78897 Xa2s_dout[21]/10:5      Xa2s_dout[21]/10:2 0.4737 $mt1
Rf78898 Xa2s_dout[20]/10:3      Xa2s_dout[20]/10:4 0.2085 $mt1
Rf78899 Xa2s_dout[20]/10:4      Xa2s_dout[20]/10:5 0.3762 $mt1
Rf78900 Xa2s_dout[20]/10:5      Xa2s_dout[20]/10:2 0.4737 $mt1
Rf78901 Xa2s_dout[19]/10:3      Xa2s_dout[19]/10:4 0.2085 $mt1
Rf78902 Xa2s_dout[19]/10:4      Xa2s_dout[19]/10:5 0.3762 $mt1

Rf79015 Xa2s_dout[21]/_clk:32   Xa2s_dout[21]/_clk:33 0.1969 $mt1
Rf79016 Xa2s_dout[21]/_clk:33   Xa2s_dout[21]/_clk:22 1.0948 $mt1
Rf79019 Xa2s_dout[20]/_clk:32   Xa2s_dout[20]/_clk:33 0.1969 $mt1
Rf79020 Xa2s_dout[20]/_clk:33   Xa2s_dout[20]/_clk:22 1.0948 $mt1
Rf79023 Xa2s_dout[19]/_clk:32   Xa2s_dout[19]/_clk:33 0.1969 $mt1
Rf79024 Xa2s_dout[19]/_clk:33   Xa2s_dout[19]/_clk:22 1.0948 $mt1

Rf79144 Xa2s_dout[21]/_clk0:56  Xa2s_dout[21]/_clk0:58 0.1119 $mt1
Rf79145 Xa2s_dout[21]/_clk0:58  Xa2s_dout[21]/_clk0:35 0.8073 $mt1
Rf79148 Xa2s_dout[20]/_clk0:56  Xa2s_dout[20]/_clk0:58 0.1119 $mt1
Rf79149 Xa2s_dout[20]/_clk0:58  Xa2s_dout[20]/_clk0:35 0.8073 $mt1
Rf79152 Xa2s_dout[19]/_clk0:56  Xa2s_dout[19]/_clk0:58 0.1119 $mt1
Rf79153 Xa2s_dout[19]/_clk0:58  Xa2s_dout[19]/_clk0:35 0.8073 $mt1

Rf79285 Xa2s_dout[21]/_R.0:33   Xa2s_dout[21]/_R.0:35 0.3848 $mt1
Rf79286 Xa2s_dout[21]/_R.0:35   Xa2s_dout[21]/_R.0:25 0.4503 $mt1
Rf79289 Xa2s_dout[20]/_R.0:34   Xa2s_dout[20]/_R.0:33 0.5720 $mt1
Rf79290 Xa2s_dout[20]/_R.0:33   Xa2s_dout[20]/_R.0:35 0.3848 $mt1
Rf79291 Xa2s_dout[20]/_R.0:35   Xa2s_dout[20]/_R.0:25 0.4503 $mt1
Rf79294 Xa2s_dout[19]/_R.0:34   Xa2s_dout[19]/_R.0:33 0.5720 $mt1
Rf79295 Xa2s_dout[19]/_R.0:33   Xa2s_dout[19]/_R.0:35 0.3848 $mt1

Rf79449 Xa2s_dout[21]/clk0:23   Xa2s_dout[21]/clk0:24 0.2364 $mt1
Rf79450 Xa2s_dout[21]/clk0:24   Xa2s_dout[21]/clk0:18 0.1876 $mt1
Rf79453 Xa2s_dout[20]/clk0:21   Xa2s_dout[20]/clk0:23 0.1768 $mt1
Rf79454 Xa2s_dout[20]/clk0:23   Xa2s_dout[20]/clk0:24 0.2364 $mt1
Rf79455 Xa2s_dout[20]/clk0:24   Xa2s_dout[20]/clk0:18 0.1876 $mt1
Rf79458 Xa2s_dout[19]/clk0:21   Xa2s_dout[19]/clk0:23 0.1768 $mt1
Rf79459 Xa2s_dout[19]/clk0:23   Xa2s_dout[19]/clk0:24 0.2364 $mt1

Rf79570 Xa2s_dout[22]/_clk0:60  Xa2s_dout[22]/_clk0:53 0.1617 $mt1
Rf79571 Xa2s_dout[21]/_clk0:60  Xa2s_dout[21]/_clk0:53 0.1617 $mt1
Rf79572 Xa2s_dout[20]/_clk0:60  Xa2s_dout[20]/_clk0:53 0.1617 $mt1
Rf79573 Xa2s_dout[19]/_clk0:60  Xa2s_dout[19]/_clk0:53 0.1617 $mt1
Rf79574 Xa2s_dout[18]/_clk0:60  Xa2s_dout[18]/_clk0:53 0.1617 $mt1

Rf79613 Xa2s_dout[21]/clk0:26   Xa2s_dout[21]/clk0:30 1.3269 $mt1
Rf79614 Xa2s_dout[21]/clk0:30   Xa2s_dout[21]/clk0:34 0.9912 $mt1
Rf79615 Xa2s_dout[20]/clk0:26   Xa2s_dout[20]/clk0:30 1.3269 $mt1
Rf79616 Xa2s_dout[20]/clk0:30   Xa2s_dout[20]/clk0:34 0.9912 $mt1
Rf79617 Xa2s_dout[19]/clk0:26   Xa2s_dout[19]/clk0:30 1.3269 $mt1
Rf79618 Xa2s_dout[19]/clk0:30   Xa2s_dout[19]/clk0:34 0.9912 $mt1

Rf79796 Xa2s_dout[22]/_clk0:62  Xa2s_dout[22]/_clk0:43 4.6008 $mt1
Rf79799 Xa2s_dout[21]/_clk0:62  Xa2s_dout[21]/_clk0:43 4.6008 $mt1
Rf79802 Xa2s_dout[20]/_clk0:62  Xa2s_dout[20]/_clk0:43 4.6008 $mt1
Rf79805 Xa2s_dout[19]/_clk0:62  Xa2s_dout[19]/_clk0:43 4.6008 $mt1
Rf79808 Xa2s_dout[18]/_clk0:62  Xa2s_dout[18]/_clk0:43 4.6008 $mt1

Re28384 Xa2s_dout[22]/_Le:1     Xa2s_dout[22]/_Le:2 6.4000 $mt2
Re28385 Xa2s_dout[21]/_Le:1     Xa2s_dout[21]/_Le:2 6.4000 $mt2
Re28386 Xa2s_dout[20]/_Le:1     Xa2s_dout[20]/_Le:2 6.4000 $mt2
Re28387 Xa2s_dout[19]/_Le:1     Xa2s_dout[19]/_Le:2 6.4000 $mt2
Re28388 Xa2s_dout[18]/_Le:1     Xa2s_dout[18]/_Le:2 6.4000 $mt2

Re28422 Xa2s_dout[22]/_R.0:4    Xa2s_dout[22]/_R.0:5 6.4000 $mt2
Re28423 Xa2s_dout[21]/_R.0:4    Xa2s_dout[21]/_R.0:5 6.4000 $mt2
Re28424 Xa2s_dout[20]/_R.0:4    Xa2s_dout[20]/_R.0:5 6.4000 $mt2
Re28425 Xa2s_dout[19]/_R.0:4    Xa2s_dout[19]/_R.0:5 6.4000 $mt2
Re28426 Xa2s_dout[18]/_R.0:4    Xa2s_dout[18]/_R.0:5 6.4000 $mt2

Re28797 Xa2s_dout[21]/_R.1:25   Xa2s_dout[21]/_R.1:22 6.4000 $mt2
Re28798 Xa2s_dout[21]/_R.1:24   Xa2s_dout[21]/_R.1:26 6.4000 $mt2
Re28799 Xa2s_dout[20]/_R.1:25   Xa2s_dout[20]/_R.1:22 6.4000 $mt2
Re28800 Xa2s_dout[20]/_R.1:24   Xa2s_dout[20]/_R.1:26 6.4000 $mt2
Re28801 Xa2s_dout[19]/_R.1:25   Xa2s_dout[19]/_R.1:22 6.4000 $mt2
Re28802 Xa2s_dout[19]/_R.1:24   Xa2s_dout[19]/_R.1:26 6.4000 $mt2

Re28876 Xa2s_dout[21]/_noR:15   Xa2s_dout[21]/_noR:1 6.6915 $mt2
Re28877 Xa2s_dout[21]/_noR:8    Xa2s_dout[21]/_noR:15 6.4000 $mt2
Re28878 Xa2s_dout[20]/_noR:14   Xa2s_dout[20]/_noR:15 7.7933 $mt2
Re28879 Xa2s_dout[20]/_noR:15   Xa2s_dout[20]/_noR:1 6.6915 $mt2
Re28880 Xa2s_dout[20]/_noR:8    Xa2s_dout[20]/_noR:15 6.4000 $mt2
Re28881 Xa2s_dout[19]/_noR:14   Xa2s_dout[19]/_noR:15 7.7933 $mt2
Re28882 Xa2s_dout[19]/_noR:15   Xa2s_dout[19]/_noR:1 6.6915 $mt2

Re29085 Xa2s_dout[21]/1:3       Xa2s_dout[21]/1:4 6.6785 $mt2
Re29086 Xa2s_dout[21]/1:2       Xa2s_dout[21]/1:3 6.4000 $mt2
Re29087 Xa2s_dout[20]/1:1       Xa2s_dout[20]/1:3 7.0100 $mt2
Re29088 Xa2s_dout[20]/1:3       Xa2s_dout[20]/1:4 6.6785 $mt2
Re29089 Xa2s_dout[20]/1:2       Xa2s_dout[20]/1:3 6.4000 $mt2
Re29090 Xa2s_dout[19]/1:1       Xa2s_dout[19]/1:3 7.0100 $mt2
Re29091 Xa2s_dout[19]/1:3       Xa2s_dout[19]/1:4 6.6785 $mt2

Re29595 Xa2s_dout[21]/0:1       Xa2s_dout[21]/0:5 6.6767 $mt2
Re29597 Xa2s_dout[21]/0:3       Xa2s_dout[21]/0:1 6.4000 $mt2
Re29598 Xa2s_dout[20]/_clk0:1   Xa2s_dout[20]/_clk0:3 6.6785 $mt2
Re29599 Xa2s_dout[20]/_clk0:3   Xa2s_dout[20]/_clk0:4 6.6785 $mt2
Re29600 Xa2s_dout[20]/_clk0:2   Xa2s_dout[20]/_clk0:3 6.4000 $mt2
Re29602 Xa2s_dout[20]/0:1       Xa2s_dout[20]/0:5 6.6767 $mt2
Re29604 Xa2s_dout[20]/0:3       Xa2s_dout[20]/0:1 6.4000 $mt2
Re29605 Xa2s_dout[19]/_clk0:1   Xa2s_dout[19]/_clk0:3 6.6785 $mt2
Re29606 Xa2s_dout[19]/_clk0:3   Xa2s_dout[19]/_clk0:4 6.6785 $mt2

Re29754 Xa2s_dout[22]/0:6       Xa2s_dout[22]/0:7 6.4000 $mt2
Re29755 Xa2s_dout[21]/0:6       Xa2s_dout[21]/0:7 6.4000 $mt2
Re29756 Xa2s_dout[20]/0:6       Xa2s_dout[20]/0:7 6.4000 $mt2
Re29757 Xa2s_dout[19]/0:6       Xa2s_dout[19]/0:7 6.4000 $mt2
Re29758 Xa2s_dout[18]/0:6       Xa2s_dout[18]/0:7 6.4000 $mt2

Re29845 Xa2s_dout[21]/_R.0:16   Xa2s_dout[21]/_R.0:1 7.1075 $mt2
Re29846 Xa2s_dout[21]/_R.0:9    Xa2s_dout[21]/_R.0:16 6.4000 $mt2
Re29847 Xa2s_dout[20]/_R.0:14   Xa2s_dout[20]/_R.0:16 7.3025 $mt2
Re29848 Xa2s_dout[20]/_R.0:16   Xa2s_dout[20]/_R.0:1 7.1075 $mt2
Re29849 Xa2s_dout[20]/_R.0:9    Xa2s_dout[20]/_R.0:16 6.4000 $mt2
Re29850 Xa2s_dout[19]/_R.0:14   Xa2s_dout[19]/_R.0:16 7.3025 $mt2
Re29851 Xa2s_dout[19]/_R.0:16   Xa2s_dout[19]/_R.0:1 7.1075 $mt2

Re29989 Xa2s_dout[21]/_R.1:32   Xa2s_dout[21]/_R.1:27 7.5288 $mt2
Re29990 Xa2s_dout[21]/_R.1:27   Xa2s_dout[21]/_R.1:19 6.7695 $mt2
Re29992 Xa2s_dout[20]/_R.1:32   Xa2s_dout[20]/_R.1:27 7.5288 $mt2
Re29993 Xa2s_dout[20]/_R.1:27   Xa2s_dout[20]/_R.1:19 6.7695 $mt2
Re29995 Xa2s_dout[19]/_R.1:32   Xa2s_dout[19]/_R.1:27 7.5288 $mt2
Re29996 Xa2s_dout[19]/_R.1:27   Xa2s_dout[19]/_R.1:19 6.7695 $mt2

Re30391 Xa2s_dout[22]/clk0:5    Xa2s_dout[22]/clk0:7 6.4000 $mt2
Re30392 Xa2s_dout[21]/clk0:7    Xa2s_dout[21]/clk0:5 6.4000 $mt2
Re30393 Xa2s_dout[20]/clk0:5    Xa2s_dout[20]/clk0:7 6.4000 $mt2
Re30394 Xa2s_dout[19]/clk0:7    Xa2s_dout[19]/clk0:5 6.4000 $mt2
Re30395 Xa2s_dout[18]/clk0:5    Xa2s_dout[18]/clk0:7 6.4000 $mt2

Re30450 Xa2s_dout[21]/_clk:11   Xa2s_dout[21]/_clk:15 6.4000 $mt2
Re30451 Xa2s_dout[21]/_clk:16   Xa2s_dout[21]/_clk:14 6.4000 $mt2
Re30452 Xa2s_dout[20]/_clk:11   Xa2s_dout[20]/_clk:15 6.4000 $mt2
Re30453 Xa2s_dout[20]/_clk:16   Xa2s_dout[20]/_clk:14 6.4000 $mt2
Re30454 Xa2s_dout[19]/_clk:11   Xa2s_dout[19]/_clk:15 6.4000 $mt2
Re30455 Xa2s_dout[19]/_clk:16   Xa2s_dout[19]/_clk:14 6.4000 $mt2

Re30605 Xa2s_dout[21]/PReset:3  Xa2s_dout[21]/PReset:4 6.4000 $mt2
Re30606 Xa2s_dout[21]/PReset:1  Xa2s_dout[21]/PReset:5 6.4000 $mt2
Re30607 Xa2s_dout[20]/PReset:3  Xa2s_dout[20]/PReset:4 6.4000 $mt2
Re30608 Xa2s_dout[20]/PReset:1  Xa2s_dout[20]/PReset:5 6.4000 $mt2
Re30609 Xa2s_dout[19]/PReset:3  Xa2s_dout[19]/PReset:4 6.4000 $mt2
Re30610 Xa2s_dout[19]/PReset:1  Xa2s_dout[19]/PReset:5 6.4000 $mt2

Re30778 Xa2s_dout[21]/_noR:29   Xa2s_dout[21]/_noR:31 6.4000 $mt2
Re30779 Xa2s_dout[21]/27:1      Xa2s_dout[21]/27:2 13.0785 $mt2
Re30780 Xa2s_dout[20]/_noR:27   Xa2s_dout[20]/_noR:31 6.8872 $mt2
Re30781 Xa2s_dout[20]/_noR:31   Xa2s_dout[20]/_noR:17 7.5105 $mt2
Re30782 Xa2s_dout[20]/_noR:29   Xa2s_dout[20]/_noR:31 6.4000 $mt2
Re30783 Xa2s_dout[20]/27:1      Xa2s_dout[20]/27:2 13.0785 $mt2
Re30784 Xa2s_dout[19]/_noR:27   Xa2s_dout[19]/_noR:31 6.8872 $mt2
Re30785 Xa2s_dout[19]/_noR:31   Xa2s_dout[19]/_noR:17 7.5105 $mt2

Re30875 Xa2s_dout[22]/_Le:7     Xa2s_dout[22]/_Le:3 9.8765 $mt2
Re30876 Xa2s_dout[21]/_Le:7     Xa2s_dout[21]/_Le:3 9.8765 $mt2
Re30877 Xa2s_dout[20]/_Le:7     Xa2s_dout[20]/_Le:3 9.8765 $mt2
Re30878 Xa2s_dout[19]/_Le:7     Xa2s_dout[19]/_Le:3 9.8765 $mt2
Re30879 Xa2s_dout[18]/_Le:7     Xa2s_dout[18]/_Le:3 9.8765 $mt2

Re31261 Xa2s_dout[22]/Rc:10     Xa2s_dout[22]/Rc:1 17.3433 $mt2
Re31262 Xa2s_dout[21]/Rc:10     Xa2s_dout[21]/Rc:1 17.3433 $mt2
Re31263 Xa2s_dout[20]/Rc:10     Xa2s_dout[20]/Rc:1 17.3433 $mt2
Re31264 Xa2s_dout[19]/Rc:10     Xa2s_dout[19]/Rc:1 17.3433 $mt2
Re31265 Xa2s_dout[18]/Rc:10     Xa2s_dout[18]/Rc:1 17.3433 $mt2

Re31432 Xa2s_dout[21]/_R.0:26   Xa2s_dout[21]/_R.0:6 4.1513 $mt2
Re31433 Xa2s_dout[21]/_R.0:25   Xa2s_dout[21]/_R.0:26 6.4000 $mt2
Re31434 Xa2s_dout[20]/_R.0:24   Xa2s_dout[20]/_R.0:26 0.2311 $mt2
Re31435 Xa2s_dout[20]/_R.0:26   Xa2s_dout[20]/_R.0:6 4.1513 $mt2
Re31436 Xa2s_dout[20]/_R.0:25   Xa2s_dout[20]/_R.0:26 6.4000 $mt2
Re31437 Xa2s_dout[19]/_R.0:24   Xa2s_dout[19]/_R.0:26 0.2311 $mt2
Re31438 Xa2s_dout[19]/_R.0:26   Xa2s_dout[19]/_R.0:6 4.1513 $mt2

Re31900 Xa2s_dout[21]/_clk:19   Xa2s_dout[21]/_clk:20 6.4000 $mt2
Re31901 Xa2s_dout[21]/_clk:9    Xa2s_dout[21]/_clk:21 6.4000 $mt2
Re31902 Xa2s_dout[20]/_clk:20   Xa2s_dout[20]/_clk:21 1.7475 $mt2
Re31903 Xa2s_dout[20]/_clk:21   Xa2s_dout[20]/_clk:1 9.4723 $mt2
Re31904 Xa2s_dout[20]/_clk:20   Xa2s_dout[20]/_clk:22 7.0848 $mt2
Re31905 Xa2s_dout[20]/_clk:19   Xa2s_dout[20]/_clk:20 6.4000 $mt2
Re31906 Xa2s_dout[20]/_clk:9    Xa2s_dout[20]/_clk:21 6.4000 $mt2
Re31907 Xa2s_dout[19]/_clk:20   Xa2s_dout[19]/_clk:21 1.7475 $mt2
Re31908 Xa2s_dout[19]/_clk:21   Xa2s_dout[19]/_clk:1 9.4723 $mt2

Re32061 Xa2s_dout[22]/_R.0:28   Xa2s_dout[22]/_R.0:27 7.2180 $mt2
Re32062 Xa2s_dout[21]/_R.0:28   Xa2s_dout[21]/_R.0:27 7.2180 $mt2
Re32063 Xa2s_dout[20]/_R.0:28   Xa2s_dout[20]/_R.0:27 7.2180 $mt2
Re32064 Xa2s_dout[19]/_R.0:28   Xa2s_dout[19]/_R.0:27 7.2180 $mt2
Re32065 Xa2s_dout[18]/_R.0:28   Xa2s_dout[18]/_R.0:27 7.2180 $mt2

Re32095 Xa2s_dout[22]/_grant:6  Xa2s_dout[22]/_grant:2 13.8065 $mt2
Re32096 Xa2s_dout[21]/_grant:6  Xa2s_dout[21]/_grant:2 13.8065 $mt2
Re32097 Xa2s_dout[20]/_grant:6  Xa2s_dout[20]/_grant:2 13.8065 $mt2
Re32098 Xa2s_dout[19]/_grant:6  Xa2s_dout[19]/_grant:2 13.8065 $mt2
Re32099 Xa2s_dout[18]/_grant:6  Xa2s_dout[18]/_grant:2 13.8065 $mt2

Re32127 Xa2s_dout[22]/_R.1:46   Xa2s_dout[22]/_R.1:41 13.9876 $mt2
Re32128 Xa2s_dout[21]/_R.1:46   Xa2s_dout[21]/_R.1:41 13.9876 $mt2
Re32129 Xa2s_dout[20]/_R.1:46   Xa2s_dout[20]/_R.1:41 13.9876 $mt2
Re32130 Xa2s_dout[19]/_R.1:46   Xa2s_dout[19]/_R.1:41 13.9876 $mt2
Re32131 Xa2s_dout[18]/_R.1:46   Xa2s_dout[18]/_R.1:41 13.9876 $mt2

Re32262 Xa2s_dout[21]/21:2      Xa2s_dout[21]/21:3 6.4000 $mt2
Re32263 Xa2s_dout[21]/21:4      Xa2s_dout[21]/21:5 6.4000 $mt2
Re32264 Xa2s_dout[20]/21:1      Xa2s_dout[20]/21:3 6.6785 $mt2
Re32265 Xa2s_dout[20]/21:3      Xa2s_dout[20]/21:5 0.4865 $mt2
Re32266 Xa2s_dout[20]/21:5      Xa2s_dout[20]/21:6 6.8865 $mt2
Re32267 Xa2s_dout[20]/21:2      Xa2s_dout[20]/21:3 6.4000 $mt2
Re32268 Xa2s_dout[20]/21:4      Xa2s_dout[20]/21:5 6.4000 $mt2
Re32269 Xa2s_dout[19]/21:1      Xa2s_dout[19]/21:3 6.6785 $mt2
Re32270 Xa2s_dout[19]/21:3      Xa2s_dout[19]/21:5 0.4865 $mt2

Re32455 Xa2s_dout[21]/15:4      Xa2s_dout[21]/15:12 6.8847 $mt2
Re32457 Xa2s_dout[21]/15:10     Xa2s_dout[21]/15:4 6.4000 $mt2
Re32458 Xa2s_dout[20]/15:5      Xa2s_dout[20]/15:1 7.2227 $mt2
Re32461 Xa2s_dout[20]/15:7      Xa2s_dout[20]/15:1 6.4000 $mt2
Re32463 Xa2s_dout[20]/15:4      Xa2s_dout[20]/15:12 6.8847 $mt2
Re32465 Xa2s_dout[20]/15:10     Xa2s_dout[20]/15:4 6.4000 $mt2
Re32466 Xa2s_dout[19]/15:5      Xa2s_dout[19]/15:1 7.2227 $mt2
Re32469 Xa2s_dout[19]/15:7      Xa2s_dout[19]/15:1 6.4000 $mt2

Re32711 Xa2s_dout[21]/_clk0:35  Xa2s_dout[21]/_clk0:33 6.4000 $mt2
Re32713 Xa2s_dout[21]/_clk0:34  Xa2s_dout[21]/_clk0:31 6.4000 $mt2
Re32714 Xa2s_dout[20]/15:13     Xa2s_dout[20]/15:2 6.4000 $mt2
Re32716 Xa2s_dout[20]/_clk0:33  Xa2s_dout[20]/_clk0:38 0.6384 $mt2
Re32717 Xa2s_dout[20]/_clk0:38  Xa2s_dout[20]/_clk0:17 7.2223 $mt2
Re32718 Xa2s_dout[20]/_clk0:38  Xa2s_dout[20]/_clk0:27 7.0093 $mt2
Re32719 Xa2s_dout[20]/_clk0:35  Xa2s_dout[20]/_clk0:33 6.4000 $mt2
Re32721 Xa2s_dout[20]/_clk0:34  Xa2s_dout[20]/_clk0:31 6.4000 $mt2
Re32722 Xa2s_dout[19]/15:13     Xa2s_dout[19]/15:2 6.4000 $mt2
Re32724 Xa2s_dout[19]/_clk0:33  Xa2s_dout[19]/_clk0:38 0.6384 $mt2

Re32928 Xa2s_dout[21]/17:7      Xa2s_dout[21]/17:3 6.8900 $mt2
Re32929 Xa2s_dout[21]/17:5      Xa2s_dout[21]/17:7 6.4000 $mt2
Re32930 Xa2s_dout[20]/17:7      Xa2s_dout[20]/17:1 6.6820 $mt2
Re32931 Xa2s_dout[20]/17:7      Xa2s_dout[20]/17:3 6.8900 $mt2
Re32932 Xa2s_dout[20]/17:5      Xa2s_dout[20]/17:7 6.4000 $mt2
Re32933 Xa2s_dout[19]/17:7      Xa2s_dout[19]/17:1 6.6820 $mt2
Re32934 Xa2s_dout[19]/17:7      Xa2s_dout[19]/17:3 6.8900 $mt2

Re33145 Xa2s_dout[21]/clk0:17   Xa2s_dout[21]/clk0:36 6.4000 $mt2
Re33146 Xa2s_dout[21]/clk0:12   Xa2s_dout[21]/clk0:37 6.4000 $mt2
Re33148 Xa2s_dout[20]/clk0:34   Xa2s_dout[20]/clk0:35 6.5463 $mt2
Re33149 Xa2s_dout[20]/clk0:35   Xa2s_dout[20]/clk0:36 1.7973 $mt2
Re33150 Xa2s_dout[20]/clk0:36   Xa2s_dout[20]/clk0:37 0.4735 $mt2
Re33151 Xa2s_dout[20]/clk0:37   Xa2s_dout[20]/clk0:8 1.5578 $mt2
Re33152 Xa2s_dout[20]/clk0:8    Xa2s_dout[20]/clk0:10 6.7442 $mt2
Re33153 Xa2s_dout[20]/clk0:35   Xa2s_dout[20]/clk0:21 7.4666 $mt2
Re33154 Xa2s_dout[20]/clk0:17   Xa2s_dout[20]/clk0:36 6.4000 $mt2
Re33155 Xa2s_dout[20]/clk0:12   Xa2s_dout[20]/clk0:37 6.4000 $mt2
Re33157 Xa2s_dout[19]/clk0:34   Xa2s_dout[19]/clk0:35 6.5463 $mt2
Re33158 Xa2s_dout[19]/clk0:35   Xa2s_dout[19]/clk0:36 1.7973 $mt2

Re33351 Xa2s_dout[22]/_clk0:62  Xa2s_dout[22]/_clk0:56 13.1695 $mt2
Re33352 Xa2s_dout[21]/_clk0:62  Xa2s_dout[21]/_clk0:56 13.1695 $mt2
Re33353 Xa2s_dout[20]/_clk0:62  Xa2s_dout[20]/_clk0:56 13.1695 $mt2
Re33354 Xa2s_dout[19]/_clk0:62  Xa2s_dout[19]/_clk0:56 13.1695 $mt2
Re33355 Xa2s_dout[18]/_clk0:62  Xa2s_dout[18]/_clk0:56 13.1695 $mt2

Rd16556 Xa2s_dout[22]/_Le:3     Xa2s_dout[22]/_Le:2 15.0740 $mt3
Rd16557 Xa2s_dout[21]/_Le:3     Xa2s_dout[21]/_Le:2 15.0740 $mt3
Rd16558 Xa2s_dout[20]/_Le:3     Xa2s_dout[20]/_Le:2 15.0740 $mt3
Rd16559 Xa2s_dout[19]/_Le:3     Xa2s_dout[19]/_Le:2 15.0740 $mt3
Rd16560 Xa2s_dout[18]/_Le:3     Xa2s_dout[18]/_Le:2 15.0740 $mt3

Rd16592 Xa2s_dout[22]/_R.0:5    Xa2s_dout[22]/_R.0:6 13.3645 $mt3
Rd16593 Xa2s_dout[21]/_R.0:5    Xa2s_dout[21]/_R.0:6 13.3645 $mt3
Rd16594 Xa2s_dout[20]/_R.0:5    Xa2s_dout[20]/_R.0:6 13.3645 $mt3
Rd16595 Xa2s_dout[19]/_R.0:5    Xa2s_dout[19]/_R.0:6 13.3645 $mt3
Rd16596 Xa2s_dout[18]/_R.0:5    Xa2s_dout[18]/_R.0:6 13.3645 $mt3

Rd16826 Xa2s_dout[21]/_R.1:28   Xa2s_dout[21]/_R.1:26 7.6015 $mt3
Rd16827 Xa2s_dout[21]/_R.1:25   Xa2s_dout[21]/_R.1:28 6.4000 $mt3
Rd16828 Xa2s_dout[20]/_R.1:27   Xa2s_dout[20]/_R.1:28 9.8635 $mt3
Rd16829 Xa2s_dout[20]/_R.1:28   Xa2s_dout[20]/_R.1:26 7.6015 $mt3
Rd16830 Xa2s_dout[20]/_R.1:25   Xa2s_dout[20]/_R.1:28 6.4000 $mt3
Rd16831 Xa2s_dout[19]/_R.1:27   Xa2s_dout[19]/_R.1:28 9.8635 $mt3
Rd16832 Xa2s_dout[19]/_R.1:28   Xa2s_dout[19]/_R.1:26 7.6015 $mt3

Rd16982 Xa2s_dout[22]/0:6       Xa2s_dout[22]/0:1 13.8065 $mt3
Rd16983 Xa2s_dout[21]/0:6       Xa2s_dout[21]/0:1 13.8065 $mt3
Rd16984 Xa2s_dout[20]/0:6       Xa2s_dout[20]/0:1 13.8065 $mt3
Rd16985 Xa2s_dout[19]/0:6       Xa2s_dout[19]/0:1 13.8065 $mt3
Rd16986 Xa2s_dout[18]/0:6       Xa2s_dout[18]/0:1 13.8065 $mt3

Rd17289 Xa2s_dout[22]/clk0:7    Xa2s_dout[22]/clk0:8 15.1975 $mt3
Rd17290 Xa2s_dout[21]/clk0:7    Xa2s_dout[21]/clk0:8 15.1975 $mt3
Rd17291 Xa2s_dout[20]/clk0:7    Xa2s_dout[20]/clk0:8 15.1975 $mt3
Rd17292 Xa2s_dout[19]/clk0:7    Xa2s_dout[19]/clk0:8 15.1975 $mt3
Rd17293 Xa2s_dout[18]/clk0:7    Xa2s_dout[18]/clk0:8 15.1975 $mt3

Rd17321 Xa2s_dout[22]/_clk:15   Xa2s_dout[22]/_clk:16 14.5475 $mt3
Rd17322 Xa2s_dout[21]/_clk:15   Xa2s_dout[21]/_clk:16 14.5475 $mt3
Rd17323 Xa2s_dout[20]/_clk:15   Xa2s_dout[20]/_clk:16 14.5475 $mt3
Rd17324 Xa2s_dout[19]/_clk:15   Xa2s_dout[19]/_clk:16 14.5475 $mt3
Rd17325 Xa2s_dout[18]/_clk:15   Xa2s_dout[18]/_clk:16 14.5475 $mt3

Rd17431 Xa2s_dout[22]/PReset:3  Xa2s_dout[22]/PReset:5 16.2570 $mt3
Rd17432 Xa2s_dout[21]/PReset:3  Xa2s_dout[21]/PReset:5 16.2570 $mt3
Rd17433 Xa2s_dout[20]/PReset:3  Xa2s_dout[20]/PReset:5 16.2570 $mt3
Rd17434 Xa2s_dout[19]/PReset:3  Xa2s_dout[19]/PReset:5 16.2570 $mt3
Rd17435 Xa2s_dout[18]/PReset:3  Xa2s_dout[18]/PReset:5 16.2570 $mt3

Rd17682 Xa2s_dout[22]/_R.0:27   Xa2s_dout[22]/_R.0:24 16.0490 $mt3
Rd17683 Xa2s_dout[21]/_R.0:27   Xa2s_dout[21]/_R.0:24 16.0490 $mt3
Rd17684 Xa2s_dout[20]/_R.0:27   Xa2s_dout[20]/_R.0:24 16.0490 $mt3
Rd17685 Xa2s_dout[19]/_R.0:27   Xa2s_dout[19]/_R.0:24 16.0490 $mt3
Rd17686 Xa2s_dout[18]/_R.0:27   Xa2s_dout[18]/_R.0:24 16.0490 $mt3

Rd17994 Xa2s_dout[21]/15:2      Xa2s_dout[21]/15:3 6.4000 $mt3
Rd17995 Xa2s_dout[21]/_clk0:33  Xa2s_dout[21]/_clk0:34 14.2875 $mt3
Rd17996 Xa2s_dout[20]/15:1      Xa2s_dout[20]/15:3 6.8865 $mt3
Rd17997 Xa2s_dout[20]/15:3      Xa2s_dout[20]/15:4 7.3415 $mt3
Rd17998 Xa2s_dout[20]/15:2      Xa2s_dout[20]/15:3 6.4000 $mt3
Rd17999 Xa2s_dout[20]/_clk0:33  Xa2s_dout[20]/_clk0:34 14.2875 $mt3
Rd18000 Xa2s_dout[19]/15:1      Xa2s_dout[19]/15:3 6.8865 $mt3
Rd18001 Xa2s_dout[19]/15:3      Xa2s_dout[19]/15:4 7.3415 $mt3
C99     init_wait.cnt[12]:30    init_wait.cnt[13]:27 8.657E-17
C100    Xa2s_dout[20]/_R.1:29   odq[20]:22 6.778E-18
C240    Xa2s_dout[27]/8:1       Xa2s_dout[27]/_R.1:39 2.105E-20
C241    GND!    Xopctrl.A2Sop/Lc[0][9].e:8 1.211E-15
C242    Xa2s_dout[20]/_R.1:28   Xa2s_dout[20]/_R.0:12 1.243E-17
C243    Xconfigure.a2s/Xdyb[6]/32:11    Xconfigure.a2s/Lc[2][6].1:9
+	 6.084E-18
C483    Xdll/Xdetect[3]/g2:3    Xdll/Xdetect[3]/g2:5 1.929E-17
C484    Xa2s_dout[20]/_R.0:25   Xa2s_dout[20]/_clk0:30 3.265E-17
C485    Xconfigure.a2s/Xdyb[6]/_lv01:1  Xconfigure.a2s/cRl[2][1].0:79
+	 1.238E-18
C680    GND!    Xopctrl.nopctrl/Xgereg/Xlatch/Xlatchv/12 3.308E-18
C681    Xa2s_dout[20]/_clk:28   Xa2s_dout[20]/21:3 3.947E-19
C682    Xopctrl.A2Sop/XbufL[6][0]/_b.0:6        
+	Xopctrl.A2Sop/XbufL[6][0]/_b.0:10 1.249E-17
C870    Xconfigure.a2s/cRl[2][2].0:69   Xconfigure.a2s/Lc[2][9].0:12
+	 1.802E-19
C871    Xa2s_dout[20]/8:2       Xa2s_dout[20]/8:5 3.957E-18
C872    Xrefresh_gen.inc0/Xincbit[2]/Xreg/Xdelay/Xdelay[2]/x:3  Vdd!
+	 6.545E-16
C947    Xdqsgen[1]/Xalt_dqs/x.0:16      Vdd! 3.779E-17
C948    Xdll/d:1290     Xdll/Xphased_fclk[0]/n[1][12]:4 4.852E-22
C949    clk:4342        Xa2s_dout[20]/Rc:12 6.649E-20
C950    Xa2s_dm[3]/_Le:8        GND! 9.155E-17
C2536   Xdll/Xctrl/Xcounter/Xcounter/cnt[4]:5   
+	Xdll/Xctrl/Xcounter/Xcounter/Xrb/_co35:6 1.368E-17
C2537   Xa2s_dout[20]/_clk0:29  clk:4975 2.864E-21
C2538   Xinit_wait.dffinit/Xolatch/Xlatchv/_v:29        
+	Xinit_wait.dffinit/Xolatch/Xlatchv/_in:11 1.383E-17
C4937   Xopconv[11]/_r.1:22     Xopconv[11]/_r.1:30 1.284E-18
C4938   Xa2s_dout[20]/8:2       Xa2s_dout[20]/9:2 4.046E-19
C4939   Xs2a_din[13]/5:4        Xs2a_din[13]/5:5 3.957E-18
C4940   Vdd!    Xopctrl.opreg[6]/x:5 4.733E-16
C5977   Xdll/Xctrl/Xcounter/Xcounter/Xincbit[4]/dq:2    
+	Xdll/Xctrl/Xcounter/Xcounter/Xincbit[4]/__rst:7 9.927E-18
C5978   Xa2s_dout[20]/_R.0:16   Xa2s_dout[20]/_r:17 6.764E-17
C5979   Xlatency_ctrl.oeD/Xvdelay[0]/Xplatch/Xlatchv/4:2        GND!
+	 1.053E-16
C6088   Xa2s_dout[20]/1:3       Xa2s_dout[20]/0:7 3.195E-17
C6089   opctrl.xop[0][25]:5     opctrl._opload:117 5.595E-16
C6090   Xopconv[5]/_r.3:12      op4[5].3:12 5.575E-17
C6642   Vdd!    Xophold[6]/Xilatch/Xlatchv/v:11 5.167E-17
C6643   Xa2s_dout[23]/_clk:23   GND! 5.764E-16
C6644   Xa2s_dout[20]/1:4       Xa2s_dout[20]/1:3 2.107E-18
C6645   refresh_gen.cnt[6]:49   _PReset!:6919 1.180E-18
C6646   Xa2s_dm[2]/clk0:24      Xa2s_dm[2]/clk0:23 1.544E-18
C7357   Xconfigure.a2s/Lc[2][11].3:3    Xconfigure.a2s/Lc[2][11].3:2
+	 4.733E-17
C7358   Xa2s_dout[20]/29:2      Xa2s_dout[20]/_clk0:17 3.221E-19
C7359   Xopctrl.A2Sop/XcL/LD4[1].0:2    Xopctrl.A2Sop/XcL/LD[4].0:6
+	 3.909E-17
C7551   Xconfigure.a2s/Xdyb[3]/r[1].0:2 _SReset!:347 5.331E-18
C7552   odq[7]  Vdd! 3.016E-16
C7553   Xa2s_dout[20]/_clk:23   GND! 5.764E-16
C7554   Xopctrl.A2Sop/XcL/XdetectL[6]/9:1       
+	Xopctrl.A2Sop/XcL/XdetectL[6]/_R:17 5.684E-17
C7623   _PReset!:915    Xconfigure.a2s/Lc[1][10].0:8 5.796E-18
C7624   Xopctrl.A2Sop/Lc[2][13].2:23    _SReset!:3114 1.203E-17
C7625   Xa2s_dout[20]/_clk:24   GND! 2.066E-16
C7626   Xa2s_dout[0]/17:3       Xa2s_dout[0]/15:1 1.093E-17
C7689   Xdll/Xphased_fclk[0]/n[7][3]:4  GND! 4.338E-16
C7690   op2[3].0:2      op2[2].1:5 1.952E-17
C7691   Xa2s_dout[20]/_clk:25   GND! 2.425E-16
C7692   Xclk_ramp/c[3]:15       clk:1922 2.312E-16
C7693   clk:886 Xopctrl.A2Sop/Xdyb[13]/_R[0]:24 2.797E-17
C7829   Xdll/Xphased_fclk[7]/Xdemux/demux._R[6]:1       GND! 2.000E-18
C7830   Xa2s_dout[20]/_grant:3  clk:4275 1.209E-17
C7831   _SReset!:2112   op4[2].3:35 9.446E-18
C7832   Xlatency_ctrl.oeD/Xvdelay[0]/Xmux/_insel[0]:14  GND! 9.996E-16
C8821   Xs2a_din[18]/go:39      Xs2a_din[18]/_clk0:11 3.551E-17
C8822   Xa2s_dout[20]/_R.0:6    Xa2s_dout[20]/Rv:4 4.288E-16
C8823   Xopctrl.A2Sop/Lc[2][10].1:6     
+	Xopctrl.A2Sop/XbufL[10][1]/_c_01:4 1.582E-17
C9820   Xdll/Xphased_fclk[1]/Xdunit[4][2]/n[1]:7        
+	Xdll/Xphased_fclk[1]/n[4][3]:7 4.938E-19
C9821   _PReset!:6825   Xa2s_dout[20]/17:1 4.053E-18
C9822   Xopctrl.A2Sop/XbufL[14][0]/_ae:15       
+	Xopctrl.A2Sop/Lc[0][14].e:19 4.422E-17
C9952   Xconfigure.a2s/Xdyb[9]/_en:19   Xconfigure.a2s/Xdyb[9]/_en:22
+	 1.757E-18
C9953   clk:4579        Xa2s_dout[20]/_clk:11 3.709E-17
C9954   op4[6].3        Xopctrl.A2Sop/XbufL[7][0]/_ce:8 2.370E-16
C9955   Xs2a_din[11]/_req:5     Xs2a_din[11]/go:11 8.042E-18
C10151  Xconfigure.a2s/Xdyb[10]/lv:2    Vdd! 7.561E-17
C10152  ddqs[0]:165     Xs2a_din[1]/_clk0:9 2.394E-17
C10153  Xa2s_dout[20]/clk0:23   Xa2s_dout[20]/_clk0:50 4.157E-17
C10154  Xopctrl.opreg[4]/Xolatch/Xlatchv/s:11   
+	Xopctrl.opreg[4]/_clk:1 7.158E-18
C10570  Xdqsgen[0]/Xalt_dqs/x.0:34      Xdqsgen[0]/async_dqs[0].e:17
+	 3.440E-21
C10571  Xa2s_dout[20]/_r:17     Xa2s_dout[20]/_r:18 7.012E-19
C10572  Xconfigure.a2s/XbufL[4][0]/_ce:12       
+	Xconfigure.a2s/XbufL[4][0]/_b.0:8 5.316E-18
C10601  Xdll/Xphased[2]/Xdunit[3][0]/n[0]:3     
+	Xdll/Xphased[2]/Xdunit[3][0]/n[1]:2 6.968E-17
C10602  dout[22].1:4    Xa2s_dout[20]/17:5 1.635E-18
C10603  Xdll/Xphased_fclk[3]/Xdunit[2][5]/n[1]:3        
+	Xdll/Xphased_fclk[3]/Xdunit[2][5]/n[1]:2 3.835E-18
C10741  Xrefresh_gen.inc0/Xincbit[3]/xnor._L[1]:9       clk:2137
+	 2.859E-19
C10742  Xa2s_dout[20]/6:1       Xa2s_dout[20]/_noR:10 6.288E-18
C11034  Xdll/d:2016     GND! 2.714E-16
C11035  Xa2s_dout[2]/_clk:11    Xa2s_dout[2]/29:1 5.696E-18
C11036  Xa2s_dout[20]/27:2      Xa2s_dout[20]/_clk0:24 9.551E-17
C11037  opctrl._opload:363      opctrl.blen[2]:1 1.680E-18
C11554  start:26        Xrefresh_gen.inc0/Xincbit0/Xtreg/Xdelay/x[3]:1
+	 4.769E-17
C11555  Xa2s_dout[20]/_R.1:27   Xa2s_dout[20]/_R.1:18 2.881E-17
C11556  Xopctrl.A2Sop/XbufL[13][0]/_b.2:1       
+	Xopctrl.A2Sop/Lc[1][13].2:14 4.702E-17
C11639  Xdqsgen[2]/Xalt_dqs/_r.0:4      Vdd! 1.304E-17
C11640  GND!    dllclk:19 8.265E-18
C11641  Xa2s_dout[20]/_R.1:16   Xa2s_dout[20]/Rv:4 2.894E-18
C11642  Xopctrl.nopctrl/Xnopcntr/Xcounter/Xincbit[2]/dq:2       
+	Xopctrl.nopctrl/Xnopcntr/Xcounter/Xincbit[2]/__rst:2 2.940E-17
C12027  Xdqsgen[0]/Xalt_dqs/_r.0:4      Vdd! 1.304E-17
C12028  Xopctrl.A2Sop/XbufL[10][1]/be:6 _SReset!:2420 3.142E-17
C12029  Xa2s_dout[20]/_Le:15    dout[22].e:6 3.258E-17
C12030  Xconfigure.a2s/Xdyb[2]/_R[1]:1  Xconfigure.a2s/Xdyb[2]/_clk:4
+	 1.867E-17
C12308  Xopctrl.opreg[18]/Xolatch/Xlatchv/s:6   GND! 1.407E-16
C12309  Xa2s_dout[20]/31:2      Xa2s_dout[20]/clk0:16 4.744E-17
C12310  Xinv[6]/x:6     Vdd! 7.738E-18
C12875  Xdll/Xctrl/Xcounter/Xcounter/Xincbit[1]/Xreg/x:13       
+	Xdll/Xctrl/Xcounter/cnt[1]:30 2.110E-17
C12876  Xa2s_dout[20]/_clk0:26  dout[22].1:5 2.410E-17
C13989  Xa2s_dout[20]/_R.1:17   Xa2s_dout[20]/Rv:4 6.375E-18
C14401  Xa2s_dout[24]/_R.1:27   Xa2s_dout[24]/_clk:1 3.802E-17
C14402  odq[30]:19      _SReset!:5089 2.729E-18
C14403  Xa2s_dout[20]/_clk:31   oe:293 1.472E-20
C14404  Vdd!    Xinv[2]/x:7 6.450E-18
C14405  Xa2s_dout[8]/8:1        Xa2s_dout[8]/_R.1:39 2.105E-20
C15228  Xa2s_dout[20]/15:7      Xa2s_dout[20]/clk0:27 4.177E-18
C15229  Xdll/Xphased_fclk[4]/Xdunit[7][3]/n[0]:3        
+	Xdll/Xphased_fclk[4]/Xdunit[7][3]/n[1]:4 2.556E-18
C15521  Xopctrl.opreg[6]/x:13   GND! 4.137E-17
C15522  Xa2s_dout[20]/__Le:3    Xa2s_dout[20]/7:5 1.478E-17
C15523  Xdll/Xctrl/Xcounter/Xcounter/Xincbit[4]/d:42    
+	Xdll/Xctrl/Xcounter/Xcounter/inc[4]:30 2.568E-18
C15583  GND!    dout[18].0:1 3.995E-16
C15584  NRFRSH[7]       Xopctrl.A2Sop/Rl.e:18 1.793E-17
C15585  Xa2s_dout[20]/_R.0:31   Xa2s_dout[20]/10:3 3.672E-20
C15586  Xdll/Xctrl/refclk:226   Xdll/Xctrl/refclk:225 2.794E-17
C17457  Xdll/Xphased_fclk[2]/Xdunit[1][8]/n[0]:3        Vdd! 1.414E-16
C17458  _PReset!:6825   Xa2s_dout[20]/_R.0:28 4.141E-17
C17459  Xlatency_ctrl.dqsenH/Xdelay/Xdelay[1]/Xdelay[0]/x:1     Vdd!
+	 1.763E-16
C17824  Xconfigure.a2s/Xdyb[4]/9:1      
+	Xconfigure.a2s/Xdyb[4]/rvb[0]:4 2.116E-20
C17825  Xa2s_dout[20]/_R.0:24   clk:4493 5.101E-17
C17826  Xdll/Xphased_fclk[2]/Xdunit[1][2]/n[0]:3        Vdd! 1.419E-16
C17827  GND!    Xramp_odqs[1]/x:22 7.163E-18
C17954  Xlatency_ctrl.ieD/Xvdelay[4]/Xplatch/Xlatchv/5:1        GND!
+	 9.296E-17
C17955  Xa2s_dout[20]/_grant:6  Xa2s_dout[20]/_clk0:35 3.009E-18
C17956  Xconfigure.a2s/XbufL[10][1]/10:5        
+	Xconfigure.a2s/Lc[2][10].0:38 5.276E-17
C18739  Xdll/d:6418     Xdll/Xphased_fclk[1]/Xdunit[3][6]/n[0]:1
+	 2.560E-17
C18740  Xa2s_dout[20]/_clk0:25  GND! 3.432E-16
C18872  Xopctrl.opreg[5]/Xolatch/Xlatchv/_out:12        sop[0][5]:27
+	 5.172E-17
C18873  Xa2s_dout[20]/_clk0:19  clk:4029 4.103E-18
C18874  init_wait.cnt[4]:21     Xinit_wait.cntr0/Xincbit[1]/6
+	 4.666E-20
C19162  Xs2a_din[21]/_Rv:4      Xs2a_din[21]/_clk0:18 9.253E-17
C19163  Xa2s_dout[20]/_R.0:27   Xa2s_dout[20]/_clk0:27 1.918E-17
C19164  _PReset!:4779   Xopctrl.rdwr_ctrl/Xbl_counter/cnt[3]:6
+	 3.796E-18
C19174  Xophold[5]/x:44 Xophold[5]/Xolatch/Xlatchv/_v:24 4.284E-18
C19175  oe:498  Xa2s_dout[20]/_clk0:43 2.519E-17
C19176  Vdd!    configure.grantinv.R 1.779E-16
C19177  sop[0][0]:4     Xopctrl.opmux[0]/_insel[0]:1 6.009E-18
C20140  Xinit_wait.cntr0/Xincbit[7]/xnor._L[0]:5        
+	init_wait.cnt[7]:22 2.228E-18
C20141  Xa2s_dout[20]/_clk0:11  Xa2s_dout[20]/PReset:1 2.528E-19
C20142  w_gol:24        Xlatency_ctrl.oeD/Xvdelay[0]/Xmux/_sel:8
+	 6.454E-17
C20296  _SReset!:3509   Xdll/Xphased[1]/n[2][13]:4 6.387E-19
C20297  clk:3212        Xophold[2]/_clk:22 9.387E-17
C20298  _PReset!:6825   Xa2s_dout[20]/17:5 2.155E-18
C20299  Xdll/d:1732     Xdll/d:1731 3.187E-17
C20300  Xopctrl.rdwr_ctrl/rw:42 GND! 1.924E-16
C20675  op2[12].0:16    op2[12].1:8 2.916E-17
C20676  Xa2s_dout[20]/clk0:23   Xa2s_dout[20]/_clk0:54 5.466E-17
C20677  Xdll/Xphased[0]/Xdunit[2][13]/n[1]:4    Xdll/r.5:107 2.996E-22
C21407  _SReset!:377    
+	Xlatency_ctrl.dqsenH/Xdelay/Xlatch[1]/Xlatchv/_in:2 1.312E-17
C21408  Xa2s_dout[20]/_clk0:14  Xa2s_dout[20]/_clk:15 1.026E-17
C21409  Xinvdm[3]/x:22  Xinvdm[3]/x:21 3.278E-17
C21410  Xs2a_din[13]/_R.0:3     Xs2a_din[13]/_skip:2 6.364E-17
C21476  clk:4756        GND! 2.258E-16
C21477  Vdd!    chan_dll.ri[7] 1.428E-16
C21478  clk:4579        Xa2s_dout[20]/31:1 2.847E-17
C21479  Xdll/Xphased_fclk[3]/n[4][4]:4  
+	Xdll/Xphased_fclk[3]/Xdunit[4][4]/n[0]:4 3.845E-17
C23361  Xconfigure.a2s/Xctrl/Lvg[1]:28  Xconfigure.a2s/Xctrl/t:20
+	 3.189E-17
C23362  Xa2s_dout[20]/21:5      Xa2s_dout[20]/clk0:33 7.340E-18
C23363  Xdll/Xphased_fclk[4]/n[3][4]:5  
+	Xdll/Xphased_fclk[4]/Xdunit[3][4]/n[1]:1 3.875E-19
C23536  Xa2s_dout[29]/_clk0:24  Xa2s_dout[29]/27:1 1.499E-16
C23537  Xdll/Xdetect[1]/g1:5    Xdll/dclk[0]:202 9.209E-19
C23538  Xa2s_dout[20]/_clk0:26  GND! 3.199E-16
C23539  Xopconv[3]/_r.0:10      Xopconv[3]/_r.1:11 4.820E-16
C23540  clk:1430        Xopctrl.opreg[3]/x:45 3.992E-18
C24315  clk:2552        _PReset!:5386 6.673E-17
C24316  Xopctrl.opreg[20]/Xolatch/Xlatchv/_out:32       GND! 2.757E-16
C24317  _SReset!:5457   Xa2s_dout[20]/17:5 1.055E-17
C24318  Xa2s_dm[2]/clk0:27      dout[26].0:6 1.643E-16
C24393  chan_dll.rden:112       Xdll/Xctrl/Xmux_r[3]/7 3.608E-18
C24394  Xa2s_dout[12]/_r:9      Xa2s_dout[12]/_r:12 1.846E-18
C24395  Xa2s_dout[20]/10:3      Xa2s_dout[20]/_clk0:50 4.882E-19
C24396  Xopctrl.A2Sop/Lc[0][9].e:8      op4[9].0:23 2.516E-17
C24397  Xinvdq[4]/x:10  Vdd! 8.336E-16
C25424  Xdll/Xphased_fclk[4]/Xdunit[3][4]/n[1]:3        
+	Xdll/Xphased_fclk[4]/Xdunit[3][4]/n[1]:2 3.835E-18
C25425  Xa2s_dout[20]/_R.0:33   Xa2s_dout[20]/_clk0:31 7.520E-17
C25426  _SReset!:5543   Xinvdq[13]/x:17 8.834E-19
C25427  Xs2a_din[0]/_clk0:17    ie[3]:549 7.684E-18
C26078  Xrefresh_gen.inc0/Xincbit[1]/Xreg/Xlatch/Xlatchv/PReset:14
+	refresh_gen.cnt[1]:28 2.370E-19
C26079  Xa2s_dout[20]/_R.0:27   Xa2s_dout[20]/_clk:28 2.591E-18
C26080  Xdll/Xphased[3]/n[6][0]:5       
+	Xdll/Xphased[3]/Xdunit[6][0]/n[1]:1 3.606E-19
C26206  GND!    Xdll/Xphased[3]/Xmux/_sl[6]:1 1.308E-16
C26207  Xdll/d:4779     Xdll/d:5013 1.886E-18
C26208  Xa2s_dout[20]/_grant:4  clk:4579 9.983E-19
C26209  Xophold[13]/Xilatch/Xlatchv/_out:42     
+	Xophold[13]/Xilatch/Xlatchv/_out:6 8.948E-18
C26631  clk:2420        Xophold[10]/Xilatch/Xlatchv/_in:11 2.061E-16
C26632  GND!    Xdqsgen[1]/Xdqs_buf/20 6.369E-18
C26633  Xa2s_dout[20]/_clk0:31  Xa2s_dout[20]/clk0:24 1.143E-17
C26634  Xophold[8]/Xilatch/Xlatchv/3:4  
+	Xophold[8]/Xilatch/Xlatchv/_v:18 1.202E-18
+	Xdll/Xctrl/start:47 1.701E-17
C27384  chan_dll.dpass:2        Xdll/__dfclk[1]:9 7.506E-19
C27385  Xa2s_dout[20]/_R.0:12   Xa2s_dout[20]/_R.1:22 1.074E-16
C27386  _SReset!:814    Xconfigure.a2s/XbufL[5][0]/_b.1:25 2.510E-18
C27387  Xconfigure.a2s/Xdyb[6]/r[1].1:8 Vdd! 2.720E-16
C27591  invdq[11].R     GND! 2.510E-16
C27592  Xinit_wait.cntr0/Xincbit0/xnor._L[1]:8  Vdd! 2.487E-17
C27593  Xa2s_dout[20]/_R.1:9    Xa2s_dout[20]/_r:12 6.972E-18
C27594  Vdd!    Xopctrl.rdwr_ctrl/Xbl_counter/cnt[3]:18 5.096E-16
C27595  Xophold[3]/x:49 Xophold[3]/Xolatch/Xlatchv/_l:13 6.888E-17
C27610  Xdll/Xphased[3]/n[2][13]:5      
+	Xdll/Xphased[3]/Xdunit[2][13]/n[0]:1 2.966E-17
C27611  Xa2s_dout[20]/_clk:19   Xa2s_dout[20]/_clk:24 1.579E-17
C27612  Xdll/Xphased_fclk[7]/Xdunit[1][14]/n[1]:4       
+	Xdll/Xphased_fclk[7]/n[1][15]:5 1.872E-21
C28032  clk:3507        Xa2s_dout[12]/_r:9 3.548E-17
C28033  _SReset!:2326   _SReset!:2312 1.060E-16
C28034  Xa2s_dout[20]/_clk0:30  Xa2s_dout[20]/clk0:18 3.588E-17
C28035  Xopctrl.A2Sop/Lc[2][9].e:29     Xopctrl.A2Sop/Lc[2][11].3:8
+	 8.574E-18
C29566  Xophold[2]/Xolatch/Xlatchv/_v:26        GND! 1.358E-16
C29567  Xa2s_dout[20]/_Le:2     Xa2s_dout[20]/55 3.955E-18
C29568  Xopctrl.A2Sop/XbufRl1[1]/la:3   Xopctrl.A2Sop/XbufRl1[1]/3:2
+	 1.124E-17
C30533  GND!    ie[3]:496 2.549E-17
C30534  Xopctrl.opreg[16]/Xolatch/Xlatchv/_v:14 Vdd! 9.208E-17
C30535  Xa2s_dout[20]/_R.1:1    Xa2s_dout[20]/_r:16 9.862E-18
C30536  _PReset!:6916   Xdll/Xphased_fclk[0]/n[3][0]:11 7.954E-19
C30537  NRFRSH[1]:7     _PReset!:4640 3.722E-17
C30805  Xconfigure.a2s/XcL/LD[3].0:8    Xconfigure.a2s/XcL/LD[1].0:6
+	 8.070E-16
C30806  Xa2s_dout[20]/clk0:15   GND! 3.236E-16
C31171  start:54        start:55 4.707E-19
C31172  Xdll/d:1839     Xdll/Xphased_fclk[2]/Xdunit[2][12]/0 8.293E-18
C31173  _SReset!:5269   Xa2s_dout[20]/PReset:6 9.483E-18
C31174  Xinit_wait.cntr1/inc[6]:2       Xinit_wait.cntr1/inc[6]:7
+	 1.747E-17
C31555  Xa2s_dout[20]/PReset:5  Xa2s_dout[20]/clk0:8 2.569E-17
C31556  Xdll/d:816      Xdll/dclk[0]:54 3.124E-17
C31557  Xdll/d:113      GND! 6.389E-16
C31663  Xopctrl.opreg[22]/x:38  GND! 1.845E-16
C31664  _PReset!:5451   Xophold[0]/Xilatch/Xlatchv/_l:11 2.147E-17
C31665  Xa2s_dout[20]/_R.0:25   clk:4493 6.674E-17
C31666  GND!    Xconfigure.a2s/Xdyb[11]/_x[1].0:30 5.442E-19
C31667  GND!    Xdll/dclk[4]:117 1.218E-18
C31882  Xopctrl.opreg[21]/Xolatch/Xlatchv/l:4   GND! 2.278E-16
C31883  opctrl.xop[1][12]:28    clk:1036 1.294E-16
C31884  Xa2s_dout[20]/__Le:7    _SReset!:5034 9.327E-18
C31885  GND!    Xconfigure.a2s/Xdyb[11]/_x[1].1:34 2.185E-17
C33399  Xophold[17]/_clk:7      Xophold[17]/Xolatch/Xlatchv/s:13
+	 7.341E-19
C33400  dout[22].1:1    Xa2s_dout[20]/8:5 3.805E-18
C33401  Xophold[16]/Xilatch/Xlatchv/_in:15      
+	Xophold[16]/Xilatch/Xlatchv/_in:6 4.319E-17
C33900  Xdll/Xphased_fclk[7]/n[6][1]:4  Xdll/d:4063 4.338E-18
C33901  Xa2s_dout[20]/clk0:28   Xa2s_dout[20]/15:7 5.908E-17
C33902  din[20].1       GND! 2.028E-17
C34825  Xdll/Xctrl/Xcounter_lock/Xincbit[3]/and._R:8    
+	Xdll/Xctrl/Xcounter_lock/inc[3]:15 7.391E-17
C34826  clk:4717        Xa2s_dout[20]/21:4 6.166E-18
C34827  Xa2s_dout[10]/_clk0:58  Xa2s_dout[10]/15:12 3.148E-18
C36558  Xs2a_din[27]/go:14      Xs2a_din[27]/go:13 6.201E-19
C36559  Xa2s_dout[20]/__Le:5    Xa2s_dout[20]/Rv:1 1.034E-19
C36560  Xopctrl.opmux[15]/_insel[0]:3   GND! 2.594E-16
C36561  clk:4353        clk:4038 7.169E-19
C36731  GND!    Xconfigure.a2s/Xdyb[5]/_lv01:13 4.254E-18
C36732  Xa2s_dout[20]/_clk:4    clk:3718 5.128E-19
C36733  Xdll/d:5921     Xdll/Xphased[3]/Xdunit[4][7]/n[1]:3 1.621E-17
C36734  Vdd!    Xdll/Xphased_fclk[1]/n[3][0]:4 2.758E-15
C37065  chan_dll.rden:32        Xdll/Xctrl/Xmux_r[0]/_insel[1]:1
+	 7.851E-17
C37066  Xa2s_dout[20]/clk0:35   dout[22].0:6 1.656E-16
C37067  odq[11]:26      odq[11]:32 1.889E-17
C38712  Xopctrl.opreg[4]/Xolatch/Xlatchv/s:7    Vdd! 8.354E-17
C38713  Xa2s_dout[20]/17:3      Xa2s_dout[20]/15:7 1.077E-16
C38714  Xdll/Xphased_fclk[5]/Xdunit[1][6]/n[0]:4        Xdll/d:4614
+	 2.455E-17
C39180  Xa2s_dout[1]/Rv:11      Xa2s_dout[1]/_R.1:30 7.246E-17
C39181  Xa2s_dout[20]/clk0:36   clk:4720 7.423E-18
C39182  Xopctrl.opreg[1]/Xolatch/Xlatchv/_l:6   Vdd! 8.330E-17
C39187  Xdll/Xphased_fclk[6]/Xdemux/demux._R[0]:2       GND! 1.682E-17
C39188  _SReset!:3269   Xopctrl.A2Sop/Lc[2][15].e:14 4.275E-18
C39189  _PReset!:5973   Xa2s_dout[20]/_R.0:12 3.218E-17
C39190  Xconfigure.a2s/Xdyb[1]/_x[1].0:2        GND! 2.234E-16
C39191  CL[3]:15        CL[3]:14 1.846E-18
C39612  Xophold[13]/Xilatch/Xlatchv/_v:32       
+	Xophold[13]/Xilatch/Xlatchv/_v:31 1.373E-18
C39613  Xa2s_dout[20]/_grant:1  GND! 1.826E-16
C39614  _SReset!:410    Xconfigure.a2s/XcpyRl0/_be_01:5 5.473E-18
C39615  chan_dll.ampsel[3]:2    Xdll/dclk[4]:239 9.884E-17
C39844  Xlatency_ctrl.ieD/X_vdelay[3]/Xnlatch/_clk:19   
+	Xlatency_ctrl.ieD/x[3]:79 3.353E-18
C39845  Xa2s_dout[20]/Rc:10     Xa2s_dout[20]/_R.0:25 3.378E-17
C39846  Xdll/d:6330     Xdll/Xphased_fclk[5]/Xdunit[3][6]/0 1.271E-18
C39847  op4[7].e:24     op4[6].1:8 1.047E-17
C40358  Xopctrl.A2Sop/Xdyb[12]/_x[1].0:8        
+	Xopctrl.A2Sop/Xdyb[12]/35:5 9.493E-17
C40359  Xa2s_dout[20]/29:2      Xa2s_dout[20]/clk0:14 9.723E-18
C40360  dout[12].e:5    dout[12].e:4 1.237E-17
C40361  _PReset!:5384   clk:2416 7.056E-17
C40510  Xa2s_dout[4]/_R.0:33    Xa2s_dout[4]/clk0:24 4.797E-18
C40511  Xa2s_dout[20]/_grant:5  Xa2s_dout[20]/31:1 1.444E-17
C40512  Xopctrl.opreg[8]/Xolatch/Xlatchv/l:1    
+	Xopctrl.opreg[8]/Xolatch/Xlatchv/l:5 3.000E-20
C40880  Xopctrl.opreg[15]/Xolatch/Xlatchv/4:1   GND! 2.090E-16
C40881  Xlatency_ctrl.ieD/x[4]:38       CL[1]:1 1.484E-17
C40882  Xa2s_dout[20]/_clk:32   Xa2s_dout[20]/clk0:35 7.336E-18
C40883  Xopctrl.A2Sop/XbufL[14][0]/12:1 _SReset!:2160 2.037E-18
C41463  Xdll/Xctrl/lcnt[1]:17   
+	Xdll/Xctrl/Xcounter_lock/Xincbit[1]/and._R:10 7.226E-19
C41464  Xa2s_dout[20]/6:3       Xa2s_dout[20]/6:6 3.244E-17
C41465  Xopctrl.rdwr_ctrl/Xbl_counter/maxL[0]:2 
+	Xopctrl.rdwr_ctrl/Xbl_counter/maxL[1]:12 7.206E-18
C42056  Xs2a_din[25]/_Rv:2      Xs2a_din[25]/3:4 1.198E-17
C42057  Xopconv[5]/_r.1:3       Xopconv[5]/4 9.048E-18
C42058  clk:4579        Xa2s_dout[20]/_clk0:14 5.697E-17
C42059  Xconfigure.a2s/XcpyRl1[0]/_be_01:8      
+	Xconfigure.a2s/Lc[2][1].e:26 1.692E-18
C42126  Xdll/Xctrl/Xcounter/Xgl4/_gg1:20        
+	Xdll/Xctrl/Xcounter/Xgl4/_A[1]:2 3.718E-18
C42127  Xa2s_dout[20]/_clk:3    Xa2s_dout[20]/_clk0:9 1.346E-17
C42128  Xopctrl.rdwr_ctrl/Xbl_counter/maxL[7]:9 
+	Xopctrl.rdwr_ctrl/Xbl_counter/maxL[7]:8 5.710E-17
C42581  Xconfigure.a2s/XcL/Lc[5].e:26   Xconfigure.a2s/XcL/LD[4].e:25
+	 3.349E-18
C42582  Xa2s_dout[20]/0:5       Xa2s_dout[20]/0:1 3.377E-18
C42583  _SReset!:3823   GND! 6.755E-16
C42928  Vdd!    Xdll/Xphased[0]/Xdunit[4][9]/n[1]:1 2.066E-16
C42929  Xopctrl.opreg[14]/Xolatch/Xlatchv/_out:5        GND! 1.237E-16
C42930  Xa2s_dout[20]/7:3       Xa2s_dout[20]/__Le:10 7.245E-17
C42931  GND!    Xconfigure.a2s/XcpyRl0/_be_01:15 9.548E-18
C44065  Xopctrl.opreg[22]/_clk:13       
+	Xopctrl.opreg[22]/Xolatch/Xlatchv/_out:16 2.873E-18
C44066  Xa2s_dout[20]/9:3       GND! 1.498E-16
C44067  Xinit_wait.dffinc0/Xdelay/Xdelay[2]/x:1 
+	Xinit_wait.dffinc0/Xdelay/Xdelay[2]/x:10 7.932E-19
C44106  sop[0][4]:24    Vdd! 6.409E-16
C44107  Xa2s_dout[20]/_clk:1    Xa2s_dout[20]/clk0:6 5.781E-17
C44108  Xdll/d:5922     Vdd! 2.427E-18
C44463  Xinit_wait.cntr0/Xincbit0/Xtreg/Xilatch/l:1     
+	Xinit_wait.cntr0/Xincbit0/Xtreg/Xilatch/10 4.734E-18
C44464  Xa2s_dout[20]/21:1      Xa2s_dout[20]/15:4 4.794E-18
C44465  Xa2s_dout[23]/_R.0:28   clk:4702 5.722E-17
C44751  Vdd!    Xdll/d:5944 1.057E-17
C44752  Xa2s_dout[20]/_R.1:4    Xa2s_dout[20]/_clk:1 5.735E-19
C44753  Xlatency_ctrl.ieD/Xvdelay[0]/Xplatch/Xlatchv/_l:10      
+	Xlatency_ctrl.ieD/Xvdelay[0]/Xplatch/Xlatchv/_out:31 6.427E-19
C45476  Xconfigure.a2s/XcL/Lc[6].e:15   
+	Xconfigure.a2s/XcL/XcpyL[6]/Xc01/_c:25 3.570E-17
C45477  Xa2s_dout[20]/_clk0:18  Xa2s_dout[20]/_noR:29 2.753E-17
C45478  Xa2s_dout[0]/9:3        GND! 1.515E-16
+	Xinit_wait.cntr0/Xincbit[5]/d:14 1.103E-17
C46259  Vdd!    Xinit_wait.cntr0/Xincbit[4]/xnor._L[0]:7 1.344E-16
C46260  Xa2s_dout[20]/_clk0:2   Xa2s_dout[20]/1:2 2.282E-16
C46261  GND!    Xopctrl.opreg[20]/Xilatch/_v:25 5.726E-17
C46262  Xdll/d:5994     Vdd! 7.762E-18
C46326  Xa2s_dout[20]/_noR:14   Xa2s_dout[20]/_noR:26 9.431E-18
C46327  _PReset!:3747   Xopctrl.A2Sop/Xdyb[13]/2 9.572E-19
C46328  Xa2s_dout[27]/Rc:9      GND! 1.810E-16
C46589  Xa2s_dout[20]/_noR:14   Xa2s_dout[20]/0:3 1.792E-17
C46590  Xopctrl.A2Sop/XbufL[14][0]/be:22        _PReset!:2627
+	 1.608E-19
C46761  clk:4028        Xa2s_dout[20]/_clk0:14 2.410E-17
C46762  Xa2s_dout[21]/Rc:9      GND! 1.810E-16
C46763  _SReset!:997    _SReset!:888 2.276E-17
C46838  Xdqsgen[1]/Xa2s_odqs/_R.1:28    clk:2045 1.018E-17
C46839  Xa2s_dout[20]/Rc:9      GND! 1.810E-16
C46840  Xopctrl.nopctrl/Xnopcntr/Xcounter/inc[3]:3      _SReset!:1266
+	 4.462E-17
C47361  Xopctrl.opreg[24]/_clk:11       
+	Xopctrl.opreg[24]/Xolatch/Xlatchv/_in:8 3.809E-18
C47362  Xa2s_dout[20]/_clk0:39  dout[22].0:4 3.294E-18
C47363  Xdqsgen[2]/Xalt_dqs/x.1:26      Xdqsgen[2]/Xalt_dqs/x.1:13
+	 1.006E-18
C47391  Xconfigure.a2s/Xdyb[11]/35:7    Vdd! 3.305E-17
C47392  Xinit_wait.cntr0/Xincbit[6]/and._R:4    Vdd! 2.379E-16
C47393  odq[20]:4       Xa2s_dout[20]/_r:17 2.609E-17
C47394  Vdd!    Xopctrl.rdwr_ctrl/Xbl_counter/cnt[5]:19 1.674E-16
C47965  _PReset!:240    _PReset!:257 1.194E-19
C47966  Vdd!    config[5].0 7.750E-17
C47967  Xa2s_dout[20]/_clk:21   Xa2s_dout[20]/PReset:4 3.397E-17
C47968  sop[0][12]:3    Xopctrl.opmux[16]/_insel[1]:5 2.176E-18
C48783  Xopconv[11]/_r.0:11     Xopconv[11]/_r.1:11 1.723E-17
C48784  Xdll/d:1315     GND! 5.760E-15
C48785  Xa2s_dout[20]/_clk:1    Xa2s_dout[20]/_r:16 3.521E-17
C48786  Xopctrl.A2Sop/XcL/XdetectL[9]/__Le:7    GND! 2.395E-16
C48787  Vdd!    Xdll/Xctrl/lcnt[1]:9 3.738E-18
C49239  Xopctrl.opreg[5]/Xolatch/Xlatchv/s:6    
+	Xopctrl.opreg[5]/Xolatch/Xlatchv/s:4 1.702E-17
C49240  Xa2s_dout[20]/8:3       GND! 1.909E-16
C49241  Xlatency_ctrl.ieD/Xvdelay[0]/Xplatch/Xlatchv/_v:19      
+	Xlatency_ctrl.ieD/Xvdelay[0]/Xplatch/Xlatchv/_v:14 3.596E-18
C49653  Xdll/Xctrl/Xcounter_lock/Xincbit0/Xtreg/Xilatch/v:1     
+	Xdll/Xctrl/Xcounter_lock/Xincbit0/Xtreg/Xilatch/v:5 6.321E-19
C49654  Xa2s_dout[20]/Rv:2      Xa2s_dout[20]/7:2 7.712E-19
C49655  Xdll/Xphased_fclk[3]/Xdunit[1][1]/n[0]:7        Xdll/d:4224
+	 2.642E-19
C49976  Xdll/Xphased[3]/Xdunit[2][8]/n[0]:1     
+	Xdll/Xphased[3]/Xdunit[2][8]/n[0]:3 5.380E-18
C49977  Xa2s_dout[20]/_r:2      odq[20]:12 5.209E-17
C49978  Xa2s_dout[14]/_clk:1    clk:3566 2.209E-17
C49979  Xopctrl.A2Sop/XcL/XdetectL[2]/__Le:4    GND! 3.062E-16
+	 3.061E-17
C50513  Vdd!    Xconfigure.a2s/Xdyb[4]/_x[1].1:16 9.027E-17
C50514  Xa2s_dout[20]/_clk:1    _SReset!:5109 1.519E-17
C50515  Xconfigure.a2s/Xctrl/Xglatch/_r.0:11    
+	Xconfigure.a2s/Xctrl/Xglatch/s:16 6.333E-18
C50798  Xconfigure.a2s/XcpyRl1[2]/Xc23/8:5      
+	Xconfigure.a2s/XcpyRl1[2]/_be_23:16 1.472E-17
C50799  Xa2s_dout[20]/_clk:1    Xa2s_dout[20]/_noR:21 5.525E-17
C50800  sop[0][19]:7    Xopctrl.opreg[23]/_clk:10 4.486E-18
C50801  Xdll/Xphased_fclk[5]/n[7][2]:7  Xdll/d:3838 3.108E-20
C51635  CL[3]   Xconfigure.a2s/XbufRl0/_rd:32 2.568E-18
C51636  opctrl.xop[1][1]:27     Xopctrl.opreg[1]/x:7 1.531E-16
C51637  Xa2s_dout[20]/_r:6      Xa2s_dout[20]/_r:3 1.846E-18
C51638  _PReset!:519    Xconfigure.a2s/Xdyb[2]/51 4.002E-18
C51639  Xconfigure.a2s/Lv[1].e:8        GND! 2.716E-16
C52179  Xconfigure.a2s/Lc[2][4].0:5     Xconfigure.a2s/cRl[2][1].0:38
+	 4.336E-18
C52180  Xa2s_dout[20]/clk0:7    clk:4579 2.062E-16
C52181  dout[24].1:1    Xa2s_dout[22]/Rv:8 2.134E-17
C52795  Xdll/Xphased[3]/Xdunit[1][4]/n[1]:3     
+	Xdll/Xphased[3]/Xdunit[1][4]/n[0]:7 3.056E-17
C52796  Xa2s_dout[20]/6:5       Xa2s_dout[20]/6:1 6.019E-18
C52797  Xdll/Xctrl/lrst:11      
+	Xdll/Xctrl/Xcounter_lock/Xincbit[3]/0:2 1.203E-18
C53112  Xdll/r.0:92     Xdll/r.0:98 3.088E-18
C53113  Vdd!    Xdll/Xphased[1]/Xdunit[4][6]/n[0]:1 2.434E-16
C53114  Xa2s_dout[20]/_noR:24   Xa2s_dout[20]/_noR:17 5.979E-18
C53115  Xa2s_dout[9]/_R.1:27    clk:4624 3.401E-17
C53116  Xconfigure.a2s/XbufL[11][0]/_b.0:2      _SReset!:681 1.062E-17
C53277  Xdll/Xgate_dclk2/Den:1  Xdll/Xgate_dclk2/Xarb/_D[0]:14
+	 2.637E-17
C53278  Xa2s_dout[20]/10:3      dout[22].0:6 4.876E-18
C53279  op2[13].1:4     op2[13].0:14 1.209E-17
C53775  Xdll/r.4:192    Xdll/Xphased_fclk[3]/n[3][7]:5 2.675E-18
C53776  Vdd!    Xdll/Xphased[0]/Xdunit[3][8]/n[0]:1 2.434E-16
C53777  Xa2s_dout[20]/clk0:29   Xa2s_dout[20]/_clk0:40 1.207E-17
C53778  Xdll/Xphased[0]/n[0][11]:5      Xdll/r.0:110 5.398E-18
C53779  Xa2s_dm[0]/_Le:13       GND! 6.304E-17
C54381  GND!    Xophold[13]/Xolatch/Xlatchv/PReset:14 6.218E-17
C54382  Xopctrl.A2Sop/XcL/Lc[8].e:28    Vdd! 8.338E-16
C54383  Xa2s_dout[20]/7:4       Xa2s_dout[20]/__Le:4 1.225E-16
C54384  Xconfigure.a2s/Xdyb[6]/rvb[0]:15        
+	Xconfigure.a2s/Xdyb[6]/_x[0].0:18 3.082E-18
C54825  Xa2s_dout[20]/_clk0:15  GND! 2.637E-16
C54826  Xopctrl.opreg[17]/Xilatch/_v:1  _SReset!:3868 3.441E-16
C54827  Xopctrl.opreg[12]/Xilatch/_out:10       GND! 2.619E-17
C55729  Xdll/Xphased_fclk[6]/n[2][4]:7  GND! 1.613E-16
C55730  _PReset!:3410   avC814:14 8.746E-18
C55731  Xa2s_dout[20]/_clk0:54  Xa2s_dout[20]/_R.0:33 4.250E-18
C55732  Xdll/r.1:105    Xdll/Xphased_fclk[0]/n[1][1]:5 3.290E-18
C55770  opctrl.xop[1][7]:24     Xopctrl.opreg[7]/Xilatch/l:6 4.281E-18
C55771  _SReset!:1454   Xopctrl.A2Sop/XcL/XdetectL[8]/_R:14 2.116E-18
C55772  clk:3618        Xa2s_dout[20]/_clk:4 4.869E-19
C55773  Xopctrl.A2Sop/Lc[2][1].0:18     Xopctrl.A2Sop/Lc[2][1].1:9
+	 4.567E-17
C56252  Xdll/Xphased[3]/n[1][0]:1       Xdll/d:4183 7.612E-18
C56253  _SReset!:5458   Xa2s_dout[20]/16 1.078E-18
C56254  Xdll/Xphased_fclk[6]/n[2][0]:11 GND! 1.624E-16
C56621  Xdll/Xphased_fclk[7]/n[2][12]:5 
+	Xdll/Xphased_fclk[7]/Xdunit[2][12]/n[1]:1 3.875E-19
C56622  Xa2s_dout[20]/29:2      Xa2s_dout[20]/clk0:37 4.272E-18
C56623  Xopctrl.opreg[5]/Xilatch/_out:6 
+	Xopctrl.opreg[5]/Xilatch/_out:22 3.288E-19
C58251  _SReset!:1407   GND! 2.379E-16
C58252  clk:4581        Xa2s_dout[20]/_r:16 1.817E-16
C58253  Xconfigure.a2s/Xctrl/PReset:10  GND! 1.558E-16
C58306  Xa2s_dout[4]/_Le:3      clk:3734 2.773E-17
C58307  Xa2s_dout[20]/26:1      Xa2s_dout[20]/PReset:6 5.437E-18
C58308  invdq[0].R:18   Xinvdq[0]/x:21 1.063E-17
C58423  Xconfigure.a2s/XcL/LD4[0].e:9   
+	Xconfigure.a2s/XcL/XdetectLD[0]/_R:14 1.396E-16
C58424  Xa2s_dout[20]/51:2      Xa2s_dout[20]/clk0:11 1.591E-17
C58425  Vdd!    Xdll/d:5100 1.031E-17
C58426  sop[1][14]:6    clk:3123 3.951E-17
C59437  sop[0][11]:47   sop[0][11]:38 4.731E-17
C59438  _PReset!:6732   Xa2s_dout[20]/PReset:4 8.571E-18
C59439  Xconfigure.a2s/Lc[2][4].3:15    GND! 4.607E-17
C59440  Vdd!    Xconfigure.a2s/Lc[2][7].2:4 5.733E-18
C74124  _PReset!:3551   Xdll/Xctrl/Xalt_r/alt.x[0].0:28 3.252E-18
C74125  clk:709 Xopctrl.A2Sop/Xdyb[11]/13:4 4.566E-17
C74126  Xa2s_dout[20]/__Le:2    Xa2s_dout[20]/_R.0:23 1.001E-19
C74127  Xdll/r.3:193    Xdll/Xphased_fclk[7]/n[3][11]:5 2.667E-18
C75466  GND!    Xdll/Xphased_fclk[1]/Xmux/sl4[0]:1 1.361E-16
C75467  Xa2s_dout[20]/_R.0:34   GND! 7.199E-17
C75468  Xdll/d:3741     Xdll/Xphased[2]/Xdunit0[3]/n[0]:2 7.309E-17
C75469  Xopctrl.A2Sop/XcL/XdetectL[7]/_L01v:5   Vdd! 2.083E-17
C86568  Xopctrl.A2Sop/Xdyb[6]/32:13     
+	Xopctrl.A2Sop/Xdyb[6]/_x[0].1:6 2.018E-17
C86569  _PReset!:6825   Xa2s_dout[20]/_R.0:27 7.671E-19
C86570  opctrl.xop[1][24]:10    GND! 2.013E-16
C90772  NRFRSH[1]:16    Xrefresh_gen.xnor[1]/_L[1]:5 1.117E-16
C90773  Xopctrl.opreg[0]/Xilatch/v:2    GND! 1.837E-16
C90774  Vdd!    Xa2s_dout[20]/_R.0:3 4.318E-18
C106439 Xopctrl.A2Sop/Lc[2][11].3:24    Xopctrl.A2Sop/Lc[2][11].0:21
+	 2.161E-17
C106440 Vdd!    Xa2s_dout[20]/_R.0:29 7.573E-18
C106441 Xopctrl.A2Sop/XcpyRl1[0]/Xc03/8:5       
+	Xopctrl.A2Sop/cRl[2][0].e:4 1.472E-17
C114625 Xconfigure.a2s/XcL/LD[2].0:14   
+	Xconfigure.a2s/XcL/XdetectLD[0]/29 5.385E-18
C114626 Xa2s_dout[20]/_R.1:27   Xa2s_dout[20]/_R.0:17 4.240E-18
C116495 Xopctrl.A2Sop/XcpyRl0/_be_23:6  Xopctrl.A2Sop/cRl[1][3].e:10
+	 1.158E-18
C116496 Xa2s_dout[20]/Rc:4      Xa2s_dout[20]/_R.0:20 6.139E-18
C118160 GND!    Xa2s_dout[20]/_R.0:29 2.056E-17
C118161 Xs2a_din[14]/go:27      Xs2a_din[14]/xnor._L[1]:5 5.205E-18
C119353 Xa2s_dout[20]/_R.0:18   Xa2s_dout[20]/0:5 4.549E-17
C119354 _ddqs[1]:13     Xdll/Xphased_fclk[2]/Xmux/_sl[3]:5 3.017E-18
C121854 Xdll/Xphased_fclk[1]/n[2][4]:7  Xdll/d:5572 1.368E-19
C121855 Xa2s_dout[10]/_R.0:19   Xa2s_dout[10]/_noR:12 2.453E-17
C121856 Xa2s_dout[20]/_R.0:16   odq[20]:19 5.754E-18
C121857 Xopctrl.A2Sop/XbufL[11][0]/_b.0:10      
+	Xopctrl.A2Sop/Lc[0][11].e:20 2.442E-17
C127287 Xdll/Xphased[0]/n[3][2]:4       Xdll/d:2749 2.049E-18
C127288 _SReset!:2323   _SReset!:2029 7.618E-18
C127289 Xa2s_dout[20]/_R.0:6    Xa2s_dout[20]/_R.1:15 5.477E-18
C127290 Xinit_wait.cntr0/Xincbit[4]/Xreg/Xlatch/Xlatchv/_out:4  
+	_PReset!:5545 5.206E-17
C132299 _PReset!:3818   Xdll/Xctrl/Xalt_r/184:1 6.767E-18
C132300 Xa2s_dout[20]/_R.0:35   Vdd! 1.354E-16
C132301 Xrefresh_gen.inc1/Xincbit[3]/Xreg/Xlatch/Xlatchv/v:1    
+	clk:3750 5.301E-17
C134696 Vdd!    Xs2a_din[22]/Rv:6 1.959E-17
C134697 Xa2s_dout[20]/_R.1:32   Xa2s_dout[20]/_R.0:17 2.828E-17
C134698 Xopctrl.A2Sop/XbufL[2][0]/12:3  _SReset!:2208 2.640E-17
C136175 Xa2s_dout[20]/_R.0:11   odq[20]:17 2.793E-17
C136176 Xinit_wait.cntr0/Xincbit[1]/Xreg/Xlatch/Xlatchv/PReset:9
+	Xinit_wait.cntr0/Xincbit[1]/d:39 3.327E-16
C139535 Xa2s_dout[20]/_grant:2  Xa2s_dout[20]/_R.0:27 1.550E-18
C139536 Xopctrl.A2Sop/Lc[1][4].e:2      
+	Xopctrl.A2Sop/XbufL[4][0]/_ae:14 1.397E-18
C139661 Xa2s_dout[20]/_R.0:21   _PReset!:6361 3.299E-18
C139662 Xdll/Xctrl/Xcounter_lock/Xincbit[2]/Xreg/Xdelay/Xdelay[0]/x:3
+	Xdll/Xctrl/Xcounter_lock/inc[2]:30 7.709E-18
C139811 _SReset!:5446   Xa2s_dout[29]/17:1 2.313E-17
C139812 Xa2s_dout[20]/_R.0:9    clk:3554 1.921E-16
C139813 opctrl.xop[0][3]:2      Xopctrl.A2Sop/Xdyb[1]/_R[1]:21
+	 3.692E-17
C144466 Xopctrl.A2Sop/Xdyb[2]/_x[0].0:15        
+	Xopctrl.A2Sop/Xdyb[2]/r[0].0:13 4.754E-18
C144467 Xa2s_dout[20]/_R.0:26   clk:4493 9.847E-18
C144468 _PReset!:4069   Xdll/dllen:24 3.775E-16
C145870 Xa2s_dout[20]/10:6      Xa2s_dout[20]/_R.0:34 1.579E-17
C164288 Xa2s_dout[8]/_clk:22    clk:4777 2.989E-18
C164289 _SReset!:843    CL[3] 1.019E-16
C164290 Xa2s_dout[20]/_R.0:24   Xa2s_dout[20]/_clk:33 2.350E-18
C171688 _PReset!:6825   Xa2s_dout[20]/_R.0:35 1.955E-17
C171689 Xdll/Xphased_fclk[7]/Xdunit[3][6]/n[1]:4        
+	Xdll/Xphased_fclk[7]/n[3][7]:4 8.823E-17
C172924 Xa2s_dout[20]/_R.0:28   Xa2s_dout[20]/21:3 1.525E-17
C172925 Xlatency_ctrl.oeH/Xdelay/Xlatch[0]/Xlatchv/v:10 
+	Xlatency_ctrl.oeH/Xdelay/Xlatch[0]/Xlatchv/_v:10 4.825E-17
C173561 Xa2s_dout[20]/_R.0:23   odq[20]:13 4.647E-18
C173562 Xrefresh_gen.inc0/Xincbit[4]/d:4        
+	Xrefresh_gen.inc0/Xincbit[4]/__rst:8 2.632E-17
C186160 Xa2s_dout[20]/_R.0:6    Xa2s_dout[20]/Rc:10 1.601E-16
C186161 opctrl.xop[0][12]:3     Xopctrl.A2Sop/Xdyb[6]/r[0].0:14
+	 2.207E-18
C187757 Xa2s_dout[20]/_R.0:3    Xa2s_dout[20]/_R.1:14 5.075E-17
C187758 op4[2].1:5      _PReset!:1411 6.516E-19
C192627 Xa2s_dout[20]/_R.0:11   GND! 5.783E-16
C192628 Xs2a_din[23]/_clk0:20   Vdd! 3.311E-16
C192629 Xopctrl.A2Sop/Xdyb[11]/_clk:10  GND! 1.134E-16
C192682 Xdll/r.7:78     Xdll/dclk[2]:14 5.791E-19
C192683 Xdll/Xphased[1]/Xmux/_sl[5]:2   Vdd! 2.689E-16
C192684 Xa2s_dout[20]/_R.0:12   GND! 3.041E-16
C192685 Xopctrl.A2Sop/Xdyb[10]/_clk:11  GND! 1.280E-16
C192686 Xdll/dclk[0]:69 chan_dll.dpass:5 3.549E-17
C197589 Xa2s_dout[20]/_R.0:14   Xa2s_dout[20]/2 2.251E-18
C197590 Xa2s_dm[1]/1:1  Xa2s_dm[1]/0:7 3.556E-17
C198857 clk:4581        Xa2s_dout[20]/_R.0:11 4.023E-17
C198858 GND!    Xopctrl.opreg[27]/Xilatch/_v:33 2.938E-18
C198859 _SReset!:127    Xconfigure.a2s/Xctrl/_done:2 1.531E-18
C202824 Xa2s_dout[20]/_R.0:30   dout[22].0:1 6.533E-19
C213588 Xa2s_dout[20]/_R.0:14   odq[20]:19 8.446E-18
C213589 Xopctrl.A2Sop/XbufL[0][1]/12:4  
+	Xopctrl.A2Sop/XbufL[0][1]/_b.0:4 1.574E-17
C215005 Xa2s_dout[20]/_R.0:11   clk:3799 2.577E-18
C215006 Xs2a_din[5]/xnor._L[0]:13       Xs2a_din[5]/_clk0:20 3.370E-18
C218555 Xa2s_dout[20]/_R.0:28   clk:4717 5.722E-17
C218556 Xa2s_dout[8]/clk0:5     Xa2s_dout[8]/_clk:21 5.591E-17
C221363 Xa2s_dout[20]/_R.0:16   GND! 3.079E-17
C222501 Xa2s_dout[20]/_R.0:33   Vdd! 1.171E-16
C226480 Xa2s_dout[20]/_clk0:46  Xa2s_dout[20]/_R.0:35 3.065E-18
C232103 Xa2s_dout[20]/_R.0:30   GND! 8.438E-17
C245799 Xa2s_dout[20]/_R.0:31   Xa2s_dout[20]/_R.0:33 3.916E-18
C245800 Xopctrl.A2Sop/Lv[0].0:16        op4[3].3:30 5.576E-16
C253614 Xa2s_dout[20]/_R.0:33   Xa2s_dout[20]/_R.0:35 1.034E-18
C257597 Xa2s_dout[20]/_R.1:15   Xa2s_dout[20]/_R.0:19 2.142E-17
C284238 Xa2s_dout[20]/_R.0:30   Xa2s_dout[20]/10:4 1.481E-17
C284239 Xrefresh_gen.s2a/Xctrl/_go:1    Xrefresh_gen.s2a/go:4
+	 6.956E-19
C287297 Xa2s_dout[20]/_R.0:27   Xa2s_dout[20]/_clk0:38 5.561E-18
C287528 Xa2s_dout[20]/_R.0:24   Xa2s_dout[20]/_R.0:25 2.181E-17
C287529 Xdll/Xphased_fclk[0]/Xdunit[4][0]/n[1]:7        
+	Xdll/Xphased_fclk[0]/n[4][1]:4 2.096E-17
C287967 Xa2s_dout[20]/_R.1:28   Xa2s_dout[20]/_R.0:11 6.037E-17
C290328 Xa2s_dout[20]/10:5      Xa2s_dout[20]/_R.0:31 1.655E-17
C292554 Xa2s_dout[20]/__Le:3    Xa2s_dout[20]/_R.0:23 5.283E-20
C301775 dout[22].0:4    Xa2s_dout[20]/_R.0:29 8.630E-18
C302114 Xa2s_dout[20]/_R.0:25   _PReset!:6825 2.275E-18
C309738 Xa2s_dout[20]/_R.0:1    Xa2s_dout[20]/_R.1:13 4.764E-19
C314876 Xa2s_dout[20]/_R.0:24   dout[22].0:2 1.166E-17
C318306 Xa2s_dout[20]/Rv:1      Xa2s_dout[20]/_R.0:23 5.542E-20
C319151 Xa2s_dout[20]/_R.0:34   Xa2s_dout[20]/clk0:23 4.798E-18
C326682 dout[22].0:2    Xa2s_dout[20]/_R.0:25 6.000E-17
C335647 Xa2s_dout[20]/_r:13     Xa2s_dout[20]/_R.0:23 6.965E-17
C338618 Xa2s_dout[20]/_R.0:33   Xa2s_dout[20]/clk0:24 4.797E-18
C343284 Xa2s_dout[20]/_R.0:26   Xa2s_dout[20]/_R.0:25 7.203E-17
C344250 Xa2s_dout[20]/10:3      Xa2s_dout[20]/_R.0:34 7.588E-17
C345254 clk:3618        Xa2s_dout[20]/_R.0:11 5.932E-17
C347109 Xa2s_dout[20]/21:2      Xa2s_dout[20]/_R.0:29 1.655E-16
C350769 Xa2s_dout[20]/_R.0:16   odq[20]:22 2.124E-16
C354085 _PReset!:6164   Xa2s_dout[20]/_R.0:21 1.596E-17
C354437 _SReset!:5270   Xa2s_dout[20]/_R.0:12 1.460E-17
C357223 Xa2s_dout[20]/_R.0:18   Xa2s_dout[20]/_noR:17 9.708E-18
C360392 Xa2s_dout[20]/_R.0:19   Xa2s_dout[20]/_noR:11 4.811E-17
C361909 Xa2s_dout[20]/_R.0:13   odq[20]:19 4.508E-17
C367177 Xa2s_dout[20]/_R.0:27   GND! 5.130E-16
C367252 Xa2s_dout[20]/_R.0:24   GND! 1.899E-16
C379447 Xa2s_dout[20]/__Le:10   Xa2s_dout[20]/_R.0:11 8.092E-18
C381039 Xa2s_dout[20]/_R.0:28   GND! 5.926E-17
C382003 Xa2s_dout[20]/_R.0:1    odq[20]:4 1.850E-16
C382628 Xa2s_dout[20]/_R.0:26   GND! 5.497E-16
C382629 _SReset!:1435   Xopctrl.A2Sop/XcL/XcpyL[15]/Xc01/_c:15
+	 2.732E-17
C383137 Xa2s_dout[20]/_R.1:39   Xa2s_dout[20]/9:5 5.038E-18
C383138 Xdll/Xctrl/Xalt_r/alt.yv[1]:3   
+	Xdll/Xctrl/Xalt_r/alt._y[2].1:9 1.365E-17
C383913 _SReset!:1206   op2[3].0:7 6.634E-18
C383914 Xa2s_dout[20]/PReset:3  GND! 1.211E-16
C383915 Xopctrl.A2Sop/Lc[2][9].1:25     GND! 1.354E-16
C383916 Xophold[19]/Xilatch/Xlatchv/v:1 sop[0][19]:54 1.427E-17
C383977 opctrl.xop[1][3]:17     Vdd! 3.123E-16
C383978 Xdll/Xctrl/Xalt_r/alt.yv[1]:1   Vdd! 9.646E-16
C383979 Xa2s_dout[20]/PReset:5  GND! 2.153E-16
C383980 Xdll/r.0:117    Xdll/Xphased_fclk[6]/Xdunit0[2]/n[0]:9
+	 2.949E-18
C384316 Xophold[16]/Xolatch/Xlatchv/_in:5       
+	Xophold[16]/Xolatch/Xlatchv/_out:23 2.389E-18
C384317 Xa2s_dout[20]/21:3      Xa2s_dout[20]/clk0:32 9.083E-18
C384318 Xopctrl.A2Sop/XbufLv[3]/_rd:8   Xopctrl.A2Sop/Lv[4].e:46
+	 6.455E-17
C384715 Xrefresh_gen.s2a/Xbufx[1]/be:8  Xrefresh_gen.s2a/Rg[0].0:17
+	 1.084E-16
C384716 clk:3491        Xa2s_dout[20]/_r:3 9.017E-18
C384717 Xconfigure.a2s/Lc[1][0].0:19    Xconfigure.a2s/Lc[1][0].1:8
+	 6.216E-17
C385283 Xophold[13]/Xolatch/Xlatchv/5:6 
+	Xophold[13]/Xolatch/Xlatchv/_out:4 1.037E-17
C385284 Xa2s_dout[20]/_noR:12   Xa2s_dout[20]/_noR:4 3.681E-19
C385285 Xconfigure.a2s/Lc[0][7].e:19    
+	Xconfigure.a2s/Xdyb[8]/_x[0].1:23 1.540E-18
C385375 Vdd!    op4[11].1:2 1.368E-17
C385376 _PReset!:5720   Xophold[12]/Xolatch/Xlatchv/_in:15 9.278E-18
C385377 Xa2s_dout[20]/8:3       Xa2s_dout[20]/_R.1:41 7.940E-17
C385378 Xconfigure.a2s/XbufL[7][1]/_b.3:6       
+	Xconfigure.a2s/Lc[2][7].3:21 3.221E-19
C385646 clk:1221        Vdd! 2.148E-16
C385647 Xa2s_dout[20]/_R.0:5    _SReset!:5034 4.932E-18
C385648 Xdll/d:2056     Xdll/Xphased_fclk[0]/n[5][4]:4 4.852E-22
C385649 Xopctrl.A2Sop/Lc[2][7].0:18     Vdd! 4.088E-17
C385684 Xa2s_dout[20]/_clk0:27  GND! 2.194E-16
C385685 odq[26]:4       Xa2s_dout[26]/_R.1:19 6.009E-17
C385897 Xdll/d:5082     Xdll/Xphased_fclk[5]/Xdunit[2][11]/n[0]:6
+	 3.242E-18
C385898 Xa2s_dout[20]/_clk:20   Xa2s_dout[20]/_clk:19 6.071E-17
C385899 Xopctrl.A2Sop/Lc[2][5].0:18     Vdd! 4.954E-17
C385900 op4[8].2:2      Vdd! 8.647E-18
C386701 Xa2s_dout[20]/_r:13     Xa2s_dout[20]/_R.0:22 1.331E-17
C386702 Xinit_wait.cntr1/Xincbit[5]/Xreg/Xlatch/Xlatchv/_out:35 GND!
+	 2.636E-16
C386820 Xopctrl.A2Sop/Lc[2][3].e:54     Xopctrl.A2Sop/Lc[2][3].2:34
+	 2.743E-16
C386821 clk:3491        Xa2s_dout[20]/_R.0:23 1.058E-17
C386858 avC792:22       avC792:17 3.707E-17
C386859 Xdll/r.1:202    Xdll/d:5083 1.855E-16
C386860 Xa2s_dout[20]/6:6       Xa2s_dout[20]/_noR:1 2.038E-19
C387207 Xdll/Xphased[1]/n[1][9]:4       Xdll/r.1:117 6.582E-18
C387208 Xa2s_dout[20]/clk0:8    clk:4341 3.209E-17
C387209 Xs2a_din[1]/1:4 ddqs[0]:15 4.359E-18
C387210 op2[7].0:4      Xopconv[3]/14:1 6.501E-19
C388300 _SReset!:1197   op4[6].e:19 4.200E-18
C388301 Xopconv[6]/_r.0:28      GND! 4.690E-16
C388302 Xa2s_dout[20]/_r:3      odq[20]:4 1.105E-17
C388303 opctrl.nopsel:6 opctrl.nops[3]:20 2.470E-17
C388557 Xa2s_dout[20]/_R.0:9    Xa2s_dout[20]/Rv:14 1.763E-18
C393016 Xa2s_dout[20]/__Le:2    Xa2s_dout[20]/_R.0:22 3.042E-21
C393017 Xdqsgen[0]/Xalt_dqs/x.1:2       Xdqsgen[0]/Xalt_dqs/_r.1:17
+	 3.644E-17
C402705 Xa2s_dout[20]/10:4      Xa2s_dout[20]/_R.0:33 1.224E-16
C403238 dout[21].1:1    Xa2s_dout[20]/_R.0:26 2.237E-17
C409697 Xa2s_dout[20]/_R.0:31   dout[22].0:1 9.490E-18
C410925 Xa2s_dout[20]/_R.0:11   Vdd! 7.526E-17
C410926 Xopctrl.opreg[8]/_clk:11        GND! 3.271E-17
C410974 Vdd!    Xa2s_dout[20]/_R.0:12 7.080E-17
C436516 Xa2s_dout[20]/_R.0:24   _SReset!:5423 5.299E-17
C436517 Vdd!    Xa2s_dout[31]/_R.1:7 4.067E-17
C440173 Xa2s_dout[20]/_R.0:31   GND! 3.378E-17
C440174 Xdll/Xphased[0]/n[2][12]:4      Xdll/Xphased[0]/n[3][10]:4
+	 5.014E-18
C440376 Xopctrl.opreg[6]/Xolatch/Xlatchv/_out:31        GND! 9.531E-17
C440377 _SReset!:1218   op4[10].e:8 4.066E-17
C440378 Xa2s_dout[20]/Rv:1      odq[20]:13 3.073E-20
C440379 Xopctrl.A2Sop/XbufL[14][1]/_c_01:5      Vdd! 2.235E-16
C440528 Xopctrl.A2Sop/Lc[2][11].e:29    
+	Xopctrl.A2Sop/XcpyRl1[2]/Xc23/8:3 1.702E-17
C440529 Xa2s_dout[20]/_R.0:5    Xa2s_dout[20]/_R.0:4 2.760E-17
C440530 Xrefresh_gen.s2a/x[2].e:10      _SReset!:4815 9.407E-19
C440531 Vdd!    Xopctrl.A2Sop/XcpyRl1[0]/_be_01:55 8.858E-18
C440906 Xdll/Xphased_fclk[3]/Xdunit0[0]/n[0]:7  
+	Xdll/Xphased_fclk[3]/Xdunit0[1]/n[0]:1 6.478E-21
C440907 Xa2s_dout[20]/PReset:3  Xa2s_dout[20]/PReset:4 4.054E-17
C440908 Xconfigure.a2s/XbufL[11][1]/16:3        
+	Xconfigure.a2s/XbufL[11][1]/_b.3:12 1.256E-17
C441134 Xopctrl.A2Sop/XbufL[12][1]/_c_01:5      Vdd! 2.250E-16
C441135 Xophold[3]/Xilatch/Xlatchv/l:6  sop[0][3]:40 3.731E-17
C441136 Xa2s_dout[20]/_R.0:9    clk:3555 6.438E-17
C441137 _PReset!:3094   Xopctrl.A2Sop/XbufL[15][1]/_ae:11 3.524E-18
C441138 Xa2s_dout[15]/26:2      Xa2s_dout[15]/Rc:12 3.381E-18
C441291 Xopconv[3]/_r.1:24      op4[3].1:4 1.201E-17
C441292 GND!    Xdll/Xphased_fclk[0]/Xdunit[1][3]/n[1]:1 1.720E-17
C441293 Xa2s_dout[20]/__Le:8    Vdd! 1.745E-16
C441294 Xdll/d:2575     Xdll/Xphased_fclk[2]/Xdunit[3][0]/0 8.198E-18
C441295 sop[0][16]:64   Xophold[16]/Xilatch/Xlatchv/_in:11 2.284E-18
C441491 Xopctrl.A2Sop/XcpyRl1[2]/_be_01:31      
+	Xopctrl.A2Sop/XcpyRl1[2]/_be_23:35 2.606E-17
C441492 Xa2s_dout[20]/8:1       Xa2s_dout[20]/_R.1:39 2.105E-20
C441493 ie[3]:99        Xs2a_din[16]/1:3 4.594E-20
C441494 Xdll/Xdetect[15]/en_n:4 Xdll/d:7002 1.696E-17
C441999 Xdll/d:3831     Xdll/Xphased_fclk[1]/n[0][1]:6 6.956E-19
C442000 Xa2s_dout[20]/9:2       Xa2s_dout[20]/Rv:10 9.389E-17
C442001 GND!    Xa2s_dout[6]/27:2 1.624E-16
C442002 Xopctrl.A2Sop/Lc[2][10].0:8     Vdd! 2.448E-16
.ENDS
