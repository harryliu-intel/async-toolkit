///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_fwd_misc_map.sv                                    
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_fwd_misc_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_FF
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_FF

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_RSTD


module rtlgen_mby_ppe_fwd_misc_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_fwd_misc_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_PH2_FF
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_FWD_MISC_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_fwd_misc_map ( //lintra s-2096
    // Clocks
    gated_clk,
    rtl_clk,

    // Resets
    rst_n,


    // Register Inputs
    load_FWD_IP,

    new_FWD_IM,
    new_FWD_IP,

    handcode_reg_rdata_FWD_LAG_CFG,
    handcode_reg_rdata_FWD_PORT_CFG_1,
    handcode_reg_rdata_FWD_PORT_CFG_2,

    handcode_rvalid_FWD_LAG_CFG,
    handcode_rvalid_FWD_PORT_CFG_1,
    handcode_rvalid_FWD_PORT_CFG_2,

    handcode_wvalid_FWD_LAG_CFG,
    handcode_wvalid_FWD_PORT_CFG_1,
    handcode_wvalid_FWD_PORT_CFG_2,

    handcode_error_FWD_LAG_CFG,
    handcode_error_FWD_PORT_CFG_1,
    handcode_error_FWD_PORT_CFG_2,


    // Register Outputs
    FWD_CPU_MAC,
    FWD_IEEE_RESERVED_MAC_ACTION,
    FWD_IEEE_RESERVED_MAC_CFG,
    FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY,
    FWD_IM,
    FWD_IP,
    FWD_QCN_MIRROR_CFG,
    FWD_RX_MIRROR_CFG,
    FWD_SYS_CFG_1,
    FWD_SYS_CFG_ROUTER,


    // Register signals for HandCoded registers
    handcode_reg_wdata_FWD_LAG_CFG,
    handcode_reg_wdata_FWD_PORT_CFG_1,
    handcode_reg_wdata_FWD_PORT_CFG_2,

    we_FWD_LAG_CFG,
    we_FWD_PORT_CFG_1,
    we_FWD_PORT_CFG_2,

    re_FWD_LAG_CFG,
    re_FWD_PORT_CFG_1,
    re_FWD_PORT_CFG_2,




    // Config Access
    req,
    ack
    

);

import mby_ppe_fwd_misc_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:0] MBY_PPE_FWD_MISC_MAP_OFFSET = {MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] FWD_MISC_SB_BAR = 3'b0;
parameter [7:0] FWD_MISC_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_SYS_CFG_1_DECODE_ADDR = FWD_SYS_CFG_1_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_CPU_MAC_DECODE_ADDR = FWD_CPU_MAC_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_SYS_CFG_ROUTER_DECODE_ADDR = FWD_SYS_CFG_ROUTER_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_RX_MIRROR_CFG_DECODE_ADDR = FWD_RX_MIRROR_CFG_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_QCN_MIRROR_CFG_DECODE_ADDR = FWD_QCN_MIRROR_CFG_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_IEEE_RESERVED_MAC_ACTION_DECODE_ADDR = FWD_IEEE_RESERVED_MAC_ACTION_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_DECODE_ADDR = FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_IEEE_RESERVED_MAC_CFG_DECODE_ADDR = FWD_IEEE_RESERVED_MAC_CFG_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_IP_DECODE_ADDR = FWD_IP_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] FWD_IM_DECODE_ADDR = FWD_IM_CR_ADDR[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_FWD_MISC_MAP_OFFSET[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];

    // Clocks
input logic  gated_clk;
input logic  rtl_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input load_FWD_IP_t  load_FWD_IP;

input new_FWD_IM_t  new_FWD_IM;
input new_FWD_IP_t  new_FWD_IP;

input FWD_LAG_CFG_t  handcode_reg_rdata_FWD_LAG_CFG;
input FWD_PORT_CFG_1_t  handcode_reg_rdata_FWD_PORT_CFG_1;
input FWD_PORT_CFG_2_t  handcode_reg_rdata_FWD_PORT_CFG_2;

input handcode_rvalid_FWD_LAG_CFG_t  handcode_rvalid_FWD_LAG_CFG;
input handcode_rvalid_FWD_PORT_CFG_1_t  handcode_rvalid_FWD_PORT_CFG_1;
input handcode_rvalid_FWD_PORT_CFG_2_t  handcode_rvalid_FWD_PORT_CFG_2;

input handcode_wvalid_FWD_LAG_CFG_t  handcode_wvalid_FWD_LAG_CFG;
input handcode_wvalid_FWD_PORT_CFG_1_t  handcode_wvalid_FWD_PORT_CFG_1;
input handcode_wvalid_FWD_PORT_CFG_2_t  handcode_wvalid_FWD_PORT_CFG_2;

input handcode_error_FWD_LAG_CFG_t  handcode_error_FWD_LAG_CFG;
input handcode_error_FWD_PORT_CFG_1_t  handcode_error_FWD_PORT_CFG_1;
input handcode_error_FWD_PORT_CFG_2_t  handcode_error_FWD_PORT_CFG_2;


    // Register Outputs
output FWD_CPU_MAC_t  FWD_CPU_MAC;
output FWD_IEEE_RESERVED_MAC_ACTION_t  FWD_IEEE_RESERVED_MAC_ACTION;
output FWD_IEEE_RESERVED_MAC_CFG_t  FWD_IEEE_RESERVED_MAC_CFG;
output FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_t  FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY;
output FWD_IM_t  FWD_IM;
output FWD_IP_t  FWD_IP;
output FWD_QCN_MIRROR_CFG_t  FWD_QCN_MIRROR_CFG;
output FWD_RX_MIRROR_CFG_t  FWD_RX_MIRROR_CFG;
output FWD_SYS_CFG_1_t  FWD_SYS_CFG_1;
output FWD_SYS_CFG_ROUTER_t  FWD_SYS_CFG_ROUTER;


    // Register signals for HandCoded registers
output FWD_LAG_CFG_t  handcode_reg_wdata_FWD_LAG_CFG;
output FWD_PORT_CFG_1_t  handcode_reg_wdata_FWD_PORT_CFG_1;
output FWD_PORT_CFG_2_t  handcode_reg_wdata_FWD_PORT_CFG_2;

output we_FWD_LAG_CFG_t  we_FWD_LAG_CFG;
output we_FWD_PORT_CFG_1_t  we_FWD_PORT_CFG_1;
output we_FWD_PORT_CFG_2_t  we_FWD_PORT_CFG_2;

output re_FWD_LAG_CFG_t  re_FWD_LAG_CFG;
output re_FWD_PORT_CFG_1_t  re_FWD_PORT_CFG_1;
output re_FWD_PORT_CFG_2_t  re_FWD_PORT_CFG_2;




    // Config Access
input mby_ppe_fwd_misc_map_cr_req_t  req;
output mby_ppe_fwd_misc_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_fwd_misc_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_FWD_MISC_MAP_MEM;
assign case_req_addr_MBY_PPE_FWD_MISC_MAP_MEM = req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_fwd_misc;
always_comb begin : sb_fid_cond_fwd_misc_BLOCK
    unique casez (req_fid) 
		FWD_MISC_SB_FID: sb_fid_cond_fwd_misc = 1;
		default: sb_fid_cond_fwd_misc = 0;
    endcase 
end


logic sb_bar_cond_fwd_misc;
always_comb begin : sb_bar_cond_fwd_misc_BLOCK
    unique casez (req_bar) 
		FWD_MISC_SB_BAR: sb_bar_cond_fwd_misc = 1;
		default: sb_bar_cond_fwd_misc = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// FWD_PORT_CFG_2 using HANDCODED_REG template.
logic addr_decode_FWD_PORT_CFG_2;
logic write_req_FWD_PORT_CFG_2;
logic read_req_FWD_PORT_CFG_2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b0???,4'h?,1'b?}: 
         addr_decode_FWD_PORT_CFG_2 = req.valid;
      default: 
         addr_decode_FWD_PORT_CFG_2 = 1'b0; 
   endcase
end

always_comb write_req_FWD_PORT_CFG_2 = f_IsMEMWr(req_opcode) && addr_decode_FWD_PORT_CFG_2 ;
always_comb read_req_FWD_PORT_CFG_2  = f_IsMEMRd(req_opcode) && addr_decode_FWD_PORT_CFG_2 ;

always_comb we_FWD_PORT_CFG_2 = {8{write_req_FWD_PORT_CFG_2}} & be;
always_comb re_FWD_PORT_CFG_2 = {8{read_req_FWD_PORT_CFG_2}} & be;
always_comb handcode_reg_wdata_FWD_PORT_CFG_2 = write_data;


// ----------------------------------------------------------------------
// FWD_LAG_CFG using HANDCODED_REG template.
logic addr_decode_FWD_LAG_CFG;
logic write_req_FWD_LAG_CFG;
logic read_req_FWD_LAG_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h10,4'b0???,1'b?},
      {44'h108,1'b0}:
          addr_decode_FWD_LAG_CFG = req.valid;
      default: 
         addr_decode_FWD_LAG_CFG = 1'b0; 
   endcase
end

always_comb write_req_FWD_LAG_CFG = f_IsMEMWr(req_opcode) && addr_decode_FWD_LAG_CFG ;
always_comb read_req_FWD_LAG_CFG  = f_IsMEMRd(req_opcode) && addr_decode_FWD_LAG_CFG ;

always_comb we_FWD_LAG_CFG = {8{write_req_FWD_LAG_CFG}} & be;
always_comb re_FWD_LAG_CFG = {8{read_req_FWD_LAG_CFG}} & be;
always_comb handcode_reg_wdata_FWD_LAG_CFG = write_data;


// ----------------------------------------------------------------------
// FWD_PORT_CFG_1 using HANDCODED_REG template.
logic addr_decode_FWD_PORT_CFG_1;
logic write_req_FWD_PORT_CFG_1;
logic read_req_FWD_PORT_CFG_1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h11,4'b0???,1'b?},
      {44'h118,1'b0}:
          addr_decode_FWD_PORT_CFG_1 = req.valid;
      default: 
         addr_decode_FWD_PORT_CFG_1 = 1'b0; 
   endcase
end

always_comb write_req_FWD_PORT_CFG_1 = f_IsMEMWr(req_opcode) && addr_decode_FWD_PORT_CFG_1 ;
always_comb read_req_FWD_PORT_CFG_1  = f_IsMEMRd(req_opcode) && addr_decode_FWD_PORT_CFG_1 ;

always_comb we_FWD_PORT_CFG_1 = {8{write_req_FWD_PORT_CFG_1}} & be;
always_comb re_FWD_PORT_CFG_1 = {8{read_req_FWD_PORT_CFG_1}} & be;
always_comb handcode_reg_wdata_FWD_PORT_CFG_1 = write_data;


//---------------------------------------------------------------------
// FWD_SYS_CFG_1 Address Decode
logic  addr_decode_FWD_SYS_CFG_1;
logic  write_req_FWD_SYS_CFG_1;
always_comb begin
   addr_decode_FWD_SYS_CFG_1 = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_SYS_CFG_1_DECODE_ADDR) && req.valid ;
   write_req_FWD_SYS_CFG_1 = IsMEMWr && addr_decode_FWD_SYS_CFG_1 && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_SYS_CFG_1.TRAP_MTU_VIOLATIONS x1 RW, using RW template.
logic [0:0] up_FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS;
always_comb begin
 up_FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS =
    ({1{write_req_FWD_SYS_CFG_1 }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS;
always_comb begin
 nxt_FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS = write_data[0:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS[0], nxt_FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS[0:0], FWD_SYS_CFG_1.TRAP_MTU_VIOLATIONS[0:0])

// ----------------------------------------------------------------------
// FWD_SYS_CFG_1.ENABLE_TRAP_PLUS_LOG x1 RW, using RW template.
logic [0:0] up_FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG;
always_comb begin
 up_FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG =
    ({1{write_req_FWD_SYS_CFG_1 }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG;
always_comb begin
 nxt_FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG = write_data[1:1];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG[0], nxt_FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG[0:0], FWD_SYS_CFG_1.ENABLE_TRAP_PLUS_LOG[0:0])

// ----------------------------------------------------------------------
// FWD_SYS_CFG_1.DROP_INVALID_SMAC x1 RW, using RW template.
logic [0:0] up_FWD_SYS_CFG_1_DROP_INVALID_SMAC;
always_comb begin
 up_FWD_SYS_CFG_1_DROP_INVALID_SMAC =
    ({1{write_req_FWD_SYS_CFG_1 }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_SYS_CFG_1_DROP_INVALID_SMAC;
always_comb begin
 nxt_FWD_SYS_CFG_1_DROP_INVALID_SMAC = write_data[2:2];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_SYS_CFG_1_DROP_INVALID_SMAC[0], nxt_FWD_SYS_CFG_1_DROP_INVALID_SMAC[0:0], FWD_SYS_CFG_1.DROP_INVALID_SMAC[0:0])

// ----------------------------------------------------------------------
// FWD_SYS_CFG_1.DROP_MAC_CTRL_ETHERTYPE x1 RW, using RW template.
logic [0:0] up_FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE;
always_comb begin
 up_FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE =
    ({1{write_req_FWD_SYS_CFG_1 }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE;
always_comb begin
 nxt_FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE = write_data[3:3];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE[0], nxt_FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE[0:0], FWD_SYS_CFG_1.DROP_MAC_CTRL_ETHERTYPE[0:0])

// ----------------------------------------------------------------------
// FWD_SYS_CFG_1.STORE_TRAP_ACTION x1 RW, using RW template.
logic [0:0] up_FWD_SYS_CFG_1_STORE_TRAP_ACTION;
always_comb begin
 up_FWD_SYS_CFG_1_STORE_TRAP_ACTION =
    ({1{write_req_FWD_SYS_CFG_1 }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_SYS_CFG_1_STORE_TRAP_ACTION;
always_comb begin
 nxt_FWD_SYS_CFG_1_STORE_TRAP_ACTION = write_data[4:4];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_SYS_CFG_1_STORE_TRAP_ACTION[0], nxt_FWD_SYS_CFG_1_STORE_TRAP_ACTION[0:0], FWD_SYS_CFG_1.STORE_TRAP_ACTION[0:0])

//---------------------------------------------------------------------
// FWD_CPU_MAC Address Decode
logic  addr_decode_FWD_CPU_MAC;
logic  write_req_FWD_CPU_MAC;
always_comb begin
   addr_decode_FWD_CPU_MAC = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_CPU_MAC_DECODE_ADDR) && req.valid ;
   write_req_FWD_CPU_MAC = IsMEMWr && addr_decode_FWD_CPU_MAC && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_CPU_MAC.MAC_ADDR x8 RW, using RW template.
logic [5:0] up_FWD_CPU_MAC_MAC_ADDR;
always_comb begin
 up_FWD_CPU_MAC_MAC_ADDR =
    ({6{write_req_FWD_CPU_MAC }} &
    be[5:0]);
end

logic [47:0] nxt_FWD_CPU_MAC_MAC_ADDR;
always_comb begin
 nxt_FWD_CPU_MAC_MAC_ADDR = write_data[47:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_CPU_MAC_MAC_ADDR[0], nxt_FWD_CPU_MAC_MAC_ADDR[7:0], FWD_CPU_MAC.MAC_ADDR[7:0])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_CPU_MAC_MAC_ADDR[1], nxt_FWD_CPU_MAC_MAC_ADDR[15:8], FWD_CPU_MAC.MAC_ADDR[15:8])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_CPU_MAC_MAC_ADDR[2], nxt_FWD_CPU_MAC_MAC_ADDR[23:16], FWD_CPU_MAC.MAC_ADDR[23:16])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_CPU_MAC_MAC_ADDR[3], nxt_FWD_CPU_MAC_MAC_ADDR[31:24], FWD_CPU_MAC.MAC_ADDR[31:24])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_CPU_MAC_MAC_ADDR[4], nxt_FWD_CPU_MAC_MAC_ADDR[39:32], FWD_CPU_MAC.MAC_ADDR[39:32])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_CPU_MAC_MAC_ADDR[5], nxt_FWD_CPU_MAC_MAC_ADDR[47:40], FWD_CPU_MAC.MAC_ADDR[47:40])

//---------------------------------------------------------------------
// FWD_SYS_CFG_ROUTER Address Decode
logic  addr_decode_FWD_SYS_CFG_ROUTER;
logic  write_req_FWD_SYS_CFG_ROUTER;
always_comb begin
   addr_decode_FWD_SYS_CFG_ROUTER = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_SYS_CFG_ROUTER_DECODE_ADDR) && req.valid ;
   write_req_FWD_SYS_CFG_ROUTER = IsMEMWr && addr_decode_FWD_SYS_CFG_ROUTER && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_SYS_CFG_ROUTER.TRAP_TTL1 x2 RW, using RW template.
logic [0:0] up_FWD_SYS_CFG_ROUTER_TRAP_TTL1;
always_comb begin
 up_FWD_SYS_CFG_ROUTER_TRAP_TTL1 =
    ({1{write_req_FWD_SYS_CFG_ROUTER }} &
    be[0:0]);
end

logic [1:0] nxt_FWD_SYS_CFG_ROUTER_TRAP_TTL1;
always_comb begin
 nxt_FWD_SYS_CFG_ROUTER_TRAP_TTL1 = write_data[1:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_FWD_SYS_CFG_ROUTER_TRAP_TTL1[0], nxt_FWD_SYS_CFG_ROUTER_TRAP_TTL1[1:0], FWD_SYS_CFG_ROUTER.TRAP_TTL1[1:0])

// ----------------------------------------------------------------------
// FWD_SYS_CFG_ROUTER.TRAP_IP_OPTIONS x1 RW, using RW template.
logic [0:0] up_FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS;
always_comb begin
 up_FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS =
    ({1{write_req_FWD_SYS_CFG_ROUTER }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS;
always_comb begin
 nxt_FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS = write_data[2:2];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS[0], nxt_FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS[0:0], FWD_SYS_CFG_ROUTER.TRAP_IP_OPTIONS[0:0])

//---------------------------------------------------------------------
// FWD_RX_MIRROR_CFG Address Decode
logic  addr_decode_FWD_RX_MIRROR_CFG;
logic  write_req_FWD_RX_MIRROR_CFG;
always_comb begin
   addr_decode_FWD_RX_MIRROR_CFG = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_RX_MIRROR_CFG_DECODE_ADDR) && req.valid ;
   write_req_FWD_RX_MIRROR_CFG = IsMEMWr && addr_decode_FWD_RX_MIRROR_CFG && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_RX_MIRROR_CFG.MIRROR_PROFILE_IDX x6 RW, using RW template.
logic [0:0] up_FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX;
always_comb begin
 up_FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX =
    ({1{write_req_FWD_RX_MIRROR_CFG }} &
    be[0:0]);
end

logic [5:0] nxt_FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX;
always_comb begin
 nxt_FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX = write_data[5:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 6'h0, up_FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX[0], nxt_FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX[5:0], FWD_RX_MIRROR_CFG.MIRROR_PROFILE_IDX[5:0])

//---------------------------------------------------------------------
// FWD_QCN_MIRROR_CFG Address Decode
logic  addr_decode_FWD_QCN_MIRROR_CFG;
logic  write_req_FWD_QCN_MIRROR_CFG;
always_comb begin
   addr_decode_FWD_QCN_MIRROR_CFG = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_QCN_MIRROR_CFG_DECODE_ADDR) && req.valid ;
   write_req_FWD_QCN_MIRROR_CFG = IsMEMWr && addr_decode_FWD_QCN_MIRROR_CFG && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_QCN_MIRROR_CFG.MIRROR_SESSION x2 RW, using RW template.
logic [0:0] up_FWD_QCN_MIRROR_CFG_MIRROR_SESSION;
always_comb begin
 up_FWD_QCN_MIRROR_CFG_MIRROR_SESSION =
    ({1{write_req_FWD_QCN_MIRROR_CFG }} &
    be[0:0]);
end

logic [1:0] nxt_FWD_QCN_MIRROR_CFG_MIRROR_SESSION;
always_comb begin
 nxt_FWD_QCN_MIRROR_CFG_MIRROR_SESSION = write_data[1:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_FWD_QCN_MIRROR_CFG_MIRROR_SESSION[0], nxt_FWD_QCN_MIRROR_CFG_MIRROR_SESSION[1:0], FWD_QCN_MIRROR_CFG.MIRROR_SESSION[1:0])

// ----------------------------------------------------------------------
// FWD_QCN_MIRROR_CFG.MIRROR_PROFILE_IDX x6 RW, using RW template.
logic [0:0] up_FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX;
always_comb begin
 up_FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX =
    ({1{write_req_FWD_QCN_MIRROR_CFG }} &
    be[0:0]);
end

logic [5:0] nxt_FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX;
always_comb begin
 nxt_FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX = write_data[7:2];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 6'h0, up_FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX[0], nxt_FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX[5:0], FWD_QCN_MIRROR_CFG.MIRROR_PROFILE_IDX[5:0])

//---------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION Address Decode
logic  addr_decode_FWD_IEEE_RESERVED_MAC_ACTION;
logic  write_req_FWD_IEEE_RESERVED_MAC_ACTION;
always_comb begin
   addr_decode_FWD_IEEE_RESERVED_MAC_ACTION = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_IEEE_RESERVED_MAC_ACTION_DECODE_ADDR) && req.valid ;
   write_req_FWD_IEEE_RESERVED_MAC_ACTION = IsMEMWr && addr_decode_FWD_IEEE_RESERVED_MAC_ACTION && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_0 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[0:0]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0 = write_data[1:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_0[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_1 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[0:0]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1 = write_data[3:2];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_1[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_2 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[0:0]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2 = write_data[5:4];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_2[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_3 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[0:0]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3 = write_data[7:6];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_3[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_4 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[1:1]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4 = write_data[9:8];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_4[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_5 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[1:1]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5 = write_data[11:10];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_5[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_6 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[1:1]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6 = write_data[13:12];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_6[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_7 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[1:1]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7 = write_data[15:14];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_7[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_8 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[2:2]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8 = write_data[17:16];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_8[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_9 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[2:2]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9 = write_data[19:18];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_9[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_10 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[2:2]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10 = write_data[21:20];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_10[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_11 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[2:2]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11 = write_data[23:22];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_11[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_12 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[3:3]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12 = write_data[25:24];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_12[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_13 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[3:3]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13 = write_data[27:26];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_13[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_14 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[3:3]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14 = write_data[29:28];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_14[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_15 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[3:3]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15 = write_data[31:30];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_15[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_16 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[4:4]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16 = write_data[33:32];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_16[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_17 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[4:4]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17 = write_data[35:34];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_17[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_18 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[4:4]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18 = write_data[37:36];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_18[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_19 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[4:4]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19 = write_data[39:38];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_19[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_20 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[5:5]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20 = write_data[41:40];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_20[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_21 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[5:5]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21 = write_data[43:42];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_21[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_22 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[5:5]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22 = write_data[45:44];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_22[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_23 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[5:5]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23 = write_data[47:46];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_23[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_24 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[6:6]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24 = write_data[49:48];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_24[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_25 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[6:6]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25 = write_data[51:50];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_25[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_26 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[6:6]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26 = write_data[53:52];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_26[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_27 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[6:6]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27 = write_data[55:54];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_27[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_28 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[7:7]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28 = write_data[57:56];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_28[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_29 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[7:7]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29 = write_data[59:58];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_29[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_30 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[7:7]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30 = write_data[61:60];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_30[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_31 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[7:7]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31 = write_data[63:62];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_31[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_32 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[8:8]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32 = write_data[65:64];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_32[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_33 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[8:8]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33 = write_data[67:66];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_33[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_34 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[8:8]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34 = write_data[69:68];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_34[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_35 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[8:8]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35 = write_data[71:70];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_35[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_36 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[9:9]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36 = write_data[73:72];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_36[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_37 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[9:9]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37 = write_data[75:74];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_37[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_38 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[9:9]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38 = write_data[77:76];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_38[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_39 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[9:9]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39 = write_data[79:78];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_39[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_40 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[10:10]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40 = write_data[81:80];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_40[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_41 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[10:10]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41 = write_data[83:82];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_41[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_42 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[10:10]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42 = write_data[85:84];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_42[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_43 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[10:10]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43 = write_data[87:86];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_43[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_44 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[11:11]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44 = write_data[89:88];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_44[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_45 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[11:11]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45 = write_data[91:90];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_45[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_46 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[11:11]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46 = write_data[93:92];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_46[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_47 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[11:11]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47 = write_data[95:94];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_47[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_48 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[12:12]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48 = write_data[97:96];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_48[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_49 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[12:12]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49 = write_data[99:98];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_49[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_50 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[12:12]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50 = write_data[101:100];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_50[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_51 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[12:12]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51 = write_data[103:102];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_51[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_52 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[13:13]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52 = write_data[105:104];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_52[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_53 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[13:13]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53 = write_data[107:106];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_53[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_54 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[13:13]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54 = write_data[109:108];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_54[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_55 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[13:13]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55 = write_data[111:110];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_55[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_56 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[14:14]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56 = write_data[113:112];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_56[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_57 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[14:14]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57 = write_data[115:114];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_57[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_58 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[14:14]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58 = write_data[117:116];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_58[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_59 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[14:14]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59 = write_data[119:118];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_59[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_60 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[15:15]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60 = write_data[121:120];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_60[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_61 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[15:15]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61 = write_data[123:122];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_61[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_62 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[15:15]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62 = write_data[125:124];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_62[1:0])

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_ACTION.ACTION_63 x2 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63 =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_ACTION }} &
    be[15:15]);
end

logic [1:0] nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63 = write_data[127:126];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 2'h2, up_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63[0], nxt_FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63[1:0], FWD_IEEE_RESERVED_MAC_ACTION.ACTION_63[1:0])

//---------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY Address Decode
logic  addr_decode_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY;
logic  write_req_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY;
always_comb begin
   addr_decode_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_DECODE_ADDR) && req.valid ;
   write_req_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY = IsMEMWr && addr_decode_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT x8 RW, using RW template.
logic [7:0] up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT =
    ({8{write_req_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY }} &
    be[7:0]);
end

logic [63:0] nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT = write_data[63:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[0], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[7:0], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[7:0])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[1], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[15:8], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[15:8])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[2], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[23:16], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[23:16])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[3], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[31:24], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[31:24])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[4], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[39:32], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[39:32])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[5], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[47:40], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[47:40])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[6], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[55:48], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[55:48])
`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[7], nxt_FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT[63:56], FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY.SELECT[63:56])

//---------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_CFG Address Decode
logic  addr_decode_FWD_IEEE_RESERVED_MAC_CFG;
logic  write_req_FWD_IEEE_RESERVED_MAC_CFG;
always_comb begin
   addr_decode_FWD_IEEE_RESERVED_MAC_CFG = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_IEEE_RESERVED_MAC_CFG_DECODE_ADDR) && req.valid ;
   write_req_FWD_IEEE_RESERVED_MAC_CFG = IsMEMWr && addr_decode_FWD_IEEE_RESERVED_MAC_CFG && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_IEEE_RESERVED_MAC_CFG.TRAP_TC x3 RW, using RW template.
logic [0:0] up_FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC;
always_comb begin
 up_FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC =
    ({1{write_req_FWD_IEEE_RESERVED_MAC_CFG }} &
    be[0:0]);
end

logic [2:0] nxt_FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC;
always_comb begin
 nxt_FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC = write_data[2:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 3'h0, up_FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC[0], nxt_FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC[2:0], FWD_IEEE_RESERVED_MAC_CFG.TRAP_TC[2:0])

//---------------------------------------------------------------------
// FWD_IP Address Decode
logic  addr_decode_FWD_IP;
logic  write_req_FWD_IP;
always_comb begin
   addr_decode_FWD_IP = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_IP_DECODE_ADDR) && req.valid ;
   write_req_FWD_IP = IsMEMWr && addr_decode_FWD_IP && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_IP.SHELL_CTRL_U_ERR x1 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [0:0] req_up_FWD_IP_SHELL_CTRL_U_ERR;
always_comb begin
 req_up_FWD_IP_SHELL_CTRL_U_ERR[0:0] = 
   {1{write_req_FWD_IP & be[0]}}
;
end

logic [0:0] clr_FWD_IP_SHELL_CTRL_U_ERR;
always_comb begin
 clr_FWD_IP_SHELL_CTRL_U_ERR = write_data[0:0] & req_up_FWD_IP_SHELL_CTRL_U_ERR;

end
logic [0:0] swwr_FWD_IP_SHELL_CTRL_U_ERR;
logic [0:0] sw_nxt_FWD_IP_SHELL_CTRL_U_ERR;
always_comb begin
 swwr_FWD_IP_SHELL_CTRL_U_ERR = clr_FWD_IP_SHELL_CTRL_U_ERR;
 sw_nxt_FWD_IP_SHELL_CTRL_U_ERR = {1{1'b0}};

end
logic [0:0] up_FWD_IP_SHELL_CTRL_U_ERR;
logic [0:0] nxt_FWD_IP_SHELL_CTRL_U_ERR;
always_comb begin
 up_FWD_IP_SHELL_CTRL_U_ERR = 
   swwr_FWD_IP_SHELL_CTRL_U_ERR | {1{load_FWD_IP.SHELL_CTRL_U_ERR}};
end
always_comb begin
 nxt_FWD_IP_SHELL_CTRL_U_ERR[0] = 
    load_FWD_IP.SHELL_CTRL_U_ERR ?
    new_FWD_IP.SHELL_CTRL_U_ERR[0] :
    sw_nxt_FWD_IP_SHELL_CTRL_U_ERR[0];
end



`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_FWD_IP_SHELL_CTRL_U_ERR[0], nxt_FWD_IP_SHELL_CTRL_U_ERR[0], FWD_IP.SHELL_CTRL_U_ERR[0])
// ----------------------------------------------------------------------
// FWD_IP.ENTRY_COUNT x1 RO/V, using RO/V template.
assign FWD_IP.ENTRY_COUNT = new_FWD_IP.ENTRY_COUNT;



// ----------------------------------------------------------------------
// FWD_IP.TCAM_ERR x1 RO/V, using RO/V template.
assign FWD_IP.TCAM_ERR = new_FWD_IP.TCAM_ERR;



// ----------------------------------------------------------------------
// FWD_IP.TRIGGER x1 RO/V, using RO/V template.
assign FWD_IP.TRIGGER = new_FWD_IP.TRIGGER;




// ----------------------------------------------------------------------
// FWD_IP.WB_FIFO_PERR x1 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [0:0] req_up_FWD_IP_WB_FIFO_PERR;
always_comb begin
 req_up_FWD_IP_WB_FIFO_PERR[0:0] = 
   {1{write_req_FWD_IP & be[0]}}
;
end

logic [0:0] clr_FWD_IP_WB_FIFO_PERR;
always_comb begin
 clr_FWD_IP_WB_FIFO_PERR = write_data[4:4] & req_up_FWD_IP_WB_FIFO_PERR;

end
logic [0:0] swwr_FWD_IP_WB_FIFO_PERR;
logic [0:0] sw_nxt_FWD_IP_WB_FIFO_PERR;
always_comb begin
 swwr_FWD_IP_WB_FIFO_PERR = clr_FWD_IP_WB_FIFO_PERR;
 sw_nxt_FWD_IP_WB_FIFO_PERR = {1{1'b0}};

end
logic [0:0] up_FWD_IP_WB_FIFO_PERR;
logic [0:0] nxt_FWD_IP_WB_FIFO_PERR;
always_comb begin
 up_FWD_IP_WB_FIFO_PERR = 
   swwr_FWD_IP_WB_FIFO_PERR | {1{load_FWD_IP.WB_FIFO_PERR}};
end
always_comb begin
 nxt_FWD_IP_WB_FIFO_PERR[0] = 
    load_FWD_IP.WB_FIFO_PERR ?
    new_FWD_IP.WB_FIFO_PERR[0] :
    sw_nxt_FWD_IP_WB_FIFO_PERR[0];
end



`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_FWD_IP_WB_FIFO_PERR[0], nxt_FWD_IP_WB_FIFO_PERR[0], FWD_IP.WB_FIFO_PERR[0])
// ----------------------------------------------------------------------
// FWD_IP.MA_TCN x1 RO/V, using RO/V template.
assign FWD_IP.MA_TCN = new_FWD_IP.MA_TCN;




//---------------------------------------------------------------------
// FWD_IM Address Decode
logic  addr_decode_FWD_IM;
logic  write_req_FWD_IM;
always_comb begin
   addr_decode_FWD_IM = (req_addr[MBY_PPE_FWD_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == FWD_IM_DECODE_ADDR) && req.valid ;
   write_req_FWD_IM = IsMEMWr && addr_decode_FWD_IM && sb_fid_cond_fwd_misc && sb_bar_cond_fwd_misc;
end

// ----------------------------------------------------------------------
// FWD_IM.SHELL_CTRL_U_ERR x1 RW, using RW template.
logic [0:0] up_FWD_IM_SHELL_CTRL_U_ERR;
always_comb begin
 up_FWD_IM_SHELL_CTRL_U_ERR =
    ({1{write_req_FWD_IM }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_IM_SHELL_CTRL_U_ERR;
always_comb begin
 nxt_FWD_IM_SHELL_CTRL_U_ERR = write_data[0:0];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_IM_SHELL_CTRL_U_ERR[0], nxt_FWD_IM_SHELL_CTRL_U_ERR[0:0], FWD_IM.SHELL_CTRL_U_ERR[0:0])

// ----------------------------------------------------------------------
// FWD_IM.ENTRY_COUNT x1 RW, using RW template.
logic [0:0] up_FWD_IM_ENTRY_COUNT;
always_comb begin
 up_FWD_IM_ENTRY_COUNT =
    ({1{write_req_FWD_IM }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_IM_ENTRY_COUNT;
always_comb begin
 nxt_FWD_IM_ENTRY_COUNT = write_data[1:1];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_IM_ENTRY_COUNT[0], nxt_FWD_IM_ENTRY_COUNT[0:0], FWD_IM.ENTRY_COUNT[0:0])

// ----------------------------------------------------------------------
// FWD_IM.TCAM_ERR x1 RW, using RW template.
logic [0:0] up_FWD_IM_TCAM_ERR;
always_comb begin
 up_FWD_IM_TCAM_ERR =
    ({1{write_req_FWD_IM }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_IM_TCAM_ERR;
always_comb begin
 nxt_FWD_IM_TCAM_ERR = write_data[2:2];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_IM_TCAM_ERR[0], nxt_FWD_IM_TCAM_ERR[0:0], FWD_IM.TCAM_ERR[0:0])

// ----------------------------------------------------------------------
// FWD_IM.TRIGGER x1 RW, using RW template.
logic [0:0] up_FWD_IM_TRIGGER;
always_comb begin
 up_FWD_IM_TRIGGER =
    ({1{write_req_FWD_IM }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_IM_TRIGGER;
always_comb begin
 nxt_FWD_IM_TRIGGER = write_data[3:3];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_IM_TRIGGER[0], nxt_FWD_IM_TRIGGER[0:0], FWD_IM.TRIGGER[0:0])

// ----------------------------------------------------------------------
// FWD_IM.WB_FIFO_PERR x1 RW, using RW template.
logic [0:0] up_FWD_IM_WB_FIFO_PERR;
always_comb begin
 up_FWD_IM_WB_FIFO_PERR =
    ({1{write_req_FWD_IM }} &
    be[0:0]);
end

logic [0:0] nxt_FWD_IM_WB_FIFO_PERR;
always_comb begin
 nxt_FWD_IM_WB_FIFO_PERR = write_data[4:4];

end


`RTLGEN_MBY_PPE_FWD_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_FWD_IM_WB_FIFO_PERR[0], nxt_FWD_IM_WB_FIFO_PERR[0:0], FWD_IM.WB_FIFO_PERR[0:0])
// ----------------------------------------------------------------------
// FWD_IM.MA_TCN x1 RO/V, using RO/V template.
assign FWD_IM.MA_TCN = new_FWD_IM.MA_TCN;




// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_FWD_MISC_MAP_MEM) 
           {40'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_FWD_PORT_CFG_2;
                    ack.read_miss = handcode_error_FWD_PORT_CFG_2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h10,4'b0???,1'b?},
           {44'h108,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_FWD_LAG_CFG;
                    ack.read_miss = handcode_error_FWD_LAG_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h11,4'b0???,1'b?},
           {44'h118,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_FWD_PORT_CFG_1;
                    ack.read_miss = handcode_error_FWD_PORT_CFG_1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_SYS_CFG_1_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_CPU_MAC_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_SYS_CFG_ROUTER_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_RX_MIRROR_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_QCN_MIRROR_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_ACTION_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           FWD_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_FWD_MISC_MAP_MEM) 
           {40'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_FWD_PORT_CFG_2;
                    ack.write_miss = handcode_error_FWD_PORT_CFG_2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h10,4'b0???,1'b?},
           {44'h108,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_FWD_LAG_CFG;
                    ack.write_miss = handcode_error_FWD_LAG_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h11,4'b0???,1'b?},
           {44'h118,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_FWD_PORT_CFG_1;
                    ack.write_miss = handcode_error_FWD_PORT_CFG_1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_SYS_CFG_1_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_CPU_MAC_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_SYS_CFG_ROUTER_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_RX_MIRROR_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_QCN_MIRROR_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_ACTION_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           FWD_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_FWD_MISC_MAP_MEM) 
           {40'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = handcode_reg_rdata_FWD_PORT_CFG_2;
                 default: read_data = '0;
              endcase
           end
           {40'h10,4'b0???,1'b?},
           {44'h108,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = handcode_reg_rdata_FWD_LAG_CFG;
                 default: read_data = '0;
              endcase
           end
           {40'h11,4'b0???,1'b?},
           {44'h118,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = handcode_reg_rdata_FWD_PORT_CFG_1;
                 default: read_data = '0;
              endcase
           end
           FWD_SYS_CFG_1_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_SYS_CFG_1};
                 default: read_data = '0;
              endcase
           end
           FWD_CPU_MAC_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_CPU_MAC};
                 default: read_data = '0;
              endcase
           end
           FWD_SYS_CFG_ROUTER_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_SYS_CFG_ROUTER};
                 default: read_data = '0;
              endcase
           end
           FWD_RX_MIRROR_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_RX_MIRROR_CFG};
                 default: read_data = '0;
              endcase
           end
           FWD_QCN_MIRROR_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_QCN_MIRROR_CFG};
                 default: read_data = '0;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_ACTION_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_IEEE_RESERVED_MAC_ACTION};
                 default: read_data = '0;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY};
                 default: read_data = '0;
              endcase
           end
           FWD_IEEE_RESERVED_MAC_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_IEEE_RESERVED_MAC_CFG};
                 default: read_data = '0;
              endcase
           end
           FWD_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_IP};
                 default: read_data = '0;
              endcase
           end
           FWD_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {FWD_MISC_SB_FID,FWD_MISC_SB_BAR}: read_data = {FWD_IM};
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    FWD_SYS_CFG_1.reserved0 = '0;
    FWD_CPU_MAC.reserved0 = '0;
    FWD_SYS_CFG_ROUTER.reserved0 = '0;
    FWD_RX_MIRROR_CFG.reserved0 = '0;
    FWD_QCN_MIRROR_CFG.reserved0 = '0;
    FWD_IEEE_RESERVED_MAC_CFG.reserved0 = '0;
    FWD_IP.reserved0 = '0;
    FWD_IM.reserved0 = '0;
end

// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
