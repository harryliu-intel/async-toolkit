
/* ----------------------------------------------------------------------


   ----------------------------------------------------------------------
   file:    mby_fuse_env.sv
   Date Created  :mby_Fuse_Map_env.svh 25/7/2016
   Author        : dbenita
   Project       : MBY IP
   ----------------------------------------------------------------------
 
  MBY Soala FUSE ENV

  This file include the MBY IP configuration for fuses
 
 In this file the IP can add constraints on fuse and addd IP
 specific code for the IP fuses
 
 

*/

//Include mby regs
import ovm_pkg::*;
import sla_pkg::*;
`include "ovm_macros.svh"
`include "sla_macros.svh"
  
class mby_fuse_env extends toplevel_fuse_env;
   `ovm_component_utils(mby_fuse_env);

`include "fusegen_api.vh"   // this file was generated by the SOCFUSEGEN tool
   
    // --------------------------
    function new( string n="mby_fuse_env", ovm_component p = null);
        super.new( n, p);
    endfunction : new

  
    // --------------------------
    //virtual function void build();
    //  super.build();
    //endfunction : build

  /*
   Function: connect()
   
   In this pahse the user can disbale the defualt constraints on the fuse
   */
   function void connect();
     super.connect();

     //Disable default fuse constraint
     mby_fuse.mby_fuse_mby_fuse_fuse_1.set_default_constraint(0);
   endfunction // void

  
  /*
   constraint: mby_fuse_1_c
   */
   constraint mby_fuse_1_c {
			    mby_fuse.mby_fuse_mby_fuse_fuse_1.cfg_val inside {8'h10,8'h15,8'h34,8'h67,8'hFF};
			    }
 
endclass : mby_fuse_env
