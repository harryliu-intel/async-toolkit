///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_mapper_map_pkg.vh                                  
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_MAPPER_MAP_PKG_VH
`define MBY_PPE_MAPPER_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_mapper_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_mapper_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_mapper_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_mapper_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [38:0] reserved0;  // RSVD
    logic [15:0] DEFAULT_SGLORT;  // RW
    logic  [0:0] DEFAULT_SGLORT_EN;  // RW
    logic  [7:0] PORT_PROFILE;  // RW
} MAP_PORT_CFG_t;

localparam MAP_PORT_CFG_REG_STRIDE = 48'h8;
localparam MAP_PORT_CFG_REG_ENTRIES = 18;
localparam MAP_PORT_CFG_CR_ADDR = 48'h0;
localparam MAP_PORT_CFG_SIZE = 64;
localparam MAP_PORT_CFG_DEFAULT_SGLORT_LO = 9;
localparam MAP_PORT_CFG_DEFAULT_SGLORT_HI = 24;
localparam MAP_PORT_CFG_DEFAULT_SGLORT_RESET = 16'h0;
localparam MAP_PORT_CFG_DEFAULT_SGLORT_EN_LO = 8;
localparam MAP_PORT_CFG_DEFAULT_SGLORT_EN_HI = 8;
localparam MAP_PORT_CFG_DEFAULT_SGLORT_EN_RESET = 1'h0;
localparam MAP_PORT_CFG_PORT_PROFILE_LO = 0;
localparam MAP_PORT_CFG_PORT_PROFILE_HI = 7;
localparam MAP_PORT_CFG_PORT_PROFILE_RESET = 8'h0;
localparam MAP_PORT_CFG_USEMASK = 64'h1FFFFFF;
localparam MAP_PORT_CFG_RO_MASK = 64'h0;
localparam MAP_PORT_CFG_WO_MASK = 64'h0;
localparam MAP_PORT_CFG_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [15:0] VALUE;  // RW
    logic  [7:0] reserved1;  // RSVD
    logic  [7:0] TARGET;  // RW
} MAP_PORT_DEFAULT_t;

localparam MAP_PORT_DEFAULT_REG_STRIDE = 48'h8;
localparam MAP_PORT_DEFAULT_REG_ENTRIES = 6;
localparam MAP_PORT_DEFAULT_REGFILE_STRIDE = 48'h40;
localparam MAP_PORT_DEFAULT_REGFILE_ENTRIES = 18;
localparam MAP_PORT_DEFAULT_CR_ADDR = 48'h200;
localparam MAP_PORT_DEFAULT_SIZE = 64;
localparam MAP_PORT_DEFAULT_VALUE_LO = 16;
localparam MAP_PORT_DEFAULT_VALUE_HI = 31;
localparam MAP_PORT_DEFAULT_VALUE_RESET = 16'h0;
localparam MAP_PORT_DEFAULT_TARGET_LO = 0;
localparam MAP_PORT_DEFAULT_TARGET_HI = 7;
localparam MAP_PORT_DEFAULT_TARGET_RESET = 8'hff;
localparam MAP_PORT_DEFAULT_USEMASK = 64'hFFFF00FF;
localparam MAP_PORT_DEFAULT_RO_MASK = 64'h0;
localparam MAP_PORT_DEFAULT_WO_MASK = 64'h0;
localparam MAP_PORT_DEFAULT_RESET = 64'hFF;

typedef struct packed {
    logic [19:0] reserved0;  // RSVD
    logic [17:0] PORT_KEY_INVERT;  // RW
    logic  [0:0] VID2_VALID_INVERT;  // RW
    logic [11:0] VID2_KEY_INVERT;  // RW
    logic  [0:0] VID1_VALID_INVERT;  // RW
    logic [11:0] VID1_KEY_INVERT;  // RW
    logic [19:0] reserved1;  // RSVD
    logic [17:0] PORT_KEY;  // RW
    logic  [0:0] VID2_VALID;  // RW
    logic [11:0] VID2_KEY;  // RW
    logic  [0:0] VID1_VALID;  // RW
    logic [11:0] VID1_KEY;  // RW
} MAP_DOMAIN_TCAM_t;

localparam MAP_DOMAIN_TCAM_REG_STRIDE = 48'h10;
localparam MAP_DOMAIN_TCAM_REG_ENTRIES = 4096;
localparam MAP_DOMAIN_TCAM_CR_ADDR = 48'h10000;
localparam MAP_DOMAIN_TCAM_SIZE = 128;
localparam MAP_DOMAIN_TCAM_PORT_KEY_INVERT_LO = 90;
localparam MAP_DOMAIN_TCAM_PORT_KEY_INVERT_HI = 107;
localparam MAP_DOMAIN_TCAM_PORT_KEY_INVERT_RESET = 18'h3ffff;
localparam MAP_DOMAIN_TCAM_VID2_VALID_INVERT_LO = 89;
localparam MAP_DOMAIN_TCAM_VID2_VALID_INVERT_HI = 89;
localparam MAP_DOMAIN_TCAM_VID2_VALID_INVERT_RESET = 1'h1;
localparam MAP_DOMAIN_TCAM_VID2_KEY_INVERT_LO = 77;
localparam MAP_DOMAIN_TCAM_VID2_KEY_INVERT_HI = 88;
localparam MAP_DOMAIN_TCAM_VID2_KEY_INVERT_RESET = 12'hfff;
localparam MAP_DOMAIN_TCAM_VID1_VALID_INVERT_LO = 76;
localparam MAP_DOMAIN_TCAM_VID1_VALID_INVERT_HI = 76;
localparam MAP_DOMAIN_TCAM_VID1_VALID_INVERT_RESET = 1'h1;
localparam MAP_DOMAIN_TCAM_VID1_KEY_INVERT_LO = 64;
localparam MAP_DOMAIN_TCAM_VID1_KEY_INVERT_HI = 75;
localparam MAP_DOMAIN_TCAM_VID1_KEY_INVERT_RESET = 12'hfff;
localparam MAP_DOMAIN_TCAM_PORT_KEY_LO = 26;
localparam MAP_DOMAIN_TCAM_PORT_KEY_HI = 43;
localparam MAP_DOMAIN_TCAM_PORT_KEY_RESET = 18'h3ffff;
localparam MAP_DOMAIN_TCAM_VID2_VALID_LO = 25;
localparam MAP_DOMAIN_TCAM_VID2_VALID_HI = 25;
localparam MAP_DOMAIN_TCAM_VID2_VALID_RESET = 1'h1;
localparam MAP_DOMAIN_TCAM_VID2_KEY_LO = 13;
localparam MAP_DOMAIN_TCAM_VID2_KEY_HI = 24;
localparam MAP_DOMAIN_TCAM_VID2_KEY_RESET = 12'hfff;
localparam MAP_DOMAIN_TCAM_VID1_VALID_LO = 12;
localparam MAP_DOMAIN_TCAM_VID1_VALID_HI = 12;
localparam MAP_DOMAIN_TCAM_VID1_VALID_RESET = 1'h1;
localparam MAP_DOMAIN_TCAM_VID1_KEY_LO = 0;
localparam MAP_DOMAIN_TCAM_VID1_KEY_HI = 11;
localparam MAP_DOMAIN_TCAM_VID1_KEY_RESET = 12'hfff;
localparam MAP_DOMAIN_TCAM_USEMASK = 128'hFFFFFFFFFFF00000FFFFFFFFFFF;
localparam MAP_DOMAIN_TCAM_RO_MASK = 128'h0;
localparam MAP_DOMAIN_TCAM_WO_MASK = 128'h0;
localparam MAP_DOMAIN_TCAM_RESET = 128'hFFFFFFFFFFF00000FFFFFFFFFFF;

typedef struct packed {
    logic [25:0] reserved0;  // RSVD
    logic  [7:0] L2_DOMAIN;  // RW
    logic  [5:0] L3_DOMAIN;  // RW
    logic  [3:0] NAD;  // RW
    logic  [0:0] UPDATE_DOMAINS;  // RW
    logic  [0:0] LEARN_EN;  // RW
    logic  [0:0] LEARN_MODE;  // RW
    logic  [4:0] PRIORITY_PROFILE;  // RW
    logic  [7:0] PRI_SOURCE;  // RW
    logic  [0:0] FORCE_DEFAULT_PRI;  // RW
    logic  [2:0] DEFAULT_PRI;  // RW
} MAP_DOMAIN_ACTION0_t;

localparam MAP_DOMAIN_ACTION0_REG_STRIDE = 48'h8;
localparam MAP_DOMAIN_ACTION0_REG_ENTRIES = 4096;
localparam MAP_DOMAIN_ACTION0_CR_ADDR = 48'h20000;
localparam MAP_DOMAIN_ACTION0_SIZE = 64;
localparam MAP_DOMAIN_ACTION0_L2_DOMAIN_LO = 30;
localparam MAP_DOMAIN_ACTION0_L2_DOMAIN_HI = 37;
localparam MAP_DOMAIN_ACTION0_L2_DOMAIN_RESET = 8'h0;
localparam MAP_DOMAIN_ACTION0_L3_DOMAIN_LO = 24;
localparam MAP_DOMAIN_ACTION0_L3_DOMAIN_HI = 29;
localparam MAP_DOMAIN_ACTION0_L3_DOMAIN_RESET = 6'h0;
localparam MAP_DOMAIN_ACTION0_NAD_LO = 20;
localparam MAP_DOMAIN_ACTION0_NAD_HI = 23;
localparam MAP_DOMAIN_ACTION0_NAD_RESET = 4'h0;
localparam MAP_DOMAIN_ACTION0_UPDATE_DOMAINS_LO = 19;
localparam MAP_DOMAIN_ACTION0_UPDATE_DOMAINS_HI = 19;
localparam MAP_DOMAIN_ACTION0_UPDATE_DOMAINS_RESET = 1'h0;
localparam MAP_DOMAIN_ACTION0_LEARN_EN_LO = 18;
localparam MAP_DOMAIN_ACTION0_LEARN_EN_HI = 18;
localparam MAP_DOMAIN_ACTION0_LEARN_EN_RESET = 1'h0;
localparam MAP_DOMAIN_ACTION0_LEARN_MODE_LO = 17;
localparam MAP_DOMAIN_ACTION0_LEARN_MODE_HI = 17;
localparam MAP_DOMAIN_ACTION0_LEARN_MODE_RESET = 1'h0;
localparam MAP_DOMAIN_ACTION0_PRIORITY_PROFILE_LO = 12;
localparam MAP_DOMAIN_ACTION0_PRIORITY_PROFILE_HI = 16;
localparam MAP_DOMAIN_ACTION0_PRIORITY_PROFILE_RESET = 5'h0;
localparam MAP_DOMAIN_ACTION0_PRI_SOURCE_LO = 4;
localparam MAP_DOMAIN_ACTION0_PRI_SOURCE_HI = 11;
localparam MAP_DOMAIN_ACTION0_PRI_SOURCE_RESET = 8'h0;
localparam MAP_DOMAIN_ACTION0_FORCE_DEFAULT_PRI_LO = 3;
localparam MAP_DOMAIN_ACTION0_FORCE_DEFAULT_PRI_HI = 3;
localparam MAP_DOMAIN_ACTION0_FORCE_DEFAULT_PRI_RESET = 1'h0;
localparam MAP_DOMAIN_ACTION0_DEFAULT_PRI_LO = 0;
localparam MAP_DOMAIN_ACTION0_DEFAULT_PRI_HI = 2;
localparam MAP_DOMAIN_ACTION0_DEFAULT_PRI_RESET = 3'h0;
localparam MAP_DOMAIN_ACTION0_USEMASK = 64'h3FFFFFFFFF;
localparam MAP_DOMAIN_ACTION0_RO_MASK = 64'h0;
localparam MAP_DOMAIN_ACTION0_WO_MASK = 64'h0;
localparam MAP_DOMAIN_ACTION0_RESET = 64'h0;

typedef struct packed {
    logic [19:0] reserved0;  // RSVD
    logic  [7:0] DOMAIN_PROFILE;  // RW
    logic [11:0] L2_POLICER;  // RW
    logic [11:0] L3_POLICER;  // RW
    logic [11:0] VLAN_COUNTER;  // RW
} MAP_DOMAIN_ACTION1_t;

localparam MAP_DOMAIN_ACTION1_REG_STRIDE = 48'h8;
localparam MAP_DOMAIN_ACTION1_REG_ENTRIES = 4096;
localparam MAP_DOMAIN_ACTION1_CR_ADDR = 48'h28000;
localparam MAP_DOMAIN_ACTION1_SIZE = 64;
localparam MAP_DOMAIN_ACTION1_DOMAIN_PROFILE_LO = 36;
localparam MAP_DOMAIN_ACTION1_DOMAIN_PROFILE_HI = 43;
localparam MAP_DOMAIN_ACTION1_DOMAIN_PROFILE_RESET = 8'h0;
localparam MAP_DOMAIN_ACTION1_L2_POLICER_LO = 24;
localparam MAP_DOMAIN_ACTION1_L2_POLICER_HI = 35;
localparam MAP_DOMAIN_ACTION1_L2_POLICER_RESET = 12'h0;
localparam MAP_DOMAIN_ACTION1_L3_POLICER_LO = 12;
localparam MAP_DOMAIN_ACTION1_L3_POLICER_HI = 23;
localparam MAP_DOMAIN_ACTION1_L3_POLICER_RESET = 12'h0;
localparam MAP_DOMAIN_ACTION1_VLAN_COUNTER_LO = 0;
localparam MAP_DOMAIN_ACTION1_VLAN_COUNTER_HI = 11;
localparam MAP_DOMAIN_ACTION1_VLAN_COUNTER_RESET = 12'h0;
localparam MAP_DOMAIN_ACTION1_USEMASK = 64'hFFFFFFFFFFF;
localparam MAP_DOMAIN_ACTION1_RO_MASK = 64'h0;
localparam MAP_DOMAIN_ACTION1_WO_MASK = 64'h0;
localparam MAP_DOMAIN_ACTION1_RESET = 64'h0;

typedef struct packed {
    logic [58:0] reserved0;  // RSVD
    logic  [4:0] PRIORITY_PROFILE;  // RW
} MAP_DOMAIN_PROFILE_t;

localparam MAP_DOMAIN_PROFILE_REG_STRIDE = 48'h8;
localparam MAP_DOMAIN_PROFILE_REG_ENTRIES = 256;
localparam MAP_DOMAIN_PROFILE_CR_ADDR = 48'h30000;
localparam MAP_DOMAIN_PROFILE_SIZE = 64;
localparam MAP_DOMAIN_PROFILE_PRIORITY_PROFILE_LO = 0;
localparam MAP_DOMAIN_PROFILE_PRIORITY_PROFILE_HI = 4;
localparam MAP_DOMAIN_PROFILE_PRIORITY_PROFILE_RESET = 5'h0;
localparam MAP_DOMAIN_PROFILE_USEMASK = 64'h1F;
localparam MAP_DOMAIN_PROFILE_RO_MASK = 64'h0;
localparam MAP_DOMAIN_PROFILE_WO_MASK = 64'h0;
localparam MAP_DOMAIN_PROFILE_RESET = 64'h0;

typedef struct packed {
    logic [55:0] reserved0;  // RSVD
    logic  [7:0] MAP_PORT;  // RW
} MAP_PORT_t;

localparam MAP_PORT_REG_STRIDE = 48'h8;
localparam MAP_PORT_REG_ENTRIES = 18;
localparam MAP_PORT_CR_ADDR = 48'h31000;
localparam MAP_PORT_SIZE = 64;
localparam MAP_PORT_MAP_PORT_LO = 0;
localparam MAP_PORT_MAP_PORT_HI = 7;
localparam MAP_PORT_MAP_PORT_RESET = 8'h0;
localparam MAP_PORT_USEMASK = 64'hFF;
localparam MAP_PORT_RO_MASK = 64'h0;
localparam MAP_PORT_WO_MASK = 64'h0;
localparam MAP_PORT_RESET = 64'h0;

typedef struct packed {
    logic [60:0] reserved0;  // RSVD
    logic  [0:0] MAC_ROUTABLE;  // RW
    logic  [7:0] MAP_MAC;  // RW
    logic  [3:0] VALID;  // RW
    logic  [5:0] IGNORE_LENGTH;  // RW
    logic [47:0] MAC;  // RW
} MAP_MAC_t;

localparam MAP_MAC_REG_STRIDE = 48'h10;
localparam MAP_MAC_REG_ENTRIES = 96;
localparam MAP_MAC_CR_ADDR = 48'h31800;
localparam MAP_MAC_SIZE = 128;
localparam MAP_MAC_MAC_ROUTABLE_LO = 66;
localparam MAP_MAC_MAC_ROUTABLE_HI = 66;
localparam MAP_MAC_MAC_ROUTABLE_RESET = 1'h0;
localparam MAP_MAC_MAP_MAC_LO = 58;
localparam MAP_MAC_MAP_MAC_HI = 65;
localparam MAP_MAC_MAP_MAC_RESET = 8'h0;
localparam MAP_MAC_VALID_LO = 54;
localparam MAP_MAC_VALID_HI = 57;
localparam MAP_MAC_VALID_RESET = 4'h0;
localparam MAP_MAC_IGNORE_LENGTH_LO = 48;
localparam MAP_MAC_IGNORE_LENGTH_HI = 53;
localparam MAP_MAC_IGNORE_LENGTH_RESET = 6'h0;
localparam MAP_MAC_MAC_LO = 0;
localparam MAP_MAC_MAC_HI = 47;
localparam MAP_MAC_MAC_RESET = 48'h0;
localparam MAP_MAC_USEMASK = 128'h7FFFFFFFFFFFFFFFF;
localparam MAP_MAC_RO_MASK = 128'h0;
localparam MAP_MAC_WO_MASK = 128'h0;
localparam MAP_MAC_RESET = 128'h0;

typedef struct packed {
    logic [63:0] IP_LO;  // RW
} MAP_IP_LO_t;

localparam MAP_IP_LO_REG_STRIDE = 48'h8;
localparam MAP_IP_LO_REG_ENTRIES = 16;
localparam MAP_IP_LO_CR_ADDR = 48'h32080;
localparam MAP_IP_LO_SIZE = 64;
localparam MAP_IP_LO_IP_LO_LO = 0;
localparam MAP_IP_LO_IP_LO_HI = 63;
localparam MAP_IP_LO_IP_LO_RESET = 64'h0;
localparam MAP_IP_LO_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam MAP_IP_LO_RO_MASK = 64'h0;
localparam MAP_IP_LO_WO_MASK = 64'h0;
localparam MAP_IP_LO_RESET = 64'h0;

typedef struct packed {
    logic [63:0] IP_HI;  // RW
} MAP_IP_HI_t;

localparam MAP_IP_HI_REG_STRIDE = 48'h8;
localparam MAP_IP_HI_REG_ENTRIES = 16;
localparam MAP_IP_HI_CR_ADDR = 48'h32100;
localparam MAP_IP_HI_SIZE = 64;
localparam MAP_IP_HI_IP_HI_LO = 0;
localparam MAP_IP_HI_IP_HI_HI = 63;
localparam MAP_IP_HI_IP_HI_RESET = 64'h0;
localparam MAP_IP_HI_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam MAP_IP_HI_RO_MASK = 64'h0;
localparam MAP_IP_HI_WO_MASK = 64'h0;
localparam MAP_IP_HI_RESET = 64'h0;

typedef struct packed {
    logic [44:0] reserved0;  // RSVD
    logic  [7:0] MATCH_LENGTH;  // RW
    logic  [3:0] VALID;  // RW
    logic  [3:0] MAP_IP;  // RW
    logic  [1:0] IP_PROFILE;  // RW
    logic  [0:0] IS_IPV6;  // RW
} MAP_IP_CFG_t;

localparam MAP_IP_CFG_REG_STRIDE = 48'h8;
localparam MAP_IP_CFG_REG_ENTRIES = 16;
localparam MAP_IP_CFG_CR_ADDR = 48'h32180;
localparam MAP_IP_CFG_SIZE = 64;
localparam MAP_IP_CFG_MATCH_LENGTH_LO = 11;
localparam MAP_IP_CFG_MATCH_LENGTH_HI = 18;
localparam MAP_IP_CFG_MATCH_LENGTH_RESET = 8'h0;
localparam MAP_IP_CFG_VALID_LO = 7;
localparam MAP_IP_CFG_VALID_HI = 10;
localparam MAP_IP_CFG_VALID_RESET = 4'h0;
localparam MAP_IP_CFG_MAP_IP_LO = 3;
localparam MAP_IP_CFG_MAP_IP_HI = 6;
localparam MAP_IP_CFG_MAP_IP_RESET = 4'h0;
localparam MAP_IP_CFG_IP_PROFILE_LO = 1;
localparam MAP_IP_CFG_IP_PROFILE_HI = 2;
localparam MAP_IP_CFG_IP_PROFILE_RESET = 2'h0;
localparam MAP_IP_CFG_IS_IPV6_LO = 0;
localparam MAP_IP_CFG_IS_IPV6_HI = 0;
localparam MAP_IP_CFG_IS_IPV6_RESET = 1'h0;
localparam MAP_IP_CFG_USEMASK = 64'h7FFFF;
localparam MAP_IP_CFG_RO_MASK = 64'h0;
localparam MAP_IP_CFG_WO_MASK = 64'h0;
localparam MAP_IP_CFG_RESET = 64'h0;

typedef struct packed {
    logic [52:0] reserved0;  // RSVD
    logic  [2:0] MAP_PROT;  // RW
    logic  [7:0] PROT;  // RW
} MAP_PROT_t;

localparam MAP_PROT_REG_STRIDE = 48'h8;
localparam MAP_PROT_REG_ENTRIES = 8;
localparam MAP_PROT_CR_ADDR = 48'h32200;
localparam MAP_PROT_SIZE = 64;
localparam MAP_PROT_MAP_PROT_LO = 8;
localparam MAP_PROT_MAP_PROT_HI = 10;
localparam MAP_PROT_MAP_PROT_RESET = 3'h0;
localparam MAP_PROT_PROT_LO = 0;
localparam MAP_PROT_PROT_HI = 7;
localparam MAP_PROT_PROT_RESET = 8'h0;
localparam MAP_PROT_USEMASK = 64'h7FF;
localparam MAP_PROT_RO_MASK = 64'h0;
localparam MAP_PROT_WO_MASK = 64'h0;
localparam MAP_PROT_RESET = 64'h0;

typedef struct packed {
    logic [26:0] reserved0;  // RSVD
    logic [15:0] MAP_L4_SRC;  // RW
    logic  [1:0] VALID;  // RW
    logic  [2:0] MAP_PROT;  // RW
    logic [15:0] L4_SRC;  // RW
} MAP_L4_SRC_t;

localparam MAP_L4_SRC_REG_STRIDE = 48'h8;
localparam MAP_L4_SRC_REG_ENTRIES = 64;
localparam MAP_L4_SRC_CR_ADDR = 48'h32400;
localparam MAP_L4_SRC_SIZE = 64;
localparam MAP_L4_SRC_MAP_L4_SRC_LO = 21;
localparam MAP_L4_SRC_MAP_L4_SRC_HI = 36;
localparam MAP_L4_SRC_MAP_L4_SRC_RESET = 16'h0;
localparam MAP_L4_SRC_VALID_LO = 19;
localparam MAP_L4_SRC_VALID_HI = 20;
localparam MAP_L4_SRC_VALID_RESET = 2'h0;
localparam MAP_L4_SRC_MAP_PROT_LO = 16;
localparam MAP_L4_SRC_MAP_PROT_HI = 18;
localparam MAP_L4_SRC_MAP_PROT_RESET = 3'h0;
localparam MAP_L4_SRC_L4_SRC_LO = 0;
localparam MAP_L4_SRC_L4_SRC_HI = 15;
localparam MAP_L4_SRC_L4_SRC_RESET = 16'h0;
localparam MAP_L4_SRC_USEMASK = 64'h1FFFFFFFFF;
localparam MAP_L4_SRC_RO_MASK = 64'h0;
localparam MAP_L4_SRC_WO_MASK = 64'h0;
localparam MAP_L4_SRC_RESET = 64'h0;

typedef struct packed {
    logic [26:0] reserved0;  // RSVD
    logic [15:0] MAP_L4_DST;  // RW
    logic  [1:0] VALID;  // RW
    logic  [2:0] MAP_PROT;  // RW
    logic [15:0] L4_DST;  // RW
} MAP_L4_DST_t;

localparam MAP_L4_DST_REG_STRIDE = 48'h8;
localparam MAP_L4_DST_REG_ENTRIES = 64;
localparam MAP_L4_DST_CR_ADDR = 48'h32600;
localparam MAP_L4_DST_SIZE = 64;
localparam MAP_L4_DST_MAP_L4_DST_LO = 21;
localparam MAP_L4_DST_MAP_L4_DST_HI = 36;
localparam MAP_L4_DST_MAP_L4_DST_RESET = 16'h0;
localparam MAP_L4_DST_VALID_LO = 19;
localparam MAP_L4_DST_VALID_HI = 20;
localparam MAP_L4_DST_VALID_RESET = 2'h0;
localparam MAP_L4_DST_MAP_PROT_LO = 16;
localparam MAP_L4_DST_MAP_PROT_HI = 18;
localparam MAP_L4_DST_MAP_PROT_RESET = 3'h0;
localparam MAP_L4_DST_L4_DST_LO = 0;
localparam MAP_L4_DST_L4_DST_HI = 15;
localparam MAP_L4_DST_L4_DST_RESET = 16'h0;
localparam MAP_L4_DST_USEMASK = 64'h1FFFFFFFFF;
localparam MAP_L4_DST_RO_MASK = 64'h0;
localparam MAP_L4_DST_WO_MASK = 64'h0;
localparam MAP_L4_DST_RESET = 64'h0;

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic [23:0] TC_BY_EXP;  // RW
} MAP_EXP_TC_t;

localparam MAP_EXP_TC_REG_STRIDE = 48'h8;
localparam MAP_EXP_TC_REG_ENTRIES = 32;
localparam MAP_EXP_TC_CR_ADDR = 48'h32800;
localparam MAP_EXP_TC_SIZE = 64;
localparam MAP_EXP_TC_TC_BY_EXP_LO = 0;
localparam MAP_EXP_TC_TC_BY_EXP_HI = 23;
localparam MAP_EXP_TC_TC_BY_EXP_RESET = 'h0;
localparam MAP_EXP_TC_USEMASK = 64'hFFFFFF;
localparam MAP_EXP_TC_RO_MASK = 64'h0;
localparam MAP_EXP_TC_WO_MASK = 64'h0;
localparam MAP_EXP_TC_RESET = 64'h0;

typedef struct packed {
    logic [54:0] reserved0;  // RSVD
    logic  [2:0] TC;  // RW
    logic  [5:0] DSCP;  // RW
} MAP_DSCP_TC_t;

localparam MAP_DSCP_TC_REG_STRIDE = 48'h8;
localparam MAP_DSCP_TC_REG_ENTRIES = 2048;
localparam MAP_DSCP_TC_CR_ADDR = 48'h34000;
localparam MAP_DSCP_TC_SIZE = 64;
localparam MAP_DSCP_TC_TC_LO = 6;
localparam MAP_DSCP_TC_TC_HI = 8;
localparam MAP_DSCP_TC_TC_RESET = 3'h0;
localparam MAP_DSCP_TC_DSCP_LO = 0;
localparam MAP_DSCP_TC_DSCP_HI = 5;
localparam MAP_DSCP_TC_DSCP_RESET = 6'h0;
localparam MAP_DSCP_TC_USEMASK = 64'h1FF;
localparam MAP_DSCP_TC_RO_MASK = 64'h0;
localparam MAP_DSCP_TC_WO_MASK = 64'h0;
localparam MAP_DSCP_TC_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] TC_BY_VPRI;  // RW
} MAP_VPRI_TC_t;

localparam MAP_VPRI_TC_REG_STRIDE = 48'h8;
localparam MAP_VPRI_TC_REG_ENTRIES = 32;
localparam MAP_VPRI_TC_CR_ADDR = 48'h38000;
localparam MAP_VPRI_TC_SIZE = 64;
localparam MAP_VPRI_TC_TC_BY_VPRI_LO = 0;
localparam MAP_VPRI_TC_TC_BY_VPRI_HI = 47;
localparam MAP_VPRI_TC_TC_BY_VPRI_RESET = 'h0;
localparam MAP_VPRI_TC_USEMASK = 64'hFFFFFFFFFFFF;
localparam MAP_VPRI_TC_RO_MASK = 64'h0;
localparam MAP_VPRI_TC_WO_MASK = 64'h0;
localparam MAP_VPRI_TC_RESET = 64'h0;

typedef struct packed {
    logic [63:0] VPRI_BY_VPRI;  // RW
} MAP_VPRI_t;

localparam MAP_VPRI_REG_STRIDE = 48'h8;
localparam MAP_VPRI_REG_ENTRIES = 32;
localparam MAP_VPRI_CR_ADDR = 48'h38100;
localparam MAP_VPRI_SIZE = 64;
localparam MAP_VPRI_VPRI_BY_VPRI_LO = 0;
localparam MAP_VPRI_VPRI_BY_VPRI_HI = 63;
localparam MAP_VPRI_VPRI_BY_VPRI_RESET = 'h0;
localparam MAP_VPRI_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam MAP_VPRI_RO_MASK = 64'h0;
localparam MAP_VPRI_WO_MASK = 64'h0;
localparam MAP_VPRI_RESET = 64'h0;

typedef struct packed {
    logic  [3:0] reserved0;  // RSVD
    logic  [0:0] PTRS_ERR;  // RW
    logic  [2:0] EX;  // RW
    logic  [1:0] CSUM;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [0:0] IHL_OK;  // RW
    logic  [0:0] IHL_FITS;  // RW
    logic [46:0] FLAGS;  // RW
    logic  [0:0] RSVD;  // RW
} MAP_PROFILE_KEY0_t;

localparam MAP_PROFILE_KEY0_REG_STRIDE = 48'h8;
localparam MAP_PROFILE_KEY0_REG_ENTRIES = 96;
localparam MAP_PROFILE_KEY0_CR_ADDR = 48'h38400;
localparam MAP_PROFILE_KEY0_SIZE = 64;
localparam MAP_PROFILE_KEY0_PTRS_ERR_LO = 59;
localparam MAP_PROFILE_KEY0_PTRS_ERR_HI = 59;
localparam MAP_PROFILE_KEY0_PTRS_ERR_RESET = 1'h1;
localparam MAP_PROFILE_KEY0_EX_LO = 56;
localparam MAP_PROFILE_KEY0_EX_HI = 58;
localparam MAP_PROFILE_KEY0_EX_RESET = 3'h7;
localparam MAP_PROFILE_KEY0_CSUM_LO = 54;
localparam MAP_PROFILE_KEY0_CSUM_HI = 55;
localparam MAP_PROFILE_KEY0_CSUM_RESET = 2'h3;
localparam MAP_PROFILE_KEY0_IHL_OK_LO = 49;
localparam MAP_PROFILE_KEY0_IHL_OK_HI = 49;
localparam MAP_PROFILE_KEY0_IHL_OK_RESET = 1'h1;
localparam MAP_PROFILE_KEY0_IHL_FITS_LO = 48;
localparam MAP_PROFILE_KEY0_IHL_FITS_HI = 48;
localparam MAP_PROFILE_KEY0_IHL_FITS_RESET = 1'h1;
localparam MAP_PROFILE_KEY0_FLAGS_LO = 1;
localparam MAP_PROFILE_KEY0_FLAGS_HI = 47;
localparam MAP_PROFILE_KEY0_FLAGS_RESET = 47'h7fffffffffff;
localparam MAP_PROFILE_KEY0_RSVD_LO = 0;
localparam MAP_PROFILE_KEY0_RSVD_HI = 0;
localparam MAP_PROFILE_KEY0_RSVD_RESET = 1'h1;
localparam MAP_PROFILE_KEY0_USEMASK = 64'hFC3FFFFFFFFFFFF;
localparam MAP_PROFILE_KEY0_RO_MASK = 64'h0;
localparam MAP_PROFILE_KEY0_WO_MASK = 64'h0;
localparam MAP_PROFILE_KEY0_RESET = 64'hFC3FFFFFFFFFFFF;

typedef struct packed {
    logic  [3:0] reserved0;  // RSVD
    logic  [0:0] PTRS_ERR;  // RW
    logic  [2:0] EX;  // RW
    logic  [1:0] CSUM;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [0:0] IHL_OK;  // RW
    logic  [0:0] IHL_FITS;  // RW
    logic [46:0] FLAGS;  // RW
    logic  [0:0] RSVD;  // RW
} MAP_PROFILE_KEY_INVERT0_t;

localparam MAP_PROFILE_KEY_INVERT0_REG_STRIDE = 48'h8;
localparam MAP_PROFILE_KEY_INVERT0_REG_ENTRIES = 96;
localparam MAP_PROFILE_KEY_INVERT0_CR_ADDR = 48'h38800;
localparam MAP_PROFILE_KEY_INVERT0_SIZE = 64;
localparam MAP_PROFILE_KEY_INVERT0_PTRS_ERR_LO = 59;
localparam MAP_PROFILE_KEY_INVERT0_PTRS_ERR_HI = 59;
localparam MAP_PROFILE_KEY_INVERT0_PTRS_ERR_RESET = 1'h1;
localparam MAP_PROFILE_KEY_INVERT0_EX_LO = 56;
localparam MAP_PROFILE_KEY_INVERT0_EX_HI = 58;
localparam MAP_PROFILE_KEY_INVERT0_EX_RESET = 3'h7;
localparam MAP_PROFILE_KEY_INVERT0_CSUM_LO = 54;
localparam MAP_PROFILE_KEY_INVERT0_CSUM_HI = 55;
localparam MAP_PROFILE_KEY_INVERT0_CSUM_RESET = 2'h3;
localparam MAP_PROFILE_KEY_INVERT0_IHL_OK_LO = 49;
localparam MAP_PROFILE_KEY_INVERT0_IHL_OK_HI = 49;
localparam MAP_PROFILE_KEY_INVERT0_IHL_OK_RESET = 1'h1;
localparam MAP_PROFILE_KEY_INVERT0_IHL_FITS_LO = 48;
localparam MAP_PROFILE_KEY_INVERT0_IHL_FITS_HI = 48;
localparam MAP_PROFILE_KEY_INVERT0_IHL_FITS_RESET = 1'h1;
localparam MAP_PROFILE_KEY_INVERT0_FLAGS_LO = 1;
localparam MAP_PROFILE_KEY_INVERT0_FLAGS_HI = 47;
localparam MAP_PROFILE_KEY_INVERT0_FLAGS_RESET = 47'h7fffffffffff;
localparam MAP_PROFILE_KEY_INVERT0_RSVD_LO = 0;
localparam MAP_PROFILE_KEY_INVERT0_RSVD_HI = 0;
localparam MAP_PROFILE_KEY_INVERT0_RSVD_RESET = 1'h1;
localparam MAP_PROFILE_KEY_INVERT0_USEMASK = 64'hFC3FFFFFFFFFFFF;
localparam MAP_PROFILE_KEY_INVERT0_RO_MASK = 64'h0;
localparam MAP_PROFILE_KEY_INVERT0_WO_MASK = 64'h0;
localparam MAP_PROFILE_KEY_INVERT0_RESET = 64'hFC3FFFFFFFFFFFF;

typedef struct packed {
    logic [13:0] reserved0;  // RSVD
    logic  [9:0] PTYPE;  // RW
    logic  [7:0] L2_DOMAIN;  // RW
    logic  [5:0] L3_DOMAIN;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [7:0] PORT_PROFILE;  // RW
    logic  [7:0] DOMAIN_PROFILE;  // RW
    logic  [3:0] MAC_ROUTABLE;  // RW
    logic  [1:0] MAC_MBCAST;  // RW
} MAP_PROFILE_KEY1_t;

localparam MAP_PROFILE_KEY1_REG_STRIDE = 48'h8;
localparam MAP_PROFILE_KEY1_REG_ENTRIES = 96;
localparam MAP_PROFILE_KEY1_CR_ADDR = 48'h38C00;
localparam MAP_PROFILE_KEY1_SIZE = 64;
localparam MAP_PROFILE_KEY1_PTYPE_LO = 40;
localparam MAP_PROFILE_KEY1_PTYPE_HI = 49;
localparam MAP_PROFILE_KEY1_PTYPE_RESET = 10'h0;
localparam MAP_PROFILE_KEY1_L2_DOMAIN_LO = 32;
localparam MAP_PROFILE_KEY1_L2_DOMAIN_HI = 39;
localparam MAP_PROFILE_KEY1_L2_DOMAIN_RESET = 8'hff;
localparam MAP_PROFILE_KEY1_L3_DOMAIN_LO = 26;
localparam MAP_PROFILE_KEY1_L3_DOMAIN_HI = 31;
localparam MAP_PROFILE_KEY1_L3_DOMAIN_RESET = 6'h3f;
localparam MAP_PROFILE_KEY1_PORT_PROFILE_LO = 14;
localparam MAP_PROFILE_KEY1_PORT_PROFILE_HI = 21;
localparam MAP_PROFILE_KEY1_PORT_PROFILE_RESET = 8'hff;
localparam MAP_PROFILE_KEY1_DOMAIN_PROFILE_LO = 6;
localparam MAP_PROFILE_KEY1_DOMAIN_PROFILE_HI = 13;
localparam MAP_PROFILE_KEY1_DOMAIN_PROFILE_RESET = 8'hff;
localparam MAP_PROFILE_KEY1_MAC_ROUTABLE_LO = 2;
localparam MAP_PROFILE_KEY1_MAC_ROUTABLE_HI = 5;
localparam MAP_PROFILE_KEY1_MAC_ROUTABLE_RESET = 4'hf;
localparam MAP_PROFILE_KEY1_MAC_MBCAST_LO = 0;
localparam MAP_PROFILE_KEY1_MAC_MBCAST_HI = 1;
localparam MAP_PROFILE_KEY1_MAC_MBCAST_RESET = 2'h3;
localparam MAP_PROFILE_KEY1_USEMASK = 64'h3FFFFFC3FFFFF;
localparam MAP_PROFILE_KEY1_RO_MASK = 64'h0;
localparam MAP_PROFILE_KEY1_WO_MASK = 64'h0;
localparam MAP_PROFILE_KEY1_RESET = 64'hFFFC3FFFFF;

typedef struct packed {
    logic [13:0] reserved0;  // RSVD
    logic  [9:0] PTYPE;  // RW
    logic  [7:0] L2_DOMAIN;  // RW
    logic  [5:0] L3_DOMAIN;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [7:0] PORT_PROFILE;  // RW
    logic  [7:0] DOMAIN_PROFILE;  // RW
    logic  [3:0] MAC_ROUTABLE;  // RW
    logic  [1:0] MAC_MBCAST;  // RW
} MAP_PROFILE_KEY_INVERT1_t;

localparam MAP_PROFILE_KEY_INVERT1_REG_STRIDE = 48'h8;
localparam MAP_PROFILE_KEY_INVERT1_REG_ENTRIES = 96;
localparam MAP_PROFILE_KEY_INVERT1_CR_ADDR = 48'h39000;
localparam MAP_PROFILE_KEY_INVERT1_SIZE = 64;
localparam MAP_PROFILE_KEY_INVERT1_PTYPE_LO = 40;
localparam MAP_PROFILE_KEY_INVERT1_PTYPE_HI = 49;
localparam MAP_PROFILE_KEY_INVERT1_PTYPE_RESET = 10'h0;
localparam MAP_PROFILE_KEY_INVERT1_L2_DOMAIN_LO = 32;
localparam MAP_PROFILE_KEY_INVERT1_L2_DOMAIN_HI = 39;
localparam MAP_PROFILE_KEY_INVERT1_L2_DOMAIN_RESET = 8'hff;
localparam MAP_PROFILE_KEY_INVERT1_L3_DOMAIN_LO = 26;
localparam MAP_PROFILE_KEY_INVERT1_L3_DOMAIN_HI = 31;
localparam MAP_PROFILE_KEY_INVERT1_L3_DOMAIN_RESET = 6'h3f;
localparam MAP_PROFILE_KEY_INVERT1_PORT_PROFILE_LO = 14;
localparam MAP_PROFILE_KEY_INVERT1_PORT_PROFILE_HI = 21;
localparam MAP_PROFILE_KEY_INVERT1_PORT_PROFILE_RESET = 8'hff;
localparam MAP_PROFILE_KEY_INVERT1_DOMAIN_PROFILE_LO = 6;
localparam MAP_PROFILE_KEY_INVERT1_DOMAIN_PROFILE_HI = 13;
localparam MAP_PROFILE_KEY_INVERT1_DOMAIN_PROFILE_RESET = 8'hff;
localparam MAP_PROFILE_KEY_INVERT1_MAC_ROUTABLE_LO = 2;
localparam MAP_PROFILE_KEY_INVERT1_MAC_ROUTABLE_HI = 5;
localparam MAP_PROFILE_KEY_INVERT1_MAC_ROUTABLE_RESET = 4'hf;
localparam MAP_PROFILE_KEY_INVERT1_MAC_MBCAST_LO = 0;
localparam MAP_PROFILE_KEY_INVERT1_MAC_MBCAST_HI = 1;
localparam MAP_PROFILE_KEY_INVERT1_MAC_MBCAST_RESET = 2'h3;
localparam MAP_PROFILE_KEY_INVERT1_USEMASK = 64'h3FFFFFC3FFFFF;
localparam MAP_PROFILE_KEY_INVERT1_RO_MASK = 64'h0;
localparam MAP_PROFILE_KEY_INVERT1_WO_MASK = 64'h0;
localparam MAP_PROFILE_KEY_INVERT1_RESET = 64'hFFFC3FFFFF;

typedef struct packed {
    logic [28:0] reserved0;  // RSVD
    logic  [0:0] PROFILE_VALID;  // RW
    logic  [5:0] PROFILE;  // RW
    logic  [3:0] REWRITE_PROFILE;  // RW
    logic  [0:0] TRIG_VALID;  // RW
    logic  [7:0] PROFILE_TRIG;  // RW
    logic  [0:0] PARSER_ERROR;  // RW
    logic  [6:0] IP_OPTIONS_MASK;  // RW
    logic  [0:0] PRIOS_VALID;  // RW
    logic  [2:0] VPRI_TGT;  // RW
    logic  [2:0] DSCP_TGT;  // RW
} MAP_PROFILE_ACTION_t;

localparam MAP_PROFILE_ACTION_REG_STRIDE = 48'h8;
localparam MAP_PROFILE_ACTION_REG_ENTRIES = 96;
localparam MAP_PROFILE_ACTION_CR_ADDR = 48'h39400;
localparam MAP_PROFILE_ACTION_SIZE = 64;
localparam MAP_PROFILE_ACTION_PROFILE_VALID_LO = 34;
localparam MAP_PROFILE_ACTION_PROFILE_VALID_HI = 34;
localparam MAP_PROFILE_ACTION_PROFILE_VALID_RESET = 1'h0;
localparam MAP_PROFILE_ACTION_PROFILE_LO = 28;
localparam MAP_PROFILE_ACTION_PROFILE_HI = 33;
localparam MAP_PROFILE_ACTION_PROFILE_RESET = 6'h0;
localparam MAP_PROFILE_ACTION_REWRITE_PROFILE_LO = 24;
localparam MAP_PROFILE_ACTION_REWRITE_PROFILE_HI = 27;
localparam MAP_PROFILE_ACTION_REWRITE_PROFILE_RESET = 4'h0;
localparam MAP_PROFILE_ACTION_TRIG_VALID_LO = 23;
localparam MAP_PROFILE_ACTION_TRIG_VALID_HI = 23;
localparam MAP_PROFILE_ACTION_TRIG_VALID_RESET = 1'h0;
localparam MAP_PROFILE_ACTION_PROFILE_TRIG_LO = 15;
localparam MAP_PROFILE_ACTION_PROFILE_TRIG_HI = 22;
localparam MAP_PROFILE_ACTION_PROFILE_TRIG_RESET = 8'h0;
localparam MAP_PROFILE_ACTION_PARSER_ERROR_LO = 14;
localparam MAP_PROFILE_ACTION_PARSER_ERROR_HI = 14;
localparam MAP_PROFILE_ACTION_PARSER_ERROR_RESET = 1'h0;
localparam MAP_PROFILE_ACTION_IP_OPTIONS_MASK_LO = 7;
localparam MAP_PROFILE_ACTION_IP_OPTIONS_MASK_HI = 13;
localparam MAP_PROFILE_ACTION_IP_OPTIONS_MASK_RESET = 7'h0;
localparam MAP_PROFILE_ACTION_PRIOS_VALID_LO = 6;
localparam MAP_PROFILE_ACTION_PRIOS_VALID_HI = 6;
localparam MAP_PROFILE_ACTION_PRIOS_VALID_RESET = 1'h0;
localparam MAP_PROFILE_ACTION_VPRI_TGT_LO = 3;
localparam MAP_PROFILE_ACTION_VPRI_TGT_HI = 5;
localparam MAP_PROFILE_ACTION_VPRI_TGT_RESET = 3'h0;
localparam MAP_PROFILE_ACTION_DSCP_TGT_LO = 0;
localparam MAP_PROFILE_ACTION_DSCP_TGT_HI = 2;
localparam MAP_PROFILE_ACTION_DSCP_TGT_RESET = 3'h0;
localparam MAP_PROFILE_ACTION_USEMASK = 64'h7FFFFFFFF;
localparam MAP_PROFILE_ACTION_RO_MASK = 64'h0;
localparam MAP_PROFILE_ACTION_WO_MASK = 64'h0;
localparam MAP_PROFILE_ACTION_RESET = 64'h0;

typedef struct packed {
    logic [57:0] reserved0;  // RSVD
    logic  [2:0] L3_COLOR_CFG;  // RW
    logic  [2:0] L2_COLOR_CFG;  // RW
} MAP_DOMAIN_POL_CFG_t;

localparam MAP_DOMAIN_POL_CFG_REG_STRIDE = 48'h8;
localparam MAP_DOMAIN_POL_CFG_REG_ENTRIES = 1;
localparam MAP_DOMAIN_POL_CFG_CR_ADDR = 48'h39800;
localparam MAP_DOMAIN_POL_CFG_SIZE = 64;
localparam MAP_DOMAIN_POL_CFG_L3_COLOR_CFG_LO = 3;
localparam MAP_DOMAIN_POL_CFG_L3_COLOR_CFG_HI = 5;
localparam MAP_DOMAIN_POL_CFG_L3_COLOR_CFG_RESET = 3'h0;
localparam MAP_DOMAIN_POL_CFG_L2_COLOR_CFG_LO = 0;
localparam MAP_DOMAIN_POL_CFG_L2_COLOR_CFG_HI = 2;
localparam MAP_DOMAIN_POL_CFG_L2_COLOR_CFG_RESET = 3'h0;
localparam MAP_DOMAIN_POL_CFG_USEMASK = 64'h3F;
localparam MAP_DOMAIN_POL_CFG_RO_MASK = 64'h0;
localparam MAP_DOMAIN_POL_CFG_WO_MASK = 64'h0;
localparam MAP_DOMAIN_POL_CFG_RESET = 64'h0;

typedef struct packed {
    logic [57:0] reserved0;  // RSVD
    logic  [5:0] SRC_ID;  // RW
} MAP_REWRITE_t;

localparam MAP_REWRITE_REG_STRIDE = 48'h8;
localparam MAP_REWRITE_REG_ENTRIES = 32;
localparam MAP_REWRITE_REGFILE_STRIDE = 48'h100;
localparam MAP_REWRITE_REGFILE_ENTRIES = 16;
localparam MAP_REWRITE_CR_ADDR = 48'h3A000;
localparam MAP_REWRITE_SIZE = 64;
localparam MAP_REWRITE_SRC_ID_LO = 0;
localparam MAP_REWRITE_SRC_ID_HI = 5;
localparam MAP_REWRITE_SRC_ID_RESET = 6'h0;
localparam MAP_REWRITE_USEMASK = 64'h3F;
localparam MAP_REWRITE_RO_MASK = 64'h0;
localparam MAP_REWRITE_WO_MASK = 64'h0;
localparam MAP_REWRITE_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_MAP_PORT_CFG_t;

typedef logic [7:0] we_MAP_PORT_DEFAULT_t;

typedef logic [15:0] we_MAP_DOMAIN_TCAM_t;

typedef logic [7:0] we_MAP_DOMAIN_ACTION0_t;

typedef logic [7:0] we_MAP_DOMAIN_ACTION1_t;

typedef logic [7:0] we_MAP_DOMAIN_PROFILE_t;

typedef logic [7:0] we_MAP_PORT_t;

typedef logic [15:0] we_MAP_MAC_t;

typedef logic [7:0] we_MAP_IP_LO_t;

typedef logic [7:0] we_MAP_IP_HI_t;

typedef logic [7:0] we_MAP_IP_CFG_t;

typedef logic [7:0] we_MAP_PROT_t;

typedef logic [7:0] we_MAP_L4_SRC_t;

typedef logic [7:0] we_MAP_L4_DST_t;

typedef logic [7:0] we_MAP_EXP_TC_t;

typedef logic [7:0] we_MAP_DSCP_TC_t;

typedef logic [7:0] we_MAP_VPRI_TC_t;

typedef logic [7:0] we_MAP_VPRI_t;

typedef logic [7:0] we_MAP_PROFILE_KEY0_t;

typedef logic [7:0] we_MAP_PROFILE_KEY_INVERT0_t;

typedef logic [7:0] we_MAP_PROFILE_KEY1_t;

typedef logic [7:0] we_MAP_PROFILE_KEY_INVERT1_t;

typedef logic [7:0] we_MAP_PROFILE_ACTION_t;

typedef logic [7:0] we_MAP_DOMAIN_POL_CFG_t;

typedef logic [7:0] we_MAP_REWRITE_t;

typedef struct packed {
    we_MAP_PORT_CFG_t MAP_PORT_CFG;
    we_MAP_PORT_DEFAULT_t MAP_PORT_DEFAULT;
    we_MAP_DOMAIN_TCAM_t MAP_DOMAIN_TCAM;
    we_MAP_DOMAIN_ACTION0_t MAP_DOMAIN_ACTION0;
    we_MAP_DOMAIN_ACTION1_t MAP_DOMAIN_ACTION1;
    we_MAP_DOMAIN_PROFILE_t MAP_DOMAIN_PROFILE;
    we_MAP_PORT_t MAP_PORT;
    we_MAP_MAC_t MAP_MAC;
    we_MAP_IP_LO_t MAP_IP_LO;
    we_MAP_IP_HI_t MAP_IP_HI;
    we_MAP_IP_CFG_t MAP_IP_CFG;
    we_MAP_PROT_t MAP_PROT;
    we_MAP_L4_SRC_t MAP_L4_SRC;
    we_MAP_L4_DST_t MAP_L4_DST;
    we_MAP_EXP_TC_t MAP_EXP_TC;
    we_MAP_DSCP_TC_t MAP_DSCP_TC;
    we_MAP_VPRI_TC_t MAP_VPRI_TC;
    we_MAP_VPRI_t MAP_VPRI;
    we_MAP_PROFILE_KEY0_t MAP_PROFILE_KEY0;
    we_MAP_PROFILE_KEY_INVERT0_t MAP_PROFILE_KEY_INVERT0;
    we_MAP_PROFILE_KEY1_t MAP_PROFILE_KEY1;
    we_MAP_PROFILE_KEY_INVERT1_t MAP_PROFILE_KEY_INVERT1;
    we_MAP_PROFILE_ACTION_t MAP_PROFILE_ACTION;
    we_MAP_DOMAIN_POL_CFG_t MAP_DOMAIN_POL_CFG;
    we_MAP_REWRITE_t MAP_REWRITE;
} mby_ppe_mapper_map_handcoded_t;

typedef logic [7:0] re_MAP_PORT_CFG_t;

typedef logic [7:0] re_MAP_PORT_DEFAULT_t;

typedef logic [15:0] re_MAP_DOMAIN_TCAM_t;

typedef logic [7:0] re_MAP_DOMAIN_ACTION0_t;

typedef logic [7:0] re_MAP_DOMAIN_ACTION1_t;

typedef logic [7:0] re_MAP_DOMAIN_PROFILE_t;

typedef logic [7:0] re_MAP_PORT_t;

typedef logic [15:0] re_MAP_MAC_t;

typedef logic [7:0] re_MAP_IP_LO_t;

typedef logic [7:0] re_MAP_IP_HI_t;

typedef logic [7:0] re_MAP_IP_CFG_t;

typedef logic [7:0] re_MAP_PROT_t;

typedef logic [7:0] re_MAP_L4_SRC_t;

typedef logic [7:0] re_MAP_L4_DST_t;

typedef logic [7:0] re_MAP_EXP_TC_t;

typedef logic [7:0] re_MAP_DSCP_TC_t;

typedef logic [7:0] re_MAP_VPRI_TC_t;

typedef logic [7:0] re_MAP_VPRI_t;

typedef logic [7:0] re_MAP_PROFILE_KEY0_t;

typedef logic [7:0] re_MAP_PROFILE_KEY_INVERT0_t;

typedef logic [7:0] re_MAP_PROFILE_KEY1_t;

typedef logic [7:0] re_MAP_PROFILE_KEY_INVERT1_t;

typedef logic [7:0] re_MAP_PROFILE_ACTION_t;

typedef logic [7:0] re_MAP_DOMAIN_POL_CFG_t;

typedef logic [7:0] re_MAP_REWRITE_t;

typedef struct packed {
    re_MAP_PORT_CFG_t MAP_PORT_CFG;
    re_MAP_PORT_DEFAULT_t MAP_PORT_DEFAULT;
    re_MAP_DOMAIN_TCAM_t MAP_DOMAIN_TCAM;
    re_MAP_DOMAIN_ACTION0_t MAP_DOMAIN_ACTION0;
    re_MAP_DOMAIN_ACTION1_t MAP_DOMAIN_ACTION1;
    re_MAP_DOMAIN_PROFILE_t MAP_DOMAIN_PROFILE;
    re_MAP_PORT_t MAP_PORT;
    re_MAP_MAC_t MAP_MAC;
    re_MAP_IP_LO_t MAP_IP_LO;
    re_MAP_IP_HI_t MAP_IP_HI;
    re_MAP_IP_CFG_t MAP_IP_CFG;
    re_MAP_PROT_t MAP_PROT;
    re_MAP_L4_SRC_t MAP_L4_SRC;
    re_MAP_L4_DST_t MAP_L4_DST;
    re_MAP_EXP_TC_t MAP_EXP_TC;
    re_MAP_DSCP_TC_t MAP_DSCP_TC;
    re_MAP_VPRI_TC_t MAP_VPRI_TC;
    re_MAP_VPRI_t MAP_VPRI;
    re_MAP_PROFILE_KEY0_t MAP_PROFILE_KEY0;
    re_MAP_PROFILE_KEY_INVERT0_t MAP_PROFILE_KEY_INVERT0;
    re_MAP_PROFILE_KEY1_t MAP_PROFILE_KEY1;
    re_MAP_PROFILE_KEY_INVERT1_t MAP_PROFILE_KEY_INVERT1;
    re_MAP_PROFILE_ACTION_t MAP_PROFILE_ACTION;
    re_MAP_DOMAIN_POL_CFG_t MAP_DOMAIN_POL_CFG;
    re_MAP_REWRITE_t MAP_REWRITE;
} mby_ppe_mapper_map_hc_re_t;

typedef logic handcode_rvalid_MAP_PORT_CFG_t;

typedef logic handcode_rvalid_MAP_PORT_DEFAULT_t;

typedef logic handcode_rvalid_MAP_DOMAIN_TCAM_t;

typedef logic handcode_rvalid_MAP_DOMAIN_ACTION0_t;

typedef logic handcode_rvalid_MAP_DOMAIN_ACTION1_t;

typedef logic handcode_rvalid_MAP_DOMAIN_PROFILE_t;

typedef logic handcode_rvalid_MAP_PORT_t;

typedef logic handcode_rvalid_MAP_MAC_t;

typedef logic handcode_rvalid_MAP_IP_LO_t;

typedef logic handcode_rvalid_MAP_IP_HI_t;

typedef logic handcode_rvalid_MAP_IP_CFG_t;

typedef logic handcode_rvalid_MAP_PROT_t;

typedef logic handcode_rvalid_MAP_L4_SRC_t;

typedef logic handcode_rvalid_MAP_L4_DST_t;

typedef logic handcode_rvalid_MAP_EXP_TC_t;

typedef logic handcode_rvalid_MAP_DSCP_TC_t;

typedef logic handcode_rvalid_MAP_VPRI_TC_t;

typedef logic handcode_rvalid_MAP_VPRI_t;

typedef logic handcode_rvalid_MAP_PROFILE_KEY0_t;

typedef logic handcode_rvalid_MAP_PROFILE_KEY_INVERT0_t;

typedef logic handcode_rvalid_MAP_PROFILE_KEY1_t;

typedef logic handcode_rvalid_MAP_PROFILE_KEY_INVERT1_t;

typedef logic handcode_rvalid_MAP_PROFILE_ACTION_t;

typedef logic handcode_rvalid_MAP_DOMAIN_POL_CFG_t;

typedef logic handcode_rvalid_MAP_REWRITE_t;

typedef struct packed {
    handcode_rvalid_MAP_PORT_CFG_t MAP_PORT_CFG;
    handcode_rvalid_MAP_PORT_DEFAULT_t MAP_PORT_DEFAULT;
    handcode_rvalid_MAP_DOMAIN_TCAM_t MAP_DOMAIN_TCAM;
    handcode_rvalid_MAP_DOMAIN_ACTION0_t MAP_DOMAIN_ACTION0;
    handcode_rvalid_MAP_DOMAIN_ACTION1_t MAP_DOMAIN_ACTION1;
    handcode_rvalid_MAP_DOMAIN_PROFILE_t MAP_DOMAIN_PROFILE;
    handcode_rvalid_MAP_PORT_t MAP_PORT;
    handcode_rvalid_MAP_MAC_t MAP_MAC;
    handcode_rvalid_MAP_IP_LO_t MAP_IP_LO;
    handcode_rvalid_MAP_IP_HI_t MAP_IP_HI;
    handcode_rvalid_MAP_IP_CFG_t MAP_IP_CFG;
    handcode_rvalid_MAP_PROT_t MAP_PROT;
    handcode_rvalid_MAP_L4_SRC_t MAP_L4_SRC;
    handcode_rvalid_MAP_L4_DST_t MAP_L4_DST;
    handcode_rvalid_MAP_EXP_TC_t MAP_EXP_TC;
    handcode_rvalid_MAP_DSCP_TC_t MAP_DSCP_TC;
    handcode_rvalid_MAP_VPRI_TC_t MAP_VPRI_TC;
    handcode_rvalid_MAP_VPRI_t MAP_VPRI;
    handcode_rvalid_MAP_PROFILE_KEY0_t MAP_PROFILE_KEY0;
    handcode_rvalid_MAP_PROFILE_KEY_INVERT0_t MAP_PROFILE_KEY_INVERT0;
    handcode_rvalid_MAP_PROFILE_KEY1_t MAP_PROFILE_KEY1;
    handcode_rvalid_MAP_PROFILE_KEY_INVERT1_t MAP_PROFILE_KEY_INVERT1;
    handcode_rvalid_MAP_PROFILE_ACTION_t MAP_PROFILE_ACTION;
    handcode_rvalid_MAP_DOMAIN_POL_CFG_t MAP_DOMAIN_POL_CFG;
    handcode_rvalid_MAP_REWRITE_t MAP_REWRITE;
} mby_ppe_mapper_map_hc_rvalid_t;

typedef logic handcode_wvalid_MAP_PORT_CFG_t;

typedef logic handcode_wvalid_MAP_PORT_DEFAULT_t;

typedef logic handcode_wvalid_MAP_DOMAIN_TCAM_t;

typedef logic handcode_wvalid_MAP_DOMAIN_ACTION0_t;

typedef logic handcode_wvalid_MAP_DOMAIN_ACTION1_t;

typedef logic handcode_wvalid_MAP_DOMAIN_PROFILE_t;

typedef logic handcode_wvalid_MAP_PORT_t;

typedef logic handcode_wvalid_MAP_MAC_t;

typedef logic handcode_wvalid_MAP_IP_LO_t;

typedef logic handcode_wvalid_MAP_IP_HI_t;

typedef logic handcode_wvalid_MAP_IP_CFG_t;

typedef logic handcode_wvalid_MAP_PROT_t;

typedef logic handcode_wvalid_MAP_L4_SRC_t;

typedef logic handcode_wvalid_MAP_L4_DST_t;

typedef logic handcode_wvalid_MAP_EXP_TC_t;

typedef logic handcode_wvalid_MAP_DSCP_TC_t;

typedef logic handcode_wvalid_MAP_VPRI_TC_t;

typedef logic handcode_wvalid_MAP_VPRI_t;

typedef logic handcode_wvalid_MAP_PROFILE_KEY0_t;

typedef logic handcode_wvalid_MAP_PROFILE_KEY_INVERT0_t;

typedef logic handcode_wvalid_MAP_PROFILE_KEY1_t;

typedef logic handcode_wvalid_MAP_PROFILE_KEY_INVERT1_t;

typedef logic handcode_wvalid_MAP_PROFILE_ACTION_t;

typedef logic handcode_wvalid_MAP_DOMAIN_POL_CFG_t;

typedef logic handcode_wvalid_MAP_REWRITE_t;

typedef struct packed {
    handcode_wvalid_MAP_PORT_CFG_t MAP_PORT_CFG;
    handcode_wvalid_MAP_PORT_DEFAULT_t MAP_PORT_DEFAULT;
    handcode_wvalid_MAP_DOMAIN_TCAM_t MAP_DOMAIN_TCAM;
    handcode_wvalid_MAP_DOMAIN_ACTION0_t MAP_DOMAIN_ACTION0;
    handcode_wvalid_MAP_DOMAIN_ACTION1_t MAP_DOMAIN_ACTION1;
    handcode_wvalid_MAP_DOMAIN_PROFILE_t MAP_DOMAIN_PROFILE;
    handcode_wvalid_MAP_PORT_t MAP_PORT;
    handcode_wvalid_MAP_MAC_t MAP_MAC;
    handcode_wvalid_MAP_IP_LO_t MAP_IP_LO;
    handcode_wvalid_MAP_IP_HI_t MAP_IP_HI;
    handcode_wvalid_MAP_IP_CFG_t MAP_IP_CFG;
    handcode_wvalid_MAP_PROT_t MAP_PROT;
    handcode_wvalid_MAP_L4_SRC_t MAP_L4_SRC;
    handcode_wvalid_MAP_L4_DST_t MAP_L4_DST;
    handcode_wvalid_MAP_EXP_TC_t MAP_EXP_TC;
    handcode_wvalid_MAP_DSCP_TC_t MAP_DSCP_TC;
    handcode_wvalid_MAP_VPRI_TC_t MAP_VPRI_TC;
    handcode_wvalid_MAP_VPRI_t MAP_VPRI;
    handcode_wvalid_MAP_PROFILE_KEY0_t MAP_PROFILE_KEY0;
    handcode_wvalid_MAP_PROFILE_KEY_INVERT0_t MAP_PROFILE_KEY_INVERT0;
    handcode_wvalid_MAP_PROFILE_KEY1_t MAP_PROFILE_KEY1;
    handcode_wvalid_MAP_PROFILE_KEY_INVERT1_t MAP_PROFILE_KEY_INVERT1;
    handcode_wvalid_MAP_PROFILE_ACTION_t MAP_PROFILE_ACTION;
    handcode_wvalid_MAP_DOMAIN_POL_CFG_t MAP_DOMAIN_POL_CFG;
    handcode_wvalid_MAP_REWRITE_t MAP_REWRITE;
} mby_ppe_mapper_map_hc_wvalid_t;

typedef logic handcode_error_MAP_PORT_CFG_t;

typedef logic handcode_error_MAP_PORT_DEFAULT_t;

typedef logic handcode_error_MAP_DOMAIN_TCAM_t;

typedef logic handcode_error_MAP_DOMAIN_ACTION0_t;

typedef logic handcode_error_MAP_DOMAIN_ACTION1_t;

typedef logic handcode_error_MAP_DOMAIN_PROFILE_t;

typedef logic handcode_error_MAP_PORT_t;

typedef logic handcode_error_MAP_MAC_t;

typedef logic handcode_error_MAP_IP_LO_t;

typedef logic handcode_error_MAP_IP_HI_t;

typedef logic handcode_error_MAP_IP_CFG_t;

typedef logic handcode_error_MAP_PROT_t;

typedef logic handcode_error_MAP_L4_SRC_t;

typedef logic handcode_error_MAP_L4_DST_t;

typedef logic handcode_error_MAP_EXP_TC_t;

typedef logic handcode_error_MAP_DSCP_TC_t;

typedef logic handcode_error_MAP_VPRI_TC_t;

typedef logic handcode_error_MAP_VPRI_t;

typedef logic handcode_error_MAP_PROFILE_KEY0_t;

typedef logic handcode_error_MAP_PROFILE_KEY_INVERT0_t;

typedef logic handcode_error_MAP_PROFILE_KEY1_t;

typedef logic handcode_error_MAP_PROFILE_KEY_INVERT1_t;

typedef logic handcode_error_MAP_PROFILE_ACTION_t;

typedef logic handcode_error_MAP_DOMAIN_POL_CFG_t;

typedef logic handcode_error_MAP_REWRITE_t;

typedef struct packed {
    handcode_error_MAP_PORT_CFG_t MAP_PORT_CFG;
    handcode_error_MAP_PORT_DEFAULT_t MAP_PORT_DEFAULT;
    handcode_error_MAP_DOMAIN_TCAM_t MAP_DOMAIN_TCAM;
    handcode_error_MAP_DOMAIN_ACTION0_t MAP_DOMAIN_ACTION0;
    handcode_error_MAP_DOMAIN_ACTION1_t MAP_DOMAIN_ACTION1;
    handcode_error_MAP_DOMAIN_PROFILE_t MAP_DOMAIN_PROFILE;
    handcode_error_MAP_PORT_t MAP_PORT;
    handcode_error_MAP_MAC_t MAP_MAC;
    handcode_error_MAP_IP_LO_t MAP_IP_LO;
    handcode_error_MAP_IP_HI_t MAP_IP_HI;
    handcode_error_MAP_IP_CFG_t MAP_IP_CFG;
    handcode_error_MAP_PROT_t MAP_PROT;
    handcode_error_MAP_L4_SRC_t MAP_L4_SRC;
    handcode_error_MAP_L4_DST_t MAP_L4_DST;
    handcode_error_MAP_EXP_TC_t MAP_EXP_TC;
    handcode_error_MAP_DSCP_TC_t MAP_DSCP_TC;
    handcode_error_MAP_VPRI_TC_t MAP_VPRI_TC;
    handcode_error_MAP_VPRI_t MAP_VPRI;
    handcode_error_MAP_PROFILE_KEY0_t MAP_PROFILE_KEY0;
    handcode_error_MAP_PROFILE_KEY_INVERT0_t MAP_PROFILE_KEY_INVERT0;
    handcode_error_MAP_PROFILE_KEY1_t MAP_PROFILE_KEY1;
    handcode_error_MAP_PROFILE_KEY_INVERT1_t MAP_PROFILE_KEY_INVERT1;
    handcode_error_MAP_PROFILE_ACTION_t MAP_PROFILE_ACTION;
    handcode_error_MAP_DOMAIN_POL_CFG_t MAP_DOMAIN_POL_CFG;
    handcode_error_MAP_REWRITE_t MAP_REWRITE;
} mby_ppe_mapper_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    MAP_PORT_CFG_t MAP_PORT_CFG;
    MAP_PORT_DEFAULT_t MAP_PORT_DEFAULT;
    MAP_DOMAIN_TCAM_t MAP_DOMAIN_TCAM;
    MAP_DOMAIN_ACTION0_t MAP_DOMAIN_ACTION0;
    MAP_DOMAIN_ACTION1_t MAP_DOMAIN_ACTION1;
    MAP_DOMAIN_PROFILE_t MAP_DOMAIN_PROFILE;
    MAP_PORT_t MAP_PORT;
    MAP_MAC_t MAP_MAC;
    MAP_IP_LO_t MAP_IP_LO;
    MAP_IP_HI_t MAP_IP_HI;
    MAP_IP_CFG_t MAP_IP_CFG;
    MAP_PROT_t MAP_PROT;
    MAP_L4_SRC_t MAP_L4_SRC;
    MAP_L4_DST_t MAP_L4_DST;
    MAP_EXP_TC_t MAP_EXP_TC;
    MAP_DSCP_TC_t MAP_DSCP_TC;
    MAP_VPRI_TC_t MAP_VPRI_TC;
    MAP_VPRI_t MAP_VPRI;
    MAP_PROFILE_KEY0_t MAP_PROFILE_KEY0;
    MAP_PROFILE_KEY_INVERT0_t MAP_PROFILE_KEY_INVERT0;
    MAP_PROFILE_KEY1_t MAP_PROFILE_KEY1;
    MAP_PROFILE_KEY_INVERT1_t MAP_PROFILE_KEY_INVERT1;
    MAP_PROFILE_ACTION_t MAP_PROFILE_ACTION;
    MAP_DOMAIN_POL_CFG_t MAP_DOMAIN_POL_CFG;
    MAP_REWRITE_t MAP_REWRITE;
} mby_ppe_mapper_map_hc_reg_read_t;

typedef struct packed {
    MAP_PORT_CFG_t MAP_PORT_CFG;
    MAP_PORT_DEFAULT_t MAP_PORT_DEFAULT;
    MAP_DOMAIN_TCAM_t MAP_DOMAIN_TCAM;
    MAP_DOMAIN_ACTION0_t MAP_DOMAIN_ACTION0;
    MAP_DOMAIN_ACTION1_t MAP_DOMAIN_ACTION1;
    MAP_DOMAIN_PROFILE_t MAP_DOMAIN_PROFILE;
    MAP_PORT_t MAP_PORT;
    MAP_MAC_t MAP_MAC;
    MAP_IP_LO_t MAP_IP_LO;
    MAP_IP_HI_t MAP_IP_HI;
    MAP_IP_CFG_t MAP_IP_CFG;
    MAP_PROT_t MAP_PROT;
    MAP_L4_SRC_t MAP_L4_SRC;
    MAP_L4_DST_t MAP_L4_DST;
    MAP_EXP_TC_t MAP_EXP_TC;
    MAP_DSCP_TC_t MAP_DSCP_TC;
    MAP_VPRI_TC_t MAP_VPRI_TC;
    MAP_VPRI_t MAP_VPRI;
    MAP_PROFILE_KEY0_t MAP_PROFILE_KEY0;
    MAP_PROFILE_KEY_INVERT0_t MAP_PROFILE_KEY_INVERT0;
    MAP_PROFILE_KEY1_t MAP_PROFILE_KEY1;
    MAP_PROFILE_KEY_INVERT1_t MAP_PROFILE_KEY_INVERT1;
    MAP_PROFILE_ACTION_t MAP_PROFILE_ACTION;
    MAP_DOMAIN_POL_CFG_t MAP_DOMAIN_POL_CFG;
    MAP_REWRITE_t MAP_REWRITE;
} mby_ppe_mapper_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_mapper_map_pkg

`endif // MBY_PPE_MAPPER_MAP_PKG_VH
