// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

// -----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Raghu P Gudla
// Created On   :  09/22/2018
// Description  :  Configuration file for HVL hierarchy
// -----------------------------------------------------------------------------
  
config `HVL_TOP_CFG;
    design `HVL_TOP_LIB.`HVL_TOP;
endconfig
/*
 *  ----------------
 *    End of file
 *  ----------------
*/
