// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

    
    `include "fc_lite_config_include.svh"

// Example reference code. To be cleaned up
//    `ifndef PMU_RTL_ENABLE
//      instance `PMU_WRAPPER use `RTL_STUB_LIB.;
//    `else
//      instance `PMU_WRAPPER use pmu_rtl_lib.;
//    `end      
