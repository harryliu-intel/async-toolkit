magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect 3 73 11 74
rect 3 65 11 70
rect 3 57 11 62
rect 3 49 11 54
rect 3 41 11 46
rect 3 37 11 38
<< pdiffusion >>
rect 27 83 35 84
rect 27 79 35 80
rect 27 70 35 71
rect 27 66 35 67
rect 27 57 35 58
rect 27 53 35 54
rect 27 44 35 45
rect 27 40 35 41
rect 27 31 35 32
rect 27 27 35 28
<< ntransistor >>
rect 3 70 11 73
rect 3 62 11 65
rect 3 54 11 57
rect 3 46 11 49
rect 3 38 11 41
<< ptransistor >>
rect 27 80 35 83
rect 27 67 35 70
rect 27 54 35 57
rect 27 41 35 44
rect 27 28 35 31
<< polysilicon >>
rect 13 80 27 83
rect 35 80 39 83
rect 13 73 16 80
rect -1 70 3 73
rect 11 70 16 73
rect 22 67 27 70
rect 35 67 39 70
rect 22 65 25 67
rect -1 62 3 65
rect 11 62 25 65
rect -1 54 3 57
rect 11 54 27 57
rect 35 54 39 57
rect -1 46 3 49
rect 11 46 25 49
rect 22 44 25 46
rect 22 41 27 44
rect 35 41 39 44
rect -1 38 3 41
rect 11 38 16 41
rect 13 31 16 38
rect 13 28 27 31
rect 35 28 39 31
<< ndcontact >>
rect 3 74 11 82
rect 3 29 11 37
<< pdcontact >>
rect 27 84 35 92
rect 27 71 35 79
rect 27 58 35 66
rect 27 45 35 53
rect 27 32 35 40
rect 27 19 35 27
<< metal1 >>
rect 15 84 35 92
rect 15 82 23 84
rect 3 74 23 82
rect 15 66 23 74
rect 27 71 35 79
rect 15 58 35 66
rect 15 40 23 58
rect 27 45 35 53
rect 3 29 11 37
rect 15 32 35 40
rect 27 19 35 27
<< labels >>
rlabel metal1 31 36 31 36 1 x
rlabel metal1 31 49 31 49 5 Vdd!
rlabel metal1 31 23 31 23 1 Vdd!
rlabel polysilicon 36 42 36 42 1 b
rlabel polysilicon 36 29 36 29 1 a
rlabel metal1 31 62 31 62 5 x
rlabel polysilicon 36 55 36 55 1 c
rlabel metal1 31 75 31 75 1 Vdd!
rlabel polysilicon 36 68 36 68 1 d
rlabel metal1 31 88 31 88 1 x
rlabel polysilicon 36 81 36 81 1 e
rlabel metal1 7 33 7 33 1 GND!
rlabel polysilicon 2 39 2 39 3 a
rlabel polysilicon 2 47 2 47 3 b
rlabel polysilicon 2 55 2 55 3 c
rlabel polysilicon 2 63 2 63 3 d
rlabel metal1 7 78 7 78 1 x
rlabel polysilicon 2 71 2 71 3 e
rlabel space -2 29 3 82 7 ^n
rlabel space 35 19 40 92 3 ^p
<< end >>
