// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

// -------------------------------------------------------------------------
// This file binds the formal assertions to the DUT 

   bind mby_top mby_checker mby_checker0 (.*);
