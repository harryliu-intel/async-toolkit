    
    `include "fc_lite_config_include.svh"

// Example reference code. To be cleaned up
//    `ifndef PMU_RTL_ENABLE
//      instance `PMU_WRAPPER use `RTL_STUB_LIB.;
//    `else
//      instance `PMU_WRAPPER use pmu_rtl_lib.;
//    `end      
