magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -220 -716 -214 -715
rect -220 -722 -214 -718
rect -220 -728 -214 -724
rect -220 -734 -214 -730
rect -220 -740 -214 -736
rect -220 -746 -214 -742
rect -220 -749 -214 -748
rect -220 -753 -218 -749
rect -220 -754 -214 -753
rect -220 -760 -214 -756
rect -220 -766 -214 -762
rect -220 -772 -214 -768
rect -220 -778 -214 -774
rect -220 -784 -214 -780
rect -220 -787 -214 -786
<< pdiffusion >>
rect -199 -706 -189 -705
rect -199 -709 -189 -708
rect -191 -713 -189 -709
rect -199 -714 -189 -713
rect -199 -717 -189 -716
rect -199 -721 -193 -717
rect -199 -722 -189 -721
rect -199 -725 -189 -724
rect -191 -729 -189 -725
rect -199 -730 -189 -729
rect -199 -733 -189 -732
rect -199 -737 -193 -733
rect -199 -738 -189 -737
rect -199 -741 -189 -740
rect -191 -745 -189 -741
rect -199 -746 -189 -745
rect -199 -749 -189 -748
rect -199 -753 -193 -749
rect -199 -754 -189 -753
rect -199 -757 -189 -756
rect -191 -761 -189 -757
rect -199 -762 -189 -761
rect -199 -765 -189 -764
rect -199 -769 -193 -765
rect -199 -770 -189 -769
rect -199 -773 -189 -772
rect -191 -777 -189 -773
rect -199 -778 -189 -777
rect -199 -781 -189 -780
rect -199 -785 -193 -781
rect -199 -786 -189 -785
rect -199 -789 -189 -788
rect -191 -793 -189 -789
rect -199 -794 -189 -793
rect -199 -797 -189 -796
<< ntransistor >>
rect -220 -718 -214 -716
rect -220 -724 -214 -722
rect -220 -730 -214 -728
rect -220 -736 -214 -734
rect -220 -742 -214 -740
rect -220 -748 -214 -746
rect -220 -756 -214 -754
rect -220 -762 -214 -760
rect -220 -768 -214 -766
rect -220 -774 -214 -772
rect -220 -780 -214 -778
rect -220 -786 -214 -784
<< ptransistor >>
rect -199 -708 -189 -706
rect -199 -716 -189 -714
rect -199 -724 -189 -722
rect -199 -732 -189 -730
rect -199 -740 -189 -738
rect -199 -748 -189 -746
rect -199 -756 -189 -754
rect -199 -764 -189 -762
rect -199 -772 -189 -770
rect -199 -780 -189 -778
rect -199 -788 -189 -786
rect -199 -796 -189 -794
<< polysilicon >>
rect -203 -708 -199 -706
rect -189 -708 -186 -706
rect -203 -714 -201 -708
rect -203 -716 -199 -714
rect -189 -716 -186 -714
rect -223 -718 -220 -716
rect -214 -718 -201 -716
rect -223 -724 -220 -722
rect -214 -724 -199 -722
rect -189 -724 -186 -722
rect -223 -730 -220 -728
rect -214 -730 -211 -728
rect -203 -732 -199 -730
rect -189 -732 -186 -730
rect -203 -734 -201 -732
rect -223 -736 -220 -734
rect -214 -736 -201 -734
rect -203 -738 -201 -736
rect -203 -740 -199 -738
rect -189 -740 -186 -738
rect -223 -742 -220 -740
rect -214 -742 -206 -740
rect -208 -746 -206 -742
rect -223 -748 -220 -746
rect -214 -748 -211 -746
rect -208 -748 -199 -746
rect -189 -748 -186 -746
rect -223 -756 -220 -754
rect -214 -756 -211 -754
rect -208 -756 -199 -754
rect -189 -756 -186 -754
rect -208 -760 -206 -756
rect -223 -762 -220 -760
rect -214 -762 -206 -760
rect -203 -764 -199 -762
rect -189 -764 -186 -762
rect -203 -766 -201 -764
rect -223 -768 -220 -766
rect -214 -768 -201 -766
rect -203 -770 -201 -768
rect -203 -772 -199 -770
rect -189 -772 -186 -770
rect -223 -774 -220 -772
rect -214 -774 -211 -772
rect -223 -780 -220 -778
rect -214 -780 -199 -778
rect -189 -780 -186 -778
rect -223 -786 -220 -784
rect -214 -786 -201 -784
rect -203 -788 -199 -786
rect -189 -788 -186 -786
rect -203 -794 -201 -788
rect -203 -796 -199 -794
rect -189 -796 -186 -794
<< ndcontact >>
rect -220 -715 -214 -711
rect -218 -753 -214 -749
rect -220 -791 -214 -787
<< pdcontact >>
rect -199 -705 -189 -701
rect -199 -713 -191 -709
rect -193 -721 -189 -717
rect -199 -729 -191 -725
rect -193 -737 -189 -733
rect -199 -745 -191 -741
rect -193 -753 -189 -749
rect -199 -761 -191 -757
rect -193 -769 -189 -765
rect -199 -777 -191 -773
rect -193 -785 -189 -781
rect -199 -793 -191 -789
rect -199 -801 -189 -797
<< metal1 >>
rect -199 -705 -189 -701
rect -220 -715 -214 -711
rect -199 -713 -191 -709
rect -199 -725 -196 -713
rect -193 -721 -189 -717
rect -199 -729 -191 -725
rect -199 -741 -196 -729
rect -193 -737 -189 -733
rect -199 -745 -191 -741
rect -199 -749 -196 -745
rect -218 -753 -196 -749
rect -193 -753 -189 -749
rect -199 -757 -196 -753
rect -199 -761 -191 -757
rect -199 -773 -196 -761
rect -193 -769 -189 -765
rect -199 -777 -191 -773
rect -220 -791 -214 -787
rect -199 -789 -196 -777
rect -193 -785 -189 -781
rect -199 -793 -191 -789
rect -199 -801 -189 -797
<< labels >>
rlabel space -192 -802 -186 -700 3 ^p
rlabel polysilicon -188 -795 -188 -795 3 a
rlabel polysilicon -188 -787 -188 -787 3 a
rlabel polysilicon -188 -779 -188 -779 3 b
rlabel polysilicon -188 -771 -188 -771 3 d
rlabel polysilicon -188 -763 -188 -763 3 d
rlabel polysilicon -188 -755 -188 -755 3 e
rlabel polysilicon -188 -747 -188 -747 3 b
rlabel polysilicon -188 -739 -188 -739 3 c
rlabel polysilicon -188 -731 -188 -731 3 c
rlabel polysilicon -188 -723 -188 -723 3 e
rlabel polysilicon -188 -715 -188 -715 3 f
rlabel polysilicon -188 -707 -188 -707 3 f
rlabel polysilicon -221 -785 -221 -785 3 a
rlabel polysilicon -221 -779 -221 -779 3 b
rlabel polysilicon -221 -773 -221 -773 3 c
rlabel polysilicon -221 -767 -221 -767 3 d
rlabel polysilicon -221 -761 -221 -761 3 e
rlabel polysilicon -221 -755 -221 -755 3 f
rlabel polysilicon -221 -747 -221 -747 3 a
rlabel polysilicon -221 -741 -221 -741 3 b
rlabel polysilicon -221 -735 -221 -735 3 c
rlabel polysilicon -221 -729 -221 -729 3 d
rlabel polysilicon -221 -723 -221 -723 3 e
rlabel polysilicon -221 -717 -221 -717 3 f
rlabel space -223 -793 -217 -710 7 ^n
rlabel pdcontact -197 -791 -197 -791 1 x
rlabel pdcontact -197 -775 -197 -775 1 x
rlabel pdcontact -197 -759 -197 -759 1 x
rlabel pdcontact -197 -743 -197 -743 1 x
rlabel pdcontact -197 -727 -197 -727 1 x
rlabel pdcontact -197 -711 -197 -711 1 x
rlabel pdcontact -191 -767 -191 -767 1 Vdd!
rlabel pdcontact -191 -783 -191 -783 1 Vdd!
rlabel pdcontact -191 -799 -191 -799 1 Vdd!
rlabel pdcontact -191 -735 -191 -735 1 Vdd!
rlabel pdcontact -191 -751 -191 -751 1 Vdd!
rlabel pdcontact -191 -719 -191 -719 1 Vdd!
rlabel pdcontact -191 -703 -191 -703 1 Vdd!
rlabel ndcontact -216 -789 -216 -789 1 GND!
rlabel ndcontact -216 -713 -216 -713 5 GND!
rlabel ndcontact -216 -751 -216 -751 1 x
<< end >>
