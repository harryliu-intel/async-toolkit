magic
tech scmos
timestamp 969760391
<< ndiffusion >>
rect 15 150 23 151
rect 45 150 53 151
rect 15 142 23 147
rect -7 129 1 134
rect 15 138 23 139
rect 15 129 23 130
rect 45 142 53 147
rect 45 138 53 139
rect 45 129 53 130
rect -7 118 1 126
rect 15 121 23 126
rect 45 121 53 126
rect 15 117 23 118
rect 15 108 23 109
rect 45 117 53 118
rect 45 108 53 109
rect 15 100 23 105
rect 45 100 53 105
rect -15 94 -7 95
rect -15 90 -7 91
rect 15 92 23 97
rect 45 92 53 97
rect 15 88 23 89
rect 15 79 23 80
rect 15 71 23 76
rect 45 88 53 89
rect 45 79 53 80
rect 45 71 53 76
rect 15 63 23 68
rect 45 63 53 68
rect 15 59 23 60
rect 15 50 23 51
rect 45 59 53 60
rect 45 50 53 51
rect -7 42 1 50
rect 15 42 23 47
rect 45 42 53 47
rect -7 34 1 39
rect 15 38 23 39
rect 15 29 23 30
rect 15 21 23 26
rect 45 38 53 39
rect 45 29 53 30
rect 45 21 53 26
rect 15 17 23 18
rect 45 17 53 18
<< pdiffusion >>
rect 69 150 77 151
rect 98 150 110 151
rect 124 150 136 151
rect 69 142 77 147
rect 98 142 110 147
rect 124 146 136 147
rect 69 138 77 139
rect 69 129 77 130
rect 69 121 77 126
rect 98 138 110 139
rect 98 129 110 130
rect 132 141 136 146
rect 98 121 110 126
rect 69 117 77 118
rect 98 117 110 118
rect 69 100 77 101
rect 123 107 139 108
rect 98 100 110 101
rect 123 103 139 104
rect 123 98 128 103
rect 69 92 77 97
rect 69 88 77 89
rect 69 79 77 80
rect 98 92 110 97
rect 136 98 139 103
rect 98 88 110 89
rect 98 79 110 80
rect 69 71 77 76
rect 98 71 110 76
rect 132 72 136 77
rect 124 71 136 72
rect 69 67 77 68
rect 69 50 77 51
rect 98 67 110 68
rect 124 67 136 68
rect 98 50 110 51
rect 69 42 77 47
rect 69 38 77 39
rect 69 29 77 30
rect 98 42 110 47
rect 98 38 110 39
rect 98 29 110 30
rect 69 21 77 26
rect 98 21 110 26
rect 132 22 136 27
rect 124 21 136 22
rect 69 17 77 18
rect 98 17 110 18
rect 124 17 136 18
<< ntransistor >>
rect 15 147 23 150
rect 45 147 53 150
rect 15 139 23 142
rect 45 139 53 142
rect -7 126 1 129
rect 15 126 23 129
rect 45 126 53 129
rect 15 118 23 121
rect 45 118 53 121
rect 15 105 23 108
rect 45 105 53 108
rect 15 97 23 100
rect 45 97 53 100
rect -15 91 -7 94
rect 15 89 23 92
rect 45 89 53 92
rect 15 76 23 79
rect 45 76 53 79
rect 15 68 23 71
rect 45 68 53 71
rect 15 60 23 63
rect 45 60 53 63
rect 15 47 23 50
rect 45 47 53 50
rect -7 39 1 42
rect 15 39 23 42
rect 45 39 53 42
rect 15 26 23 29
rect 45 26 53 29
rect 15 18 23 21
rect 45 18 53 21
<< ptransistor >>
rect 69 147 77 150
rect 98 147 110 150
rect 124 147 136 150
rect 69 139 77 142
rect 98 139 110 142
rect 69 126 77 129
rect 98 126 110 129
rect 69 118 77 121
rect 98 118 110 121
rect 69 97 77 100
rect 123 104 139 107
rect 98 97 110 100
rect 69 89 77 92
rect 98 89 110 92
rect 69 76 77 79
rect 98 76 110 79
rect 69 68 77 71
rect 98 68 110 71
rect 124 68 136 71
rect 69 47 77 50
rect 98 47 110 50
rect 69 39 77 42
rect 98 39 110 42
rect 69 26 77 29
rect 98 26 110 29
rect 69 18 77 21
rect 98 18 110 21
rect 124 18 136 21
<< polysilicon >>
rect 11 147 15 150
rect 23 147 45 150
rect 53 147 69 150
rect 77 147 98 150
rect 110 147 114 150
rect 120 147 124 150
rect 136 147 141 150
rect 11 139 15 142
rect 23 139 28 142
rect 11 134 13 139
rect 10 129 13 134
rect 33 129 36 147
rect 41 139 45 142
rect 53 139 69 142
rect 77 139 89 142
rect 94 139 98 142
rect 110 139 114 142
rect -9 126 -7 129
rect 1 126 5 129
rect 10 126 15 129
rect 23 126 28 129
rect 33 126 45 129
rect 53 126 69 129
rect 77 126 81 129
rect 86 121 89 139
rect 112 134 114 139
rect 138 134 141 147
rect 112 129 115 134
rect 94 126 98 129
rect 110 126 115 129
rect 136 131 141 134
rect 11 118 15 121
rect 23 118 45 121
rect 53 118 69 121
rect 77 118 98 121
rect 110 118 114 121
rect 11 105 15 108
rect 23 105 45 108
rect 53 105 57 108
rect 11 97 15 100
rect 23 97 45 100
rect 53 97 69 100
rect 77 97 84 100
rect 119 104 123 107
rect 139 104 143 107
rect 92 97 98 100
rect 110 97 114 100
rect -19 91 -15 94
rect -7 91 -3 94
rect 10 89 15 92
rect 23 89 28 92
rect 33 89 45 92
rect 53 89 69 92
rect 77 89 81 92
rect 10 84 13 89
rect 11 79 13 84
rect 11 76 15 79
rect 23 76 28 79
rect 33 71 36 89
rect 86 79 89 97
rect 94 89 98 92
rect 110 89 115 92
rect 112 84 115 89
rect 136 84 141 87
rect 112 79 114 84
rect 41 76 45 79
rect 53 76 69 79
rect 77 76 89 79
rect 94 76 98 79
rect 110 76 114 79
rect 138 71 141 84
rect -9 68 15 71
rect 23 68 45 71
rect 53 68 69 71
rect 77 68 98 71
rect 110 68 114 71
rect 120 68 124 71
rect 136 68 141 71
rect 11 60 15 63
rect 23 60 45 63
rect 53 60 57 63
rect 11 47 15 50
rect 23 47 45 50
rect 53 47 69 50
rect 77 47 98 50
rect 110 47 114 50
rect -9 39 -7 42
rect 1 39 5 42
rect 10 39 15 42
rect 23 39 28 42
rect 33 39 45 42
rect 53 39 69 42
rect 77 39 81 42
rect 10 34 13 39
rect 11 29 13 34
rect 11 26 15 29
rect 23 26 28 29
rect 33 21 36 39
rect 86 29 89 47
rect 94 39 98 42
rect 110 39 115 42
rect 112 34 115 39
rect 136 34 141 37
rect 112 29 114 34
rect 41 26 45 29
rect 53 26 69 29
rect 77 26 89 29
rect 94 26 98 29
rect 110 26 114 29
rect 138 21 141 34
rect 11 18 15 21
rect 23 18 45 21
rect 53 18 69 21
rect 77 18 98 21
rect 110 18 114 21
rect 120 18 124 21
rect 136 18 141 21
<< ndcontact >>
rect 15 151 23 159
rect 45 151 53 159
rect -7 134 1 142
rect 15 130 23 138
rect 45 130 53 138
rect -7 110 1 118
rect 15 109 23 117
rect 45 109 53 117
rect -15 95 -7 103
rect -15 82 -7 90
rect 15 80 23 88
rect 45 80 53 88
rect -7 50 1 58
rect 15 51 23 59
rect 45 51 53 59
rect -7 26 1 34
rect 15 30 23 38
rect 45 30 53 38
rect 15 9 23 17
rect 45 9 53 17
<< pdcontact >>
rect 69 151 77 159
rect 98 151 110 159
rect 124 151 136 159
rect 69 130 77 138
rect 98 130 110 138
rect 124 138 132 146
rect 69 101 77 117
rect 98 101 110 117
rect 123 108 139 116
rect 69 80 77 88
rect 128 95 136 103
rect 98 80 110 88
rect 124 72 132 80
rect 69 51 77 67
rect 98 51 110 67
rect 124 59 136 67
rect 69 30 77 38
rect 98 30 110 38
rect 124 22 132 30
rect 69 9 77 17
rect 98 9 110 17
rect 124 9 136 17
<< polycontact >>
rect 3 134 11 142
rect -17 122 -9 130
rect 114 134 122 142
rect 128 126 136 134
rect 84 97 92 105
rect -3 89 5 97
rect 3 76 11 84
rect -17 68 -9 76
rect 128 84 136 92
rect 114 76 122 84
rect -17 38 -9 46
rect 3 26 11 34
rect 128 34 136 42
rect 114 26 122 34
<< metal1 >>
rect 15 151 53 159
rect 69 151 136 159
rect 6 146 128 147
rect 6 142 132 146
rect -7 134 11 142
rect 114 138 132 142
rect 15 130 110 138
rect 114 134 122 138
rect 128 130 136 134
rect -17 122 23 130
rect -7 117 1 118
rect -15 110 53 117
rect -15 95 -7 110
rect 15 109 53 110
rect 58 97 64 130
rect 106 126 136 130
rect 69 116 110 117
rect 69 109 139 116
rect 69 101 77 109
rect 84 97 92 105
rect 98 101 110 109
rect 123 108 139 109
rect -3 95 5 97
rect -15 84 -7 90
rect -3 89 23 95
rect 58 92 89 97
rect 128 92 136 103
rect 15 88 23 89
rect 106 88 136 92
rect -15 82 11 84
rect -14 80 11 82
rect 15 80 110 88
rect 128 84 136 88
rect 114 80 122 84
rect 3 76 11 80
rect 114 76 132 80
rect -17 68 -9 76
rect 6 72 132 76
rect 6 71 128 72
rect -17 46 -11 68
rect 69 59 136 67
rect 15 58 53 59
rect -7 51 53 58
rect 69 51 77 59
rect 98 51 110 59
rect -7 50 1 51
rect -17 38 23 46
rect 106 38 136 42
rect -7 26 11 34
rect 15 30 110 38
rect 128 34 136 38
rect 114 30 122 34
rect 114 26 132 30
rect 6 22 132 26
rect 6 21 128 22
rect 15 9 53 17
rect 69 9 136 17
<< labels >>
rlabel metal1 104 155 104 155 5 Vdd!
rlabel metal1 19 155 19 155 5 GND!
rlabel metal1 73 155 73 155 5 Vdd!
rlabel metal1 49 155 49 155 5 GND!
rlabel metal1 104 34 104 34 1 _ab
rlabel metal1 73 34 73 34 1 _ab
rlabel metal1 49 34 49 34 1 _ab
rlabel metal1 19 34 19 34 1 _ab
rlabel polysilicon 111 48 111 48 1 b
rlabel polysilicon 14 19 14 19 1 a
rlabel metal1 130 13 130 13 1 Vdd!
rlabel metal1 104 13 104 13 1 Vdd!
rlabel metal1 19 13 19 13 1 GND!
rlabel metal1 73 13 73 13 1 Vdd!
rlabel metal1 49 13 49 13 1 GND!
rlabel metal1 19 55 19 55 1 GND!
rlabel metal1 49 55 49 55 1 GND!
rlabel metal1 19 113 19 113 5 GND!
rlabel metal1 49 113 49 113 5 GND!
rlabel metal1 132 88 132 88 1 x
rlabel polysilicon 14 61 14 61 1 _SReset!
rlabel polysilicon 14 106 14 106 1 _SReset!
rlabel metal1 130 63 130 63 1 Vdd!
rlabel metal1 104 63 104 63 1 Vdd!
rlabel metal1 104 84 104 84 5 x
rlabel metal1 19 84 19 84 1 x
rlabel metal1 73 63 73 63 1 Vdd!
rlabel metal1 73 84 73 84 1 x
rlabel metal1 49 84 49 84 1 x
rlabel metal1 104 113 104 113 5 Vdd!
rlabel metal1 73 113 73 113 5 Vdd!
rlabel polysilicon 14 149 14 149 5 c
rlabel polysilicon 111 120 111 120 5 d
rlabel metal1 49 134 49 134 5 _cd
rlabel metal1 19 134 19 134 5 _cd
rlabel metal1 73 134 73 134 5 _cd
rlabel metal1 104 134 104 134 5 _cd
rlabel metal1 130 155 130 155 1 Vdd!
rlabel metal1 128 113 128 113 1 Vdd!
rlabel metal1 88 101 88 101 1 _cd
rlabel metal1 1 93 1 93 5 x
rlabel ndcontact -3 114 -3 114 5 GND!
rlabel metal1 -11 99 -11 99 1 GND!
rlabel metal1 -13 72 -13 72 1 _ab
rlabel metal1 -3 54 -3 54 1 GND!
rlabel polysilicon 140 105 140 105 7 _PReset!
rlabel space -20 8 46 160 7 ^n
rlabel space 76 8 144 160 3 ^p
rlabel space 32 16 45 52 3 ^nab
rlabel space 77 16 90 52 7 ^pab
rlabel space 32 58 45 110 3 ^nx
rlabel space 77 66 93 106 7 ^px
rlabel space 32 116 45 152 3 ^ncd
rlabel space 77 116 90 152 7 ^pcd
<< end >>
