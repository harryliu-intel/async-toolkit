///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Mike Jarvis <michael.a.jarvis.com> 
// -- Project Name : MBY 
// -- Description  : mgp (MeGaPort) netlist. 
// ------------------------------------------------------------------- 

module mgp (
//Input List
input                   arst_n,                                   //Asynchronous negedge reset    
input                   clk,                                      
input            [7:0]  grp_A_rx_data_valid,                      
input         [0:7][71:0]  grp_A_rx_data_w_ecc,                      
input            [7:0]  grp_A_rx_ecc,                             
input            [2:0]  grp_A_rx_flow_control_tc,                 
input           [23:0]  grp_A_rx_metadata,                        
input                   grp_A_rx_pfc_xoff,                        
input            [1:0]  grp_A_rx_port_num,                        
input           [35:0]  grp_A_rx_time_stamp,                      
input            [7:0]  grp_B_rx_data_valid,                      
input         [0:7][71:0]  grp_B_rx_data_w_ecc,                      
input            [7:0]  grp_B_rx_ecc,                             
input            [2:0]  grp_B_rx_flow_control_tc,                 
input           [23:0]  grp_B_rx_metadata,                        
input                   grp_B_rx_pfc_xoff,                        
input            [1:0]  grp_B_rx_port_num,                        
input           [35:0]  grp_B_rx_time_stamp,                      
input            [7:0]  grp_C_rx_data_valid,                      
input         [0:7][71:0]  grp_C_rx_data_w_ecc,                      
input            [7:0]  grp_C_rx_ecc,                             
input            [2:0]  grp_C_rx_flow_control_tc,                 
input           [23:0]  grp_C_rx_metadata,                        
input                   grp_C_rx_pfc_xoff,                        
input            [1:0]  grp_C_rx_port_num,                        
input           [35:0]  grp_C_rx_time_stamp,                      
input            [7:0]  grp_D_rx_data_valid,                      
input         [0:7][71:0]  grp_D_rx_data_w_ecc,                      
input            [7:0]  grp_D_rx_ecc,                             
input            [2:0]  grp_D_rx_flow_control_tc,                 
input           [23:0]  grp_D_rx_metadata,                        
input                   grp_D_rx_pfc_xoff,                        
input            [1:0]  grp_D_rx_port_num,                        
input           [35:0]  grp_D_rx_time_stamp,                      
input                   rst_n,                                    //taken from HLP active low for MBY? 
input           [19:0]  vp_cpp_rx_metadata,                       
input            [7:0]  vp_rx_data_valid,                         
input         [0:7][71:0]  vp_rx_data_w_ecc,                         
input            [7:0]  vp_rx_ecc,                                
input            [2:0]  vp_rx_flow_control_tc,                    
input           [23:0]  vp_rx_metadata,                           
input            [1:0]  vp_rx_port_num,                           
input           [35:0]  vp_rx_time_stamp,                         

//Interface List
egr_ahb_if.egr                    ahb_if,  //EGR-AHB and DFx Interface 
egr_epl_if.egr                    epl_if0,  //EGR-EPL 0 Interface 
egr_epl_if.egr                    epl_if1,  //EGR-EPL 1 Interface 
egr_epl_if.egr                    epl_if2,  //EGR-EPL 2 Interface 
egr_epl_if.egr                    epl_if3,  //EGR-EPL 3 Interface 
egr_igr_if.egr                    igr_if,  //EGR-IGR Pointer Interface 
igr_rx_ppe_if.igr                 igr_rx_ppe,  
egr_mc_table_if.egr               mc_table_if0,  //EGR-MultiCast Shared Table 0 Interface 
egr_mc_table_if.egr               mc_table_if1,  //EGR-MultiCast Shared Table 1 Interface 
egr_pod_if.egr                    pod_if,  //EGR-Pod Ring Interface 
egr_ppe_stm_if.egr                ppe_stm_if0,  //EGR-PPE Shared Table Memory 0 Interface  
egr_ppe_stm_if.egr                ppe_stm_if1,  //EGR-PPE Shared Table Memory 1 Interface 
rx_ppe_igr_if.igr                 rx_ppe_igr,  
egr_smm_readarb_if.egr            smm_readarb_if,  //EGR-SMM_Read_Arb Interface 
egr_smm_writearb_if.egr           smm_writearb_if,  //EGR-SMM_Write_Arb Interface 
egr_statsmgmt_if.egr              statsmgmt_if,  //EGR-Stats Management Interface 
egr_tagring_if.egr                tagring_if,  //EGR-Tag Ring Interface 
egr_tx_ppe_if.egr                 tx_ppe_if0,  //EGR-TxPPE 0 Interface 
egr_tx_ppe_if.egr                 tx_ppe_if1,  //EGR-TxPPE 1 Interface 
egr_vp_if.egr                     vp_if0,  //EGR-VP0 Interface 
egr_vp_if.egr                     vp_if1,  //EGR-VP1 Interface 

//Output List
output                  vp_tx_pfc_xoff                            //FIXME should this be [1:0] for 2 VP  
);



// module igr    from igr_top using igr.map 
igr_top    igr(
/* input  logic                */ .clk                      (clk),                                
/* input  logic                */ .rst_n                    (rst_n),                              //taken from HLP active low for MBY? 
/* input  logic          [7:0] */ .grp_A_rx_ecc             (grp_A_rx_ecc),                       
/* input  logic          [7:0] */ .grp_B_rx_ecc             (grp_B_rx_ecc),                       
/* input  logic          [7:0] */ .grp_C_rx_ecc             (grp_C_rx_ecc),                       
/* input  logic          [7:0] */ .grp_D_rx_ecc             (grp_D_rx_ecc),                       
/* input  logic          [1:0] */ .grp_A_rx_port_num        (grp_A_rx_port_num),                  
/* input  logic          [1:0] */ .grp_B_rx_port_num        (grp_B_rx_port_num),                  
/* input  logic          [1:0] */ .grp_C_rx_port_num        (grp_C_rx_port_num),                  
/* input  logic          [1:0] */ .grp_D_rx_port_num        (grp_D_rx_port_num),                  
/* input  logic          [7:0] */ .grp_A_rx_data_valid      (grp_A_rx_data_valid),                
/* input  logic          [7:0] */ .grp_B_rx_data_valid      (grp_B_rx_data_valid),                
/* input  logic          [7:0] */ .grp_C_rx_data_valid      (grp_C_rx_data_valid),                
/* input  logic          [7:0] */ .grp_D_rx_data_valid      (grp_D_rx_data_valid),                
/* input  logic         [23:0] */ .grp_A_rx_metadata        (grp_A_rx_metadata),                  
/* input  logic         [23:0] */ .grp_B_rx_metadata        (grp_B_rx_metadata),                  
/* input  logic         [23:0] */ .grp_C_rx_metadata        (grp_C_rx_metadata),                  
/* input  logic         [23:0] */ .grp_D_rx_metadata        (grp_D_rx_metadata),                  
/* input  logic         [35:0] */ .grp_A_rx_time_stamp      (grp_A_rx_time_stamp),                
/* input  logic         [35:0] */ .grp_B_rx_time_stamp      (grp_B_rx_time_stamp),                
/* input  logic         [35:0] */ .grp_C_rx_time_stamp      (grp_C_rx_time_stamp),                
/* input  logic         [35:0] */ .grp_D_rx_time_stamp      (grp_D_rx_time_stamp),                
/* input  logic    [0:7][71:0] */ .grp_A_rx_data_w_ecc      (grp_A_rx_data_w_ecc),                
/* input  logic    [0:7][71:0] */ .grp_B_rx_data_w_ecc      (grp_B_rx_data_w_ecc),                
/* input  logic    [0:7][71:0] */ .grp_C_rx_data_w_ecc      (grp_C_rx_data_w_ecc),                
/* input  logic    [0:7][71:0] */ .grp_D_rx_data_w_ecc      (grp_D_rx_data_w_ecc),                
/* input  logic                */ .grp_A_rx_pfc_xoff        (grp_A_rx_pfc_xoff),                  
/* input  logic                */ .grp_B_rx_pfc_xoff        (grp_B_rx_pfc_xoff),                  
/* input  logic                */ .grp_C_rx_pfc_xoff        (grp_C_rx_pfc_xoff),                  
/* input  logic                */ .grp_D_rx_pfc_xoff        (grp_D_rx_pfc_xoff),                  
/* input  logic          [2:0] */ .grp_A_rx_flow_control_tc (grp_A_rx_flow_control_tc),           
/* input  logic          [2:0] */ .grp_B_rx_flow_control_tc (grp_B_rx_flow_control_tc),           
/* input  logic          [2:0] */ .grp_C_rx_flow_control_tc (grp_C_rx_flow_control_tc),           
/* input  logic          [2:0] */ .grp_D_rx_flow_control_tc (grp_D_rx_flow_control_tc),           
/* input  logic          [7:0] */ .vp_rx_ecc                (vp_rx_ecc),                          
/* input  logic          [1:0] */ .vp_rx_port_num           (vp_rx_port_num),                     
/* input  logic          [7:0] */ .vp_rx_data_valid         (vp_rx_data_valid),                   
/* input  logic         [23:0] */ .vp_rx_metadata           (vp_rx_metadata),                     
/* input  logic         [35:0] */ .vp_rx_time_stamp         (vp_rx_time_stamp),                   
/* input  logic         [19:0] */ .vp_cpp_rx_metadata       (vp_cpp_rx_metadata),                 
/* input  logic    [0:7][71:0] */ .vp_rx_data_w_ecc         (vp_rx_data_w_ecc),                   
/* input  logic          [2:0] */ .vp_rx_flow_control_tc    (vp_rx_flow_control_tc),              
/* output logic                */ .vp_tx_pfc_xoff           (vp_tx_pfc_xoff),                     //FIXME should this be [1:0] for 2 VP  
/* Interface rx_ppe_igr_if.igr */ .rx_ppe_igr               (rx_ppe_igr),                         
/* Interface igr_rx_ppe_if.igr */ .igr_rx_ppe               (igr_rx_ppe));                         
// End of module igr from igr_top


// module egr    from egr_top using egr.map 
egr_top    egr(
/* input  logic                      */ .clk                      (clk),                                
/* input  logic                      */ .arst_n                   (arst_n),                             //Asynchronous negedge reset    
/* Interface egr_igr_if.egr          */ .igr_if                   (igr_if),                             
/* Interface egr_pod_if.egr          */ .pod_if                   (pod_if),                             
/* Interface egr_ahb_if.egr          */ .ahb_if                   (ahb_if),                             
/* Interface egr_smm_writearb_if.egr */ .smm_writearb_if          (smm_writearb_if),                    
/* Interface egr_smm_readarb_if.egr  */ .smm_readarb_if           (smm_readarb_if),                     
/* Interface egr_tagring_if.egr      */ .tagring_if               (tagring_if),                         
/* Interface egr_statsmgmt_if.egr    */ .statsmgmt_if             (statsmgmt_if),                       
/* Interface egr_tx_ppe_if.egr       */ .tx_ppe_if0               (tx_ppe_if0),                         
/* Interface egr_tx_ppe_if.egr       */ .tx_ppe_if1               (tx_ppe_if1),                         
/* Interface egr_ppe_stm_if.egr      */ .ppe_stm_if0              (ppe_stm_if0),                        
/* Interface egr_ppe_stm_if.egr      */ .ppe_stm_if1              (ppe_stm_if1),                        
/* Interface egr_epl_if.egr          */ .epl_if0                  (epl_if0),                            
/* Interface egr_epl_if.egr          */ .epl_if1                  (epl_if1),                            
/* Interface egr_epl_if.egr          */ .epl_if2                  (epl_if2),                            
/* Interface egr_epl_if.egr          */ .epl_if3                  (epl_if3),                            
/* Interface egr_vp_if.egr           */ .vp_if0                   (vp_if0),                             
/* Interface egr_vp_if.egr           */ .vp_if1                   (vp_if1),                             
/* Interface egr_mc_table_if.egr     */ .mc_table_if0             (mc_table_if0),                       
/* Interface egr_mc_table_if.egr     */ .mc_table_if1             (mc_table_if1));                       
// End of module egr from egr_top

endmodule // mgp
