magic
tech scmos
timestamp 988943070
<< nselect >>
rect -46 23 0 58
<< pselect >>
rect 0 23 70 58
<< ndiffusion >>
rect -42 44 -38 47
rect -16 37 -8 38
rect -42 33 -38 36
rect -16 33 -8 34
<< pdiffusion >>
rect 29 44 33 47
rect 58 46 66 47
rect 8 37 16 38
rect 8 33 16 34
rect 29 33 33 40
rect 58 42 66 43
<< ntransistor >>
rect -42 36 -38 44
rect -16 34 -8 37
<< ptransistor >>
rect 29 40 33 44
rect 8 34 16 37
rect 58 43 66 46
<< polysilicon >>
rect -46 36 -42 44
rect -38 37 -33 44
rect -2 37 2 46
rect 25 40 29 44
rect 33 40 37 44
rect -38 36 -25 37
rect -20 34 -16 37
rect -8 34 8 37
rect 16 34 20 37
rect 54 43 58 46
rect 66 43 70 46
<< ndcontact >>
rect -45 47 -37 55
rect -16 38 -8 46
rect -42 25 -34 33
rect -16 25 -8 33
<< pdcontact >>
rect 25 47 33 55
rect 8 38 16 46
rect 58 47 66 55
rect 58 34 66 42
rect 8 25 16 33
rect 25 25 33 33
<< polycontact >>
rect -4 46 4 54
rect -33 37 -25 45
rect 37 38 45 46
<< metal1 >>
rect -45 50 66 55
rect -45 47 -37 50
rect -4 46 4 50
rect 25 47 33 50
rect 58 47 66 50
rect -25 45 -8 46
rect -33 42 -8 45
rect 8 43 16 46
rect 37 43 45 46
rect 8 42 45 43
rect -33 41 45 42
rect -33 37 -25 41
rect -16 39 45 41
rect -16 38 16 39
rect 37 38 45 39
rect 58 33 66 42
rect -42 25 -8 33
rect 8 25 66 33
<< labels >>
rlabel metal1 -45 50 66 55 1 x
rlabel space 66 23 71 58 3 ^p
rlabel polysilicon 54 43 58 46 1 a|pin|w|3|poly
rlabel polysilicon 66 43 70 46 1 a|pin|w|3|poly
rlabel metal1 -42 25 -8 33 1 GND!
rlabel metal1 58 25 66 42 1 Vdd!
rlabel metal1 8 25 66 33 1 Vdd!
<< end >>
