magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect -1 45 7 46
rect -1 37 7 42
rect -1 29 7 34
rect -1 21 7 26
rect -1 17 7 18
<< pdiffusion >>
rect 23 50 31 51
rect 23 46 31 47
rect 23 37 31 38
rect 23 33 31 34
rect 23 24 31 25
rect 23 20 31 21
rect 31 12 39 17
rect 23 11 39 12
rect 23 7 39 8
<< ntransistor >>
rect -1 42 7 45
rect -1 34 7 37
rect -1 26 7 29
rect -1 18 7 21
<< ptransistor >>
rect 23 47 31 50
rect 23 34 31 37
rect 23 21 31 24
rect 23 8 39 11
<< polysilicon >>
rect 18 47 23 50
rect 31 47 35 50
rect 18 45 21 47
rect -5 42 -1 45
rect 7 42 21 45
rect -5 34 -1 37
rect 7 34 23 37
rect 31 34 35 37
rect -5 26 -1 29
rect 7 26 21 29
rect 18 24 21 26
rect 18 21 23 24
rect 31 21 35 24
rect -5 18 -1 21
rect 7 18 11 21
rect 19 8 23 11
rect 39 8 43 11
<< ndcontact >>
rect -1 46 7 54
rect -1 9 7 17
<< pdcontact >>
rect 23 51 31 59
rect 23 38 31 46
rect 23 25 31 33
rect 23 12 31 20
rect 23 -1 39 7
<< metal1 >>
rect -1 46 7 54
rect 23 51 31 59
rect -1 38 31 46
rect 11 20 19 38
rect 23 25 31 33
rect -1 9 7 17
rect 11 12 31 20
rect 23 -1 39 7
<< labels >>
rlabel metal1 27 16 27 16 1 x
rlabel metal1 27 55 27 55 5 Vdd!
rlabel metal1 27 29 27 29 1 Vdd!
rlabel metal1 27 42 27 42 5 x
rlabel metal1 3 13 3 13 1 GND!
rlabel metal1 3 50 3 50 1 x
rlabel polysilicon -2 43 -2 43 3 c
rlabel polysilicon -2 35 -2 35 3 b
rlabel polysilicon -2 27 -2 27 3 a
rlabel polysilicon -2 19 -2 19 3 _SReset!
rlabel polysilicon 32 48 32 48 1 c
rlabel polysilicon 32 22 32 22 1 a
rlabel polysilicon 32 35 32 35 1 b
rlabel metal1 27 3 27 3 1 Vdd!
rlabel space -6 9 -1 54 7 ^n
rlabel polysilicon 40 10 40 10 5 _PReset!
rlabel space 31 19 36 59 3 ^p
<< end >>
