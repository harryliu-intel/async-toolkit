///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_mesh_row_map_pkg.vh                                    
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_MESH_ROW_MAP_PKG_VH
`define MBY_MESH_ROW_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_mesh_row_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_mesh_row_map_cr_req_t;
typedef cfg_ack_64bit_t mby_mesh_row_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_mesh_row_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic  [7:0] WB_TO_NB;  // RW
    logic  [7:0] EB_TO_NB;  // RW
    logic  [7:0] NB_TO_NB;  // RW
    logic  [7:0] WB_TO_SB;  // RW
    logic  [7:0] EB_TO_SB;  // RW
    logic  [7:0] SB_TO_SB;  // RW
} MESH_ARB_RREQ_Y_t;

localparam MESH_ARB_RREQ_Y_REG_STRIDE = 48'h8;
localparam MESH_ARB_RREQ_Y_REG_ENTRIES = 8;
localparam [7:0][47:0] MESH_ARB_RREQ_Y_CR_ADDR = {48'h38, 48'h30, 48'h28, 48'h20, 48'h18, 48'h10, 48'h8, 48'h0};
localparam MESH_ARB_RREQ_Y_SIZE = 64;
localparam MESH_ARB_RREQ_Y_WB_TO_NB_LO = 40;
localparam MESH_ARB_RREQ_Y_WB_TO_NB_HI = 47;
localparam MESH_ARB_RREQ_Y_WB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_RREQ_Y_EB_TO_NB_LO = 32;
localparam MESH_ARB_RREQ_Y_EB_TO_NB_HI = 39;
localparam MESH_ARB_RREQ_Y_EB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_RREQ_Y_NB_TO_NB_LO = 24;
localparam MESH_ARB_RREQ_Y_NB_TO_NB_HI = 31;
localparam MESH_ARB_RREQ_Y_NB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_RREQ_Y_WB_TO_SB_LO = 16;
localparam MESH_ARB_RREQ_Y_WB_TO_SB_HI = 23;
localparam MESH_ARB_RREQ_Y_WB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_RREQ_Y_EB_TO_SB_LO = 8;
localparam MESH_ARB_RREQ_Y_EB_TO_SB_HI = 15;
localparam MESH_ARB_RREQ_Y_EB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_RREQ_Y_SB_TO_SB_LO = 0;
localparam MESH_ARB_RREQ_Y_SB_TO_SB_HI = 7;
localparam MESH_ARB_RREQ_Y_SB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_RREQ_Y_USEMASK = 64'hFFFFFFFFFFFF;
localparam MESH_ARB_RREQ_Y_RO_MASK = 64'h0;
localparam MESH_ARB_RREQ_Y_WO_MASK = 64'h0;
localparam MESH_ARB_RREQ_Y_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic  [7:0] WB_TO_NB;  // RW
    logic  [7:0] EB_TO_NB;  // RW
    logic  [7:0] NB_TO_NB;  // RW
    logic  [7:0] WB_TO_SB;  // RW
    logic  [7:0] EB_TO_SB;  // RW
    logic  [7:0] SB_TO_SB;  // RW
} MESH_ARB_WREQ_Y_t;

localparam MESH_ARB_WREQ_Y_REG_STRIDE = 48'h8;
localparam MESH_ARB_WREQ_Y_REG_ENTRIES = 8;
localparam [7:0][47:0] MESH_ARB_WREQ_Y_CR_ADDR = {48'h78, 48'h70, 48'h68, 48'h60, 48'h58, 48'h50, 48'h48, 48'h40};
localparam MESH_ARB_WREQ_Y_SIZE = 64;
localparam MESH_ARB_WREQ_Y_WB_TO_NB_LO = 40;
localparam MESH_ARB_WREQ_Y_WB_TO_NB_HI = 47;
localparam MESH_ARB_WREQ_Y_WB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_WREQ_Y_EB_TO_NB_LO = 32;
localparam MESH_ARB_WREQ_Y_EB_TO_NB_HI = 39;
localparam MESH_ARB_WREQ_Y_EB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_WREQ_Y_NB_TO_NB_LO = 24;
localparam MESH_ARB_WREQ_Y_NB_TO_NB_HI = 31;
localparam MESH_ARB_WREQ_Y_NB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_WREQ_Y_WB_TO_SB_LO = 16;
localparam MESH_ARB_WREQ_Y_WB_TO_SB_HI = 23;
localparam MESH_ARB_WREQ_Y_WB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_WREQ_Y_EB_TO_SB_LO = 8;
localparam MESH_ARB_WREQ_Y_EB_TO_SB_HI = 15;
localparam MESH_ARB_WREQ_Y_EB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_WREQ_Y_SB_TO_SB_LO = 0;
localparam MESH_ARB_WREQ_Y_SB_TO_SB_HI = 7;
localparam MESH_ARB_WREQ_Y_SB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_WREQ_Y_USEMASK = 64'hFFFFFFFFFFFF;
localparam MESH_ARB_WREQ_Y_RO_MASK = 64'h0;
localparam MESH_ARB_WREQ_Y_WO_MASK = 64'h0;
localparam MESH_ARB_WREQ_Y_RESET = 64'h0;

typedef struct packed {
    logic  [7:0] WB_TO_NB;  // RW
    logic  [7:0] EB_TO_NB;  // RW
    logic  [7:0] NB_TO_NB;  // RW
    logic  [7:0] MEM_TO_NB;  // RW
    logic  [7:0] WB_TO_SB;  // RW
    logic  [7:0] EB_TO_SB;  // RW
    logic  [7:0] SB_TO_SB;  // RW
    logic  [7:0] MEM_TO_SB;  // RW
} MESH_ARB_RRSP_Y_t;

localparam MESH_ARB_RRSP_Y_REG_STRIDE = 48'h8;
localparam MESH_ARB_RRSP_Y_REG_ENTRIES = 8;
localparam [7:0][47:0] MESH_ARB_RRSP_Y_CR_ADDR = {48'hB8, 48'hB0, 48'hA8, 48'hA0, 48'h98, 48'h90, 48'h88, 48'h80};
localparam MESH_ARB_RRSP_Y_SIZE = 64;
localparam MESH_ARB_RRSP_Y_WB_TO_NB_LO = 56;
localparam MESH_ARB_RRSP_Y_WB_TO_NB_HI = 63;
localparam MESH_ARB_RRSP_Y_WB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_EB_TO_NB_LO = 48;
localparam MESH_ARB_RRSP_Y_EB_TO_NB_HI = 55;
localparam MESH_ARB_RRSP_Y_EB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_NB_TO_NB_LO = 40;
localparam MESH_ARB_RRSP_Y_NB_TO_NB_HI = 47;
localparam MESH_ARB_RRSP_Y_NB_TO_NB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_MEM_TO_NB_LO = 32;
localparam MESH_ARB_RRSP_Y_MEM_TO_NB_HI = 39;
localparam MESH_ARB_RRSP_Y_MEM_TO_NB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_WB_TO_SB_LO = 24;
localparam MESH_ARB_RRSP_Y_WB_TO_SB_HI = 31;
localparam MESH_ARB_RRSP_Y_WB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_EB_TO_SB_LO = 16;
localparam MESH_ARB_RRSP_Y_EB_TO_SB_HI = 23;
localparam MESH_ARB_RRSP_Y_EB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_SB_TO_SB_LO = 8;
localparam MESH_ARB_RRSP_Y_SB_TO_SB_HI = 15;
localparam MESH_ARB_RRSP_Y_SB_TO_SB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_MEM_TO_SB_LO = 0;
localparam MESH_ARB_RRSP_Y_MEM_TO_SB_HI = 7;
localparam MESH_ARB_RRSP_Y_MEM_TO_SB_RESET = 8'h0;
localparam MESH_ARB_RRSP_Y_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam MESH_ARB_RRSP_Y_RO_MASK = 64'h0;
localparam MESH_ARB_RRSP_Y_WO_MASK = 64'h0;
localparam MESH_ARB_RRSP_Y_RESET = 64'h0;

typedef struct packed {
    logic  [7:0] NB_TO_WB;  // RW
    logic  [7:0] SB_TO_WB;  // RW
    logic  [7:0] WB_TO_WB;  // RW
    logic  [7:0] MEM_TO_WB;  // RW
    logic  [7:0] NB_TO_EB;  // RW
    logic  [7:0] SB_TO_EB;  // RW
    logic  [7:0] EB_TO_EB;  // RW
    logic  [7:0] MEM_TO_EB;  // RW
} MESH_ARB_RRSP_X_t;

localparam MESH_ARB_RRSP_X_REG_STRIDE = 48'h8;
localparam MESH_ARB_RRSP_X_REG_ENTRIES = 8;
localparam [7:0][47:0] MESH_ARB_RRSP_X_CR_ADDR = {48'hF8, 48'hF0, 48'hE8, 48'hE0, 48'hD8, 48'hD0, 48'hC8, 48'hC0};
localparam MESH_ARB_RRSP_X_SIZE = 64;
localparam MESH_ARB_RRSP_X_NB_TO_WB_LO = 56;
localparam MESH_ARB_RRSP_X_NB_TO_WB_HI = 63;
localparam MESH_ARB_RRSP_X_NB_TO_WB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_SB_TO_WB_LO = 48;
localparam MESH_ARB_RRSP_X_SB_TO_WB_HI = 55;
localparam MESH_ARB_RRSP_X_SB_TO_WB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_WB_TO_WB_LO = 40;
localparam MESH_ARB_RRSP_X_WB_TO_WB_HI = 47;
localparam MESH_ARB_RRSP_X_WB_TO_WB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_MEM_TO_WB_LO = 32;
localparam MESH_ARB_RRSP_X_MEM_TO_WB_HI = 39;
localparam MESH_ARB_RRSP_X_MEM_TO_WB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_NB_TO_EB_LO = 24;
localparam MESH_ARB_RRSP_X_NB_TO_EB_HI = 31;
localparam MESH_ARB_RRSP_X_NB_TO_EB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_SB_TO_EB_LO = 16;
localparam MESH_ARB_RRSP_X_SB_TO_EB_HI = 23;
localparam MESH_ARB_RRSP_X_SB_TO_EB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_EB_TO_EB_LO = 8;
localparam MESH_ARB_RRSP_X_EB_TO_EB_HI = 15;
localparam MESH_ARB_RRSP_X_EB_TO_EB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_MEM_TO_EB_LO = 0;
localparam MESH_ARB_RRSP_X_MEM_TO_EB_HI = 7;
localparam MESH_ARB_RRSP_X_MEM_TO_EB_RESET = 8'h0;
localparam MESH_ARB_RRSP_X_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam MESH_ARB_RRSP_X_RO_MASK = 64'h0;
localparam MESH_ARB_RRSP_X_WO_MASK = 64'h0;
localparam MESH_ARB_RRSP_X_RESET = 64'h0;

typedef struct packed {
    MESH_ARB_RREQ_Y_t [7:0] MESH_ARB_RREQ_Y;
    MESH_ARB_WREQ_Y_t [7:0] MESH_ARB_WREQ_Y;
    MESH_ARB_RRSP_Y_t [7:0] MESH_ARB_RRSP_Y;
    MESH_ARB_RRSP_X_t [7:0] MESH_ARB_RRSP_X;
} mby_mesh_row_map_registers_t;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_mesh_row_map_pkg

`endif // MBY_MESH_ROW_MAP_PKG_VH
