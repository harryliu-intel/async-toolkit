magic
tech scmos
timestamp 965071348
<< ndiffusion >>
rect -52 33 -44 34
rect -78 19 -66 20
rect -52 29 -44 30
rect -52 20 -44 21
rect -78 11 -66 16
rect -78 7 -66 8
rect -78 -2 -66 -1
rect -52 16 -44 17
rect -52 7 -44 8
rect -52 3 -44 4
rect -52 -6 -44 -5
rect -52 -10 -44 -9
<< pdiffusion >>
rect -122 33 -112 34
rect -28 33 -20 34
rect -122 29 -112 30
rect -122 20 -112 21
rect -122 16 -112 17
rect -28 29 -20 30
rect -28 20 -20 21
rect -114 8 -112 16
rect -98 13 -94 16
rect -122 7 -112 8
rect -98 7 -94 10
rect -122 3 -112 4
rect -122 -6 -112 -5
rect -102 -2 -94 -1
rect -122 -10 -112 -9
rect -28 16 -20 17
rect -28 7 -20 8
rect -28 3 -20 4
rect -28 -6 -20 -5
rect -28 -10 -20 -9
<< ntransistor >>
rect -52 30 -44 33
rect -78 16 -66 19
rect -52 17 -44 20
rect -78 8 -66 11
rect -52 4 -44 7
rect -52 -9 -44 -6
<< ptransistor >>
rect -122 30 -112 33
rect -122 17 -112 20
rect -28 30 -20 33
rect -28 17 -20 20
rect -98 10 -94 13
rect -122 4 -112 7
rect -122 -9 -112 -6
rect -28 4 -20 7
rect -28 -9 -20 -6
<< polysilicon >>
rect -127 30 -122 33
rect -112 30 -80 33
rect -57 32 -52 33
rect -127 20 -124 30
rect -127 17 -122 20
rect -112 17 -108 20
rect -127 7 -124 17
rect -83 19 -80 30
rect -56 30 -52 32
rect -44 30 -28 33
rect -20 30 -16 33
rect -56 24 -54 30
rect -57 20 -54 24
rect -83 16 -78 19
rect -66 16 -62 19
rect -57 17 -52 20
rect -44 17 -28 20
rect -20 17 -16 20
rect -102 10 -98 13
rect -94 11 -88 13
rect -94 10 -90 11
rect -91 7 -90 10
rect -127 4 -122 7
rect -112 4 -108 7
rect -127 -6 -124 4
rect -82 8 -78 11
rect -66 8 -62 11
rect -127 -9 -122 -6
rect -112 -9 -108 -6
rect -57 7 -54 17
rect -57 4 -52 7
rect -44 4 -28 7
rect -20 4 -16 7
rect -57 -6 -54 4
rect -57 -9 -52 -6
rect -44 -9 -28 -6
rect -20 -9 -16 -6
<< ndcontact >>
rect -52 34 -44 42
rect -78 20 -66 28
rect -52 21 -44 29
rect -78 -1 -66 7
rect -52 8 -44 16
rect -52 -5 -44 3
rect -52 -18 -44 -10
<< pdcontact >>
rect -122 34 -112 42
rect -28 34 -20 42
rect -122 21 -112 29
rect -102 16 -94 24
rect -28 21 -20 29
rect -122 8 -114 16
rect -122 -5 -112 3
rect -102 -1 -94 7
rect -28 8 -20 16
rect -28 -5 -20 3
rect -122 -18 -112 -10
rect -28 -18 -20 -10
<< psubstratepcontact >>
rect -78 -10 -66 -2
<< nsubstratencontact >>
rect -102 -10 -94 -2
<< polycontact >>
rect -64 24 -56 32
rect -90 3 -82 11
<< metal1 >>
rect -122 34 -112 42
rect -52 34 -44 42
rect -28 34 -20 42
rect -122 25 -112 29
rect -64 28 -56 32
rect -78 25 -56 28
rect -122 24 -56 25
rect -122 23 -57 24
rect -122 21 -66 23
rect -52 21 -20 29
rect -110 20 -66 21
rect -110 17 -94 20
rect -122 8 -114 16
rect -110 3 -106 17
rect -102 16 -94 17
rect -86 11 -57 15
rect -122 -1 -106 3
rect -122 -5 -112 -1
rect -102 -10 -94 7
rect -90 3 -82 11
rect -122 -18 -94 -10
rect -78 -10 -66 7
rect -61 3 -57 11
rect -52 8 -44 16
rect -40 3 -32 21
rect -28 8 -20 16
rect -61 -1 -20 3
rect -52 -5 -20 -1
rect -78 -18 -44 -10
rect -28 -18 -20 -10
<< labels >>
rlabel metal1 -74 -6 -74 -6 1 GND!
rlabel metal1 -74 3 -74 3 1 GND!
rlabel metal1 -98 -6 -98 -6 1 Vdd!
rlabel metal1 -98 3 -98 3 1 Vdd!
rlabel polysilicon -99 11 -99 11 1 x
rlabel metal1 -74 24 -74 24 1 _x
rlabel polysilicon -79 9 -79 9 1 x
rlabel polysilicon -79 17 -79 17 1 a
rlabel polysilicon -123 -7 -123 -7 5 a
rlabel polysilicon -123 6 -123 6 5 a
rlabel metal1 -118 -14 -118 -14 1 Vdd!
rlabel polysilicon -123 31 -123 31 1 a
rlabel polysilicon -123 18 -123 18 1 a
rlabel metal1 -118 38 -118 38 5 Vdd!
rlabel metal1 -118 12 -118 12 1 Vdd!
rlabel metal1 -117 25 -117 25 1 _x
rlabel metal1 -117 -1 -117 -1 5 _x
rlabel pdcontact -24 -1 -24 -1 5 x
rlabel pdcontact -24 -14 -24 -14 1 Vdd!
rlabel polysilicon -19 -7 -19 -7 5 _x
rlabel polysilicon -19 6 -19 6 5 _x
rlabel polysilicon -53 -7 -53 -7 3 _x
rlabel polysilicon -53 6 -53 6 3 _x
rlabel ndcontact -48 -14 -48 -14 1 GND!
rlabel ndcontact -48 -1 -48 -1 5 x
rlabel pdcontact -24 12 -24 12 1 Vdd!
rlabel pdcontact -24 25 -24 25 1 x
rlabel pdcontact -24 38 -24 38 5 Vdd!
rlabel polysilicon -19 31 -19 31 1 _x
rlabel polysilicon -19 18 -19 18 1 _x
rlabel polysilicon -53 31 -53 31 3 _x
rlabel polysilicon -53 18 -53 18 3 _x
rlabel ndcontact -48 38 -48 38 5 GND!
rlabel ndcontact -48 12 -48 12 1 GND!
rlabel ndcontact -48 25 -48 25 1 x
rlabel metal1 -98 20 -98 20 1 _x
rlabel space -128 -18 -122 42 7 ^p1
rlabel space -20 -18 -15 42 3 ^p2
rlabel space -44 -19 -14 43 3 ^n2
<< end >>
