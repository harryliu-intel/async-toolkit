magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect -191 -696 -183 -695
rect -191 -704 -183 -699
rect -191 -712 -183 -707
rect -191 -720 -183 -715
rect -191 -728 -183 -723
rect -191 -732 -183 -731
rect -191 -741 -183 -740
rect -191 -749 -183 -744
rect -191 -757 -183 -752
rect -191 -765 -183 -760
rect -191 -773 -183 -768
rect -191 -777 -183 -776
<< pdiffusion >>
rect -167 -676 -159 -675
rect -167 -680 -159 -679
rect -167 -689 -159 -688
rect -167 -693 -159 -692
rect -167 -702 -159 -701
rect -167 -706 -159 -705
rect -167 -715 -159 -714
rect -167 -719 -159 -718
rect -167 -728 -159 -727
rect -167 -732 -159 -731
rect -167 -741 -159 -740
rect -167 -745 -159 -744
rect -167 -754 -159 -753
rect -167 -758 -159 -757
rect -167 -767 -159 -766
rect -167 -771 -159 -770
rect -167 -780 -159 -779
rect -167 -784 -159 -783
rect -167 -793 -159 -792
rect -167 -797 -159 -796
<< ntransistor >>
rect -191 -699 -183 -696
rect -191 -707 -183 -704
rect -191 -715 -183 -712
rect -191 -723 -183 -720
rect -191 -731 -183 -728
rect -191 -744 -183 -741
rect -191 -752 -183 -749
rect -191 -760 -183 -757
rect -191 -768 -183 -765
rect -191 -776 -183 -773
<< ptransistor >>
rect -167 -679 -159 -676
rect -167 -692 -159 -689
rect -167 -705 -159 -702
rect -167 -718 -159 -715
rect -167 -731 -159 -728
rect -167 -744 -159 -741
rect -167 -757 -159 -754
rect -167 -770 -159 -767
rect -167 -783 -159 -780
rect -167 -796 -159 -793
<< polysilicon >>
rect -181 -679 -167 -676
rect -159 -679 -155 -676
rect -181 -696 -178 -679
rect -195 -699 -191 -696
rect -183 -699 -178 -696
rect -172 -692 -167 -689
rect -159 -692 -155 -689
rect -172 -702 -169 -692
rect -172 -704 -167 -702
rect -195 -707 -191 -704
rect -183 -705 -167 -704
rect -159 -705 -155 -702
rect -183 -707 -169 -705
rect -195 -715 -191 -712
rect -183 -715 -169 -712
rect -172 -718 -167 -715
rect -159 -718 -155 -715
rect -195 -723 -191 -720
rect -183 -723 -179 -720
rect -195 -731 -191 -728
rect -183 -731 -167 -728
rect -159 -731 -155 -728
rect -195 -744 -191 -741
rect -183 -744 -167 -741
rect -159 -744 -155 -741
rect -195 -752 -191 -749
rect -183 -752 -179 -749
rect -172 -757 -167 -754
rect -159 -757 -155 -754
rect -195 -760 -191 -757
rect -183 -760 -169 -757
rect -195 -768 -191 -765
rect -183 -767 -169 -765
rect -183 -768 -167 -767
rect -172 -770 -167 -768
rect -159 -770 -155 -767
rect -195 -776 -191 -773
rect -183 -776 -178 -773
rect -181 -793 -178 -776
rect -172 -780 -169 -770
rect -172 -783 -167 -780
rect -159 -783 -155 -780
rect -181 -796 -167 -793
rect -159 -796 -155 -793
<< ndcontact >>
rect -191 -695 -183 -687
rect -191 -740 -183 -732
rect -191 -785 -183 -777
<< pdcontact >>
rect -167 -675 -159 -667
rect -167 -688 -159 -680
rect -167 -701 -159 -693
rect -167 -714 -159 -706
rect -167 -727 -159 -719
rect -167 -740 -159 -732
rect -167 -753 -159 -745
rect -167 -766 -159 -758
rect -167 -779 -159 -771
rect -167 -792 -159 -784
rect -167 -805 -159 -797
<< metal1 >>
rect -167 -675 -159 -667
rect -191 -695 -183 -687
rect -179 -688 -159 -680
rect -179 -706 -171 -688
rect -167 -701 -159 -693
rect -179 -714 -159 -706
rect -179 -732 -171 -714
rect -167 -727 -159 -719
rect -191 -740 -159 -732
rect -179 -758 -171 -740
rect -167 -753 -159 -745
rect -179 -766 -159 -758
rect -191 -785 -183 -777
rect -179 -784 -171 -766
rect -167 -779 -159 -771
rect -179 -792 -159 -784
rect -167 -805 -159 -797
<< labels >>
rlabel metal1 -163 -722 -163 -722 5 Vdd!
rlabel metal1 -163 -748 -163 -748 5 Vdd!
rlabel metal1 -163 -801 -163 -801 1 Vdd!
rlabel metal1 -163 -710 -163 -710 5 x
rlabel metal1 -163 -672 -163 -672 1 Vdd!
rlabel metal1 -163 -684 -163 -684 5 x
rlabel polysilicon -192 -730 -192 -730 3 a
rlabel polysilicon -192 -722 -192 -722 3 b
rlabel polysilicon -192 -714 -192 -714 3 c
rlabel metal1 -187 -736 -187 -736 5 x
rlabel polysilicon -192 -706 -192 -706 1 d
rlabel metal1 -187 -691 -187 -691 5 GND!
rlabel metal1 -187 -781 -187 -781 1 GND!
rlabel polysilicon -192 -759 -192 -759 3 c
rlabel polysilicon -192 -767 -192 -767 3 b
rlabel polysilicon -192 -775 -192 -775 3 a
rlabel polysilicon -192 -751 -192 -751 1 d
rlabel polysilicon -192 -743 -192 -743 3 e
rlabel polysilicon -192 -698 -192 -698 3 e
rlabel metal1 -163 -697 -163 -697 1 Vdd!
rlabel metal1 -163 -736 -163 -736 1 x
rlabel metal1 -163 -762 -163 -762 5 x
rlabel metal1 -163 -788 -163 -788 1 x
rlabel metal1 -163 -775 -163 -775 1 Vdd!
rlabel polysilicon -158 -678 -158 -678 7 e
rlabel polysilicon -158 -743 -158 -743 7 e
rlabel polysilicon -158 -795 -158 -795 7 a
rlabel polysilicon -158 -730 -158 -730 7 a
rlabel polysilicon -158 -717 -158 -717 7 c
rlabel polysilicon -158 -756 -158 -756 7 c
rlabel polysilicon -158 -782 -158 -782 7 b
rlabel polysilicon -158 -769 -158 -769 7 b
rlabel polysilicon -158 -704 -158 -704 7 d
rlabel polysilicon -158 -691 -158 -691 7 d
rlabel space -196 -785 -191 -687 7 ^n
rlabel space -159 -805 -154 -667 3 ^p
<< end >>
