magic
tech scmos
timestamp 970031125
<< ndiffusion >>
rect -25 22 -13 23
rect -25 14 -13 19
rect -25 10 -13 11
rect -25 2 -23 10
rect -25 1 -13 2
rect -47 -7 -39 -6
rect -25 -7 -13 -2
rect -47 -11 -39 -10
rect -25 -11 -13 -10
<< pdiffusion >>
rect 8 22 24 23
rect 8 14 24 19
rect 55 21 59 24
rect 55 15 59 18
rect 8 10 24 11
rect 8 1 24 2
rect 8 -7 24 -2
rect 53 -7 61 -6
rect 8 -11 24 -10
rect 53 -11 61 -10
<< ntransistor >>
rect -25 19 -13 22
rect -25 11 -13 14
rect -25 -2 -13 1
rect -47 -10 -39 -7
rect -25 -10 -13 -7
<< ptransistor >>
rect 8 19 24 22
rect 55 18 59 21
rect 8 11 24 14
rect 8 -2 24 1
rect 8 -10 24 -7
rect 53 -10 61 -7
<< polysilicon >>
rect -29 19 -25 22
rect -13 19 8 22
rect 24 19 33 22
rect 51 18 55 21
rect 59 18 63 21
rect -30 11 -25 14
rect -13 11 -9 14
rect -52 -7 -49 10
rect -30 6 -27 11
rect 4 11 8 14
rect 24 11 28 14
rect -27 -2 -25 1
rect -13 -2 -9 1
rect -4 -7 -1 6
rect 33 1 36 14
rect 4 -2 8 1
rect 24 -2 36 1
rect 46 -7 49 1
rect -52 -10 -47 -7
rect -39 -10 -35 -7
rect -29 -10 -25 -7
rect -13 -10 8 -7
rect 24 -10 28 -7
rect 46 -10 53 -7
rect 61 -10 65 -7
<< ndcontact >>
rect -25 23 -13 31
rect -47 -6 -39 2
rect -23 2 -13 10
rect -47 -19 -39 -11
rect -25 -19 -13 -11
<< pdcontact >>
rect 8 23 24 31
rect 51 24 59 32
rect 8 2 24 10
rect 51 7 59 15
rect 53 -6 61 2
rect 8 -19 24 -11
rect 53 -19 61 -11
<< psubstratepcontact >>
rect -42 23 -34 31
<< nsubstratencontact >>
rect 33 -19 41 -11
<< polycontact >>
rect -52 10 -44 18
rect 33 14 41 22
rect -35 -2 -27 6
rect -4 6 4 14
rect 41 1 49 9
rect 63 13 71 21
<< metal1 >>
rect -42 27 -21 31
rect 51 31 59 32
rect 21 27 59 31
rect -42 23 -13 27
rect 8 26 59 27
rect 8 23 24 26
rect 51 24 59 26
rect 33 21 41 22
rect -52 14 -44 18
rect -52 10 -19 14
rect -23 9 -13 10
rect -35 2 -27 6
rect -4 6 4 15
rect 33 14 41 15
rect 51 11 59 15
rect 8 9 24 10
rect 45 9 59 11
rect -23 2 -13 3
rect 8 2 24 3
rect 49 7 59 9
rect 63 13 71 21
rect -47 -2 -27 2
rect 41 1 49 3
rect 63 2 67 13
rect -47 -6 -39 -2
rect -31 -3 -27 -2
rect 53 -2 67 2
rect 53 -3 61 -2
rect -31 -6 61 -3
rect -31 -7 58 -6
rect -47 -15 -13 -11
rect -47 -19 -21 -15
rect 8 -15 61 -11
rect 21 -19 61 -15
<< m2contact >>
rect -21 27 -3 33
rect 3 27 21 33
rect -4 15 4 21
rect -23 3 -13 9
rect 33 15 41 21
rect 8 3 24 9
rect 41 3 49 9
rect -21 -21 -13 -15
rect 8 -21 21 -15
<< metal2 >>
rect -27 15 4 21
rect 27 15 41 21
rect -23 3 49 9
<< m3contact >>
rect -21 27 -3 33
rect 3 27 21 33
rect -21 -21 -3 -15
rect 3 -21 21 -15
<< metal3 >>
rect -21 -24 -3 36
rect 3 -24 21 36
<< labels >>
rlabel metal1 -19 -15 -19 -15 1 GND!
rlabel metal1 -19 27 -19 27 5 GND!
rlabel metal1 -43 -15 -43 -15 1 GND!
rlabel polysilicon -38 -9 -38 -9 1 x
rlabel metal1 20 27 20 27 5 Vdd!
rlabel metal1 20 -15 20 -15 1 Vdd!
rlabel polysilicon 25 -9 25 -9 1 a
rlabel polysilicon 25 -1 25 -1 1 b
rlabel polysilicon 25 12 25 12 1 a
rlabel polysilicon 25 20 25 20 1 b
rlabel polysilicon 49 -8 49 -8 5 x
rlabel metal1 55 11 55 11 5 x
rlabel metal1 57 -15 57 -15 5 Vdd!
rlabel metal1 37 -15 37 -15 1 Vdd!
rlabel metal1 -38 27 -38 27 1 GND!
rlabel metal2 0 3 0 9 1 x
rlabel metal2 37 18 37 18 1 b
rlabel metal2 -27 15 -27 21 3 a
rlabel metal1 55 28 55 28 5 Vdd!
rlabel space 23 -20 72 33 3 ^p
rlabel metal2 27 15 27 21 7 ^p
rlabel metal2 45 6 45 6 1 x
<< end >>
