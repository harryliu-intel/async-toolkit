magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 51 44 57 45
rect 51 41 57 42
rect 51 37 53 41
rect 51 36 57 37
rect 51 33 57 34
rect 51 28 57 29
rect 51 25 57 26
rect 51 21 53 25
rect 51 20 57 21
rect 51 17 57 18
rect 51 12 57 13
rect 51 9 57 10
rect 51 5 53 9
rect 51 4 57 5
rect 51 1 57 2
<< pdiffusion >>
rect 69 44 79 45
rect 69 41 79 42
rect 77 37 79 41
rect 69 36 79 37
rect 69 33 79 34
rect 69 29 75 33
rect 69 28 79 29
rect 69 25 79 26
rect 77 21 79 25
rect 69 20 79 21
rect 69 17 79 18
rect 69 13 75 17
rect 69 12 79 13
rect 69 9 79 10
rect 77 5 79 9
rect 69 4 79 5
rect 69 1 79 2
<< ntransistor >>
rect 51 42 57 44
rect 51 34 57 36
rect 51 26 57 28
rect 51 18 57 20
rect 51 10 57 12
rect 51 2 57 4
<< ptransistor >>
rect 69 42 79 44
rect 69 34 79 36
rect 69 26 79 28
rect 69 18 79 20
rect 69 10 79 12
rect 69 2 79 4
<< polysilicon >>
rect 47 42 51 44
rect 57 42 69 44
rect 79 42 83 44
rect 47 36 49 42
rect 62 36 64 42
rect 81 36 83 42
rect 47 34 51 36
rect 57 34 69 36
rect 79 34 83 36
rect 47 28 49 34
rect 62 28 64 34
rect 81 28 83 34
rect 47 26 51 28
rect 57 26 69 28
rect 79 26 83 28
rect 47 20 49 26
rect 62 20 64 26
rect 81 20 83 26
rect 47 18 51 20
rect 57 18 69 20
rect 79 18 83 20
rect 47 12 49 18
rect 62 12 64 18
rect 81 12 83 18
rect 47 10 51 12
rect 57 10 69 12
rect 79 10 83 12
rect 47 4 49 10
rect 62 4 64 10
rect 81 4 83 10
rect 47 2 51 4
rect 57 2 69 4
rect 79 2 83 4
<< ndcontact >>
rect 51 45 57 49
rect 53 37 57 41
rect 51 29 57 33
rect 53 21 57 25
rect 51 13 57 17
rect 53 5 57 9
rect 51 -3 57 1
<< pdcontact >>
rect 69 45 79 49
rect 69 37 77 41
rect 75 29 79 33
rect 69 21 77 25
rect 75 13 79 17
rect 69 5 77 9
rect 69 -3 79 1
<< metal1 >>
rect 51 45 57 49
rect 69 45 79 49
rect 53 37 77 41
rect 51 29 57 33
rect 69 25 72 37
rect 75 29 79 33
rect 53 21 77 25
rect 51 13 57 17
rect 69 9 72 21
rect 75 13 79 17
rect 53 5 77 9
rect 51 -3 57 1
rect 69 -3 79 1
<< labels >>
rlabel space 47 -4 54 50 7 ^n
rlabel space 76 -4 83 50 3 ^p
rlabel polysilicon 48 3 48 3 3 a
rlabel polysilicon 48 43 48 43 3 a
rlabel polysilicon 82 3 82 3 7 a
rlabel polysilicon 82 43 82 43 7 a
rlabel ndcontact 55 15 55 15 5 GND!
rlabel ndcontact 55 -1 55 -1 1 GND!
rlabel ndcontact 55 23 55 23 1 x
rlabel ndcontact 55 7 55 7 1 x
rlabel ndcontact 55 31 55 31 5 GND!
rlabel ndcontact 55 47 55 47 5 GND!
rlabel ndcontact 55 39 55 39 1 x
rlabel pdcontact 71 23 71 23 1 x
rlabel pdcontact 71 39 71 39 1 x
rlabel pdcontact 71 7 71 7 1 x
rlabel pdcontact 77 15 77 15 5 Vdd!
rlabel pdcontact 77 31 77 31 5 Vdd!
rlabel pdcontact 77 -1 77 -1 1 Vdd!
rlabel pdcontact 77 47 77 47 5 Vdd!
<< end >>
