///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_nexthop_map_pkg.vh                                 
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_NEXTHOP_MAP_PKG_VH
`define MBY_PPE_NEXTHOP_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_nexthop_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_nexthop_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_nexthop_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_nexthop_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [53:0] reserved0;  // RSVD
    logic  [7:0] SWEEPER_RATE;  // RW
    logic  [0:0] FLOWLET_INT_EN;  // RW
    logic  [0:0] FLOWLET_ENABLE;  // RW
} NH_CONFIG_t;

localparam NH_CONFIG_REG_STRIDE = 48'h8;
localparam NH_CONFIG_REG_ENTRIES = 1;
localparam NH_CONFIG_CR_ADDR = 48'h0;
localparam NH_CONFIG_SIZE = 64;
localparam NH_CONFIG_SWEEPER_RATE_LO = 2;
localparam NH_CONFIG_SWEEPER_RATE_HI = 9;
localparam NH_CONFIG_SWEEPER_RATE_RESET = 8'h0;
localparam NH_CONFIG_FLOWLET_INT_EN_LO = 1;
localparam NH_CONFIG_FLOWLET_INT_EN_HI = 1;
localparam NH_CONFIG_FLOWLET_INT_EN_RESET = 1'h0;
localparam NH_CONFIG_FLOWLET_ENABLE_LO = 0;
localparam NH_CONFIG_FLOWLET_ENABLE_HI = 0;
localparam NH_CONFIG_FLOWLET_ENABLE_RESET = 1'h0;
localparam NH_CONFIG_USEMASK = 64'h3FF;
localparam NH_CONFIG_RO_MASK = 64'h0;
localparam NH_CONFIG_WO_MASK = 64'h0;
localparam NH_CONFIG_RESET = 64'h0;

typedef struct packed {
    logic [49:0] reserved0;  // RSVD
    logic [13:0] FLOWLET;  // RW
} NH_STATUS_t;

localparam NH_STATUS_REG_STRIDE = 48'h8;
localparam NH_STATUS_REG_ENTRIES = 1;
localparam NH_STATUS_CR_ADDR = 48'h8;
localparam NH_STATUS_SIZE = 64;
localparam NH_STATUS_FLOWLET_LO = 0;
localparam NH_STATUS_FLOWLET_HI = 13;
localparam NH_STATUS_FLOWLET_RESET = 14'h0;
localparam NH_STATUS_USEMASK = 64'h3FFF;
localparam NH_STATUS_RO_MASK = 64'h0;
localparam NH_STATUS_WO_MASK = 64'h0;
localparam NH_STATUS_RESET = 64'h0;

typedef struct packed {
    logic [15:0] DGLORT;  // RW
    logic [47:0] DST_MAC;  // RW
} NH_NEIGHBORS_0_t;

localparam NH_NEIGHBORS_0_REG_STRIDE = 48'h8;
localparam NH_NEIGHBORS_0_REG_ENTRIES = 16384;
localparam NH_NEIGHBORS_0_CR_ADDR = 48'h20000;
localparam NH_NEIGHBORS_0_SIZE = 64;
localparam NH_NEIGHBORS_0_DGLORT_LO = 48;
localparam NH_NEIGHBORS_0_DGLORT_HI = 63;
localparam NH_NEIGHBORS_0_DGLORT_RESET = 16'h0;
localparam NH_NEIGHBORS_0_DST_MAC_LO = 0;
localparam NH_NEIGHBORS_0_DST_MAC_HI = 47;
localparam NH_NEIGHBORS_0_DST_MAC_RESET = 48'h0;
localparam NH_NEIGHBORS_0_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam NH_NEIGHBORS_0_RO_MASK = 64'h0;
localparam NH_NEIGHBORS_0_WO_MASK = 64'h0;
localparam NH_NEIGHBORS_0_RESET = 64'h0;

typedef struct packed {
    logic  [5:0] reserved0;  // RSVD
    logic  [0:0] ENTRY_TYPE;  // RW
    logic  [0:0] IPV6_ENTRY;  // RW
    logic  [0:0] MARK_ROUTED;  // RW
    logic  [0:0] UPDATE_L3_DOMAIN;  // RW
    logic  [0:0] UPDATE_L2_DOMAIN;  // RW
    logic  [5:0] L3_DOMAIN;  // RW
    logic  [7:0] L2_DOMAIN;  // RW
    logic [23:0] MOD_IDX;  // RW
    logic  [2:0] MTU_INDEX;  // RW
    logic [11:0] EVID;  // RW
} NH_NEIGHBORS_1_t;

localparam NH_NEIGHBORS_1_REG_STRIDE = 48'h8;
localparam NH_NEIGHBORS_1_REG_ENTRIES = 16384;
localparam NH_NEIGHBORS_1_CR_ADDR = 48'h40000;
localparam NH_NEIGHBORS_1_SIZE = 64;
localparam NH_NEIGHBORS_1_ENTRY_TYPE_LO = 57;
localparam NH_NEIGHBORS_1_ENTRY_TYPE_HI = 57;
localparam NH_NEIGHBORS_1_ENTRY_TYPE_RESET = 1'h0;
localparam NH_NEIGHBORS_1_IPV6_ENTRY_LO = 56;
localparam NH_NEIGHBORS_1_IPV6_ENTRY_HI = 56;
localparam NH_NEIGHBORS_1_IPV6_ENTRY_RESET = 1'h0;
localparam NH_NEIGHBORS_1_MARK_ROUTED_LO = 55;
localparam NH_NEIGHBORS_1_MARK_ROUTED_HI = 55;
localparam NH_NEIGHBORS_1_MARK_ROUTED_RESET = 1'h0;
localparam NH_NEIGHBORS_1_UPDATE_L3_DOMAIN_LO = 54;
localparam NH_NEIGHBORS_1_UPDATE_L3_DOMAIN_HI = 54;
localparam NH_NEIGHBORS_1_UPDATE_L3_DOMAIN_RESET = 1'h0;
localparam NH_NEIGHBORS_1_UPDATE_L2_DOMAIN_LO = 53;
localparam NH_NEIGHBORS_1_UPDATE_L2_DOMAIN_HI = 53;
localparam NH_NEIGHBORS_1_UPDATE_L2_DOMAIN_RESET = 1'h0;
localparam NH_NEIGHBORS_1_L3_DOMAIN_LO = 47;
localparam NH_NEIGHBORS_1_L3_DOMAIN_HI = 52;
localparam NH_NEIGHBORS_1_L3_DOMAIN_RESET = 6'h0;
localparam NH_NEIGHBORS_1_L2_DOMAIN_LO = 39;
localparam NH_NEIGHBORS_1_L2_DOMAIN_HI = 46;
localparam NH_NEIGHBORS_1_L2_DOMAIN_RESET = 8'h0;
localparam NH_NEIGHBORS_1_MOD_IDX_LO = 15;
localparam NH_NEIGHBORS_1_MOD_IDX_HI = 38;
localparam NH_NEIGHBORS_1_MOD_IDX_RESET = 24'h0;
localparam NH_NEIGHBORS_1_MTU_INDEX_LO = 12;
localparam NH_NEIGHBORS_1_MTU_INDEX_HI = 14;
localparam NH_NEIGHBORS_1_MTU_INDEX_RESET = 3'h0;
localparam NH_NEIGHBORS_1_EVID_LO = 0;
localparam NH_NEIGHBORS_1_EVID_HI = 11;
localparam NH_NEIGHBORS_1_EVID_RESET = 12'h0;
localparam NH_NEIGHBORS_1_USEMASK = 64'h3FFFFFFFFFFFFFF;
localparam NH_NEIGHBORS_1_RO_MASK = 64'h0;
localparam NH_NEIGHBORS_1_WO_MASK = 64'h0;
localparam NH_NEIGHBORS_1_RESET = 64'h0;

typedef struct packed {
    logic [23:0] reserved0;  // RSVD
    logic  [5:0] WEIGHT_ROW_OFFSET;  // RW
    logic [10:0] WEIGHT_ROW;  // RW
    logic  [5:0] N_GROUP_SIZE;  // RW
    logic  [0:0] N_GROUP_SZ_TYPE;  // RW
    logic [13:0] BASE_INDEX;  // RW
    logic  [1:0] GROUP_TYPE;  // RW
} NH_GROUPS_0_t;

localparam NH_GROUPS_0_REG_STRIDE = 48'h8;
localparam NH_GROUPS_0_REG_ENTRIES = 4096;
localparam NH_GROUPS_0_CR_ADDR = 48'h60000;
localparam NH_GROUPS_0_SIZE = 64;
localparam NH_GROUPS_0_WEIGHT_ROW_OFFSET_LO = 34;
localparam NH_GROUPS_0_WEIGHT_ROW_OFFSET_HI = 39;
localparam NH_GROUPS_0_WEIGHT_ROW_OFFSET_RESET = 6'h0;
localparam NH_GROUPS_0_WEIGHT_ROW_LO = 23;
localparam NH_GROUPS_0_WEIGHT_ROW_HI = 33;
localparam NH_GROUPS_0_WEIGHT_ROW_RESET = 11'h0;
localparam NH_GROUPS_0_N_GROUP_SIZE_LO = 17;
localparam NH_GROUPS_0_N_GROUP_SIZE_HI = 22;
localparam NH_GROUPS_0_N_GROUP_SIZE_RESET = 6'h0;
localparam NH_GROUPS_0_N_GROUP_SZ_TYPE_LO = 16;
localparam NH_GROUPS_0_N_GROUP_SZ_TYPE_HI = 16;
localparam NH_GROUPS_0_N_GROUP_SZ_TYPE_RESET = 1'h0;
localparam NH_GROUPS_0_BASE_INDEX_LO = 2;
localparam NH_GROUPS_0_BASE_INDEX_HI = 15;
localparam NH_GROUPS_0_BASE_INDEX_RESET = 14'h0;
localparam NH_GROUPS_0_GROUP_TYPE_LO = 0;
localparam NH_GROUPS_0_GROUP_TYPE_HI = 1;
localparam NH_GROUPS_0_GROUP_TYPE_RESET = 2'h0;
localparam NH_GROUPS_0_USEMASK = 64'hFFFFFFFFFF;
localparam NH_GROUPS_0_RO_MASK = 64'h0;
localparam NH_GROUPS_0_WO_MASK = 64'h0;
localparam NH_GROUPS_0_RESET = 64'h0;

typedef struct packed {
    logic [34:0] reserved0;  // RSVD
    logic [10:0] GROUP_MIN_INDEX;  // RW
    logic  [7:0] FLOWLET_AGE_RESET;  // RW
    logic  [2:0] FLOWLET_POLICY;  // RW
    logic  [5:0] R_GROUP_SIZE;  // RW
    logic  [0:0] R_GROUP_SZ_TYPE;  // RW
} NH_GROUPS_1_t;

localparam NH_GROUPS_1_REG_STRIDE = 48'h8;
localparam NH_GROUPS_1_REG_ENTRIES = 4096;
localparam NH_GROUPS_1_CR_ADDR = 48'h68000;
localparam NH_GROUPS_1_SIZE = 64;
localparam NH_GROUPS_1_GROUP_MIN_INDEX_LO = 18;
localparam NH_GROUPS_1_GROUP_MIN_INDEX_HI = 28;
localparam NH_GROUPS_1_GROUP_MIN_INDEX_RESET = 11'h0;
localparam NH_GROUPS_1_FLOWLET_AGE_RESET_LO = 10;
localparam NH_GROUPS_1_FLOWLET_AGE_RESET_HI = 17;
localparam NH_GROUPS_1_FLOWLET_AGE_RESET_RESET = 8'h0;
localparam NH_GROUPS_1_FLOWLET_POLICY_LO = 7;
localparam NH_GROUPS_1_FLOWLET_POLICY_HI = 9;
localparam NH_GROUPS_1_FLOWLET_POLICY_RESET = 3'h0;
localparam NH_GROUPS_1_R_GROUP_SIZE_LO = 1;
localparam NH_GROUPS_1_R_GROUP_SIZE_HI = 6;
localparam NH_GROUPS_1_R_GROUP_SIZE_RESET = 6'h0;
localparam NH_GROUPS_1_R_GROUP_SZ_TYPE_LO = 0;
localparam NH_GROUPS_1_R_GROUP_SZ_TYPE_HI = 0;
localparam NH_GROUPS_1_R_GROUP_SZ_TYPE_RESET = 1'h0;
localparam NH_GROUPS_1_USEMASK = 64'h1FFFFFFF;
localparam NH_GROUPS_1_RO_MASK = 64'h0;
localparam NH_GROUPS_1_WO_MASK = 64'h0;
localparam NH_GROUPS_1_RESET = 64'h0;

typedef struct packed {
    logic [29:0] reserved0;  // RSVD
    logic  [7:0] AGE_COUNTER;  // RW
    logic [11:0] GROUP_IDX;  // RW
    logic [13:0] NEIGHBOR_IDX;  // RW
} NH_ROUTES_t;

localparam NH_ROUTES_REG_STRIDE = 48'h8;
localparam NH_ROUTES_REG_ENTRIES = 16384;
localparam NH_ROUTES_CR_ADDR = 48'h80000;
localparam NH_ROUTES_SIZE = 64;
localparam NH_ROUTES_AGE_COUNTER_LO = 26;
localparam NH_ROUTES_AGE_COUNTER_HI = 33;
localparam NH_ROUTES_AGE_COUNTER_RESET = 8'h0;
localparam NH_ROUTES_GROUP_IDX_LO = 14;
localparam NH_ROUTES_GROUP_IDX_HI = 25;
localparam NH_ROUTES_GROUP_IDX_RESET = 12'h0;
localparam NH_ROUTES_NEIGHBOR_IDX_LO = 0;
localparam NH_ROUTES_NEIGHBOR_IDX_HI = 13;
localparam NH_ROUTES_NEIGHBOR_IDX_RESET = 14'h0;
localparam NH_ROUTES_USEMASK = 64'h3FFFFFFFF;
localparam NH_ROUTES_RO_MASK = 64'h0;
localparam NH_ROUTES_WO_MASK = 64'h0;
localparam NH_ROUTES_RESET = 64'h0;

typedef struct packed {
    logic  [7:0] WEIGHT_7;  // RW
    logic  [7:0] WEIGHT_6;  // RW
    logic  [7:0] WEIGHT_5;  // RW
    logic  [7:0] WEIGHT_4;  // RW
    logic  [7:0] WEIGHT_3;  // RW
    logic  [7:0] WEIGHT_2;  // RW
    logic  [7:0] WEIGHT_1;  // RW
    logic  [7:0] WEIGHT_0;  // RW
} NH_WEIGHTS_t;

localparam NH_WEIGHTS_REG_STRIDE = 48'h8;
localparam NH_WEIGHTS_REG_ENTRIES = 8;
localparam NH_WEIGHTS_REGFILE_STRIDE = 48'h40;
localparam NH_WEIGHTS_REGFILE_ENTRIES = 2048;
localparam NH_WEIGHTS_CR_ADDR = 48'hA0000;
localparam NH_WEIGHTS_SIZE = 64;
localparam NH_WEIGHTS_WEIGHT_7_LO = 56;
localparam NH_WEIGHTS_WEIGHT_7_HI = 63;
localparam NH_WEIGHTS_WEIGHT_7_RESET = 8'h0;
localparam NH_WEIGHTS_WEIGHT_6_LO = 48;
localparam NH_WEIGHTS_WEIGHT_6_HI = 55;
localparam NH_WEIGHTS_WEIGHT_6_RESET = 8'h0;
localparam NH_WEIGHTS_WEIGHT_5_LO = 40;
localparam NH_WEIGHTS_WEIGHT_5_HI = 47;
localparam NH_WEIGHTS_WEIGHT_5_RESET = 8'h0;
localparam NH_WEIGHTS_WEIGHT_4_LO = 32;
localparam NH_WEIGHTS_WEIGHT_4_HI = 39;
localparam NH_WEIGHTS_WEIGHT_4_RESET = 8'h0;
localparam NH_WEIGHTS_WEIGHT_3_LO = 24;
localparam NH_WEIGHTS_WEIGHT_3_HI = 31;
localparam NH_WEIGHTS_WEIGHT_3_RESET = 8'h0;
localparam NH_WEIGHTS_WEIGHT_2_LO = 16;
localparam NH_WEIGHTS_WEIGHT_2_HI = 23;
localparam NH_WEIGHTS_WEIGHT_2_RESET = 8'h0;
localparam NH_WEIGHTS_WEIGHT_1_LO = 8;
localparam NH_WEIGHTS_WEIGHT_1_HI = 15;
localparam NH_WEIGHTS_WEIGHT_1_RESET = 8'h0;
localparam NH_WEIGHTS_WEIGHT_0_LO = 0;
localparam NH_WEIGHTS_WEIGHT_0_HI = 7;
localparam NH_WEIGHTS_WEIGHT_0_RESET = 8'h0;
localparam NH_WEIGHTS_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam NH_WEIGHTS_RO_MASK = 64'h0;
localparam NH_WEIGHTS_WO_MASK = 64'h0;
localparam NH_WEIGHTS_RESET = 64'h0;

typedef struct packed {
    logic [44:0] reserved0;  // RSVD
    logic  [0:0] TRAP_IGMP;  // RW
    logic  [0:0] REFLECT;  // RW
    logic [16:0] MEMBERSHIP;  // RW
} INGRESS_VID_TABLE_t;

localparam INGRESS_VID_TABLE_REG_STRIDE = 48'h8;
localparam INGRESS_VID_TABLE_REG_ENTRIES = 4096;
localparam INGRESS_VID_TABLE_CR_ADDR = 48'hC0000;
localparam INGRESS_VID_TABLE_SIZE = 64;
localparam INGRESS_VID_TABLE_TRAP_IGMP_LO = 18;
localparam INGRESS_VID_TABLE_TRAP_IGMP_HI = 18;
localparam INGRESS_VID_TABLE_TRAP_IGMP_RESET = 1'h0;
localparam INGRESS_VID_TABLE_REFLECT_LO = 17;
localparam INGRESS_VID_TABLE_REFLECT_HI = 17;
localparam INGRESS_VID_TABLE_REFLECT_RESET = 1'h0;
localparam INGRESS_VID_TABLE_MEMBERSHIP_LO = 0;
localparam INGRESS_VID_TABLE_MEMBERSHIP_HI = 16;
localparam INGRESS_VID_TABLE_MEMBERSHIP_RESET = 17'h0;
localparam INGRESS_VID_TABLE_USEMASK = 64'h7FFFF;
localparam INGRESS_VID_TABLE_RO_MASK = 64'h0;
localparam INGRESS_VID_TABLE_WO_MASK = 64'h0;
localparam INGRESS_VID_TABLE_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [15:0] BROADCAST_GLORT;  // RW
    logic [15:0] FLOOD_MULTICAST_GLORT;  // RW
    logic [15:0] FLOOD_UNICAST_GLORT;  // RW
} FLOOD_GLORT_TABLE_t;

localparam FLOOD_GLORT_TABLE_REG_STRIDE = 48'h8;
localparam FLOOD_GLORT_TABLE_REG_ENTRIES = 256;
localparam FLOOD_GLORT_TABLE_CR_ADDR = 48'hC8000;
localparam FLOOD_GLORT_TABLE_SIZE = 64;
localparam FLOOD_GLORT_TABLE_BROADCAST_GLORT_LO = 32;
localparam FLOOD_GLORT_TABLE_BROADCAST_GLORT_HI = 47;
localparam FLOOD_GLORT_TABLE_BROADCAST_GLORT_RESET = 16'h0;
localparam FLOOD_GLORT_TABLE_FLOOD_MULTICAST_GLORT_LO = 16;
localparam FLOOD_GLORT_TABLE_FLOOD_MULTICAST_GLORT_HI = 31;
localparam FLOOD_GLORT_TABLE_FLOOD_MULTICAST_GLORT_RESET = 16'h0;
localparam FLOOD_GLORT_TABLE_FLOOD_UNICAST_GLORT_LO = 0;
localparam FLOOD_GLORT_TABLE_FLOOD_UNICAST_GLORT_HI = 15;
localparam FLOOD_GLORT_TABLE_FLOOD_UNICAST_GLORT_RESET = 16'h0;
localparam FLOOD_GLORT_TABLE_USEMASK = 64'hFFFFFFFFFFFF;
localparam FLOOD_GLORT_TABLE_RO_MASK = 64'h0;
localparam FLOOD_GLORT_TABLE_WO_MASK = 64'h0;
localparam FLOOD_GLORT_TABLE_RESET = 64'h0;

typedef struct packed {
    logic [63:0] USED;  // RW/1C/V
} NH_USED_t;

localparam NH_USED_REG_STRIDE = 48'h8;
localparam NH_USED_REG_ENTRIES = 256;
localparam NH_USED_CR_ADDR = 48'hC8800;
localparam NH_USED_SIZE = 64;
localparam NH_USED_USED_LO = 0;
localparam NH_USED_USED_HI = 63;
localparam NH_USED_USED_RESET = 64'h0;
localparam NH_USED_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam NH_USED_RO_MASK = 64'h0;
localparam NH_USED_WO_MASK = 64'h0;
localparam NH_USED_RESET = 64'h0;

typedef struct packed {
    logic [63:0] BYTES;  // RW
} NH_PATH_CTRS_t;

localparam NH_PATH_CTRS_REG_STRIDE = 48'h8;
localparam NH_PATH_CTRS_REG_ENTRIES = 16384;
localparam NH_PATH_CTRS_CR_ADDR = 48'hE0000;
localparam NH_PATH_CTRS_SIZE = 64;
localparam NH_PATH_CTRS_BYTES_LO = 0;
localparam NH_PATH_CTRS_BYTES_HI = 63;
localparam NH_PATH_CTRS_BYTES_RESET = 64'h0;
localparam NH_PATH_CTRS_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam NH_PATH_CTRS_RO_MASK = 64'h0;
localparam NH_PATH_CTRS_WO_MASK = 64'h0;
localparam NH_PATH_CTRS_RESET = 64'h0;

typedef struct packed {
    logic [15:0] MIN_3;  // RW
    logic [15:0] MIN_2;  // RW
    logic [15:0] MIN_1;  // RW
    logic [15:0] MIN_0;  // RW
} NH_GROUP_MIN_t;

localparam NH_GROUP_MIN_REG_STRIDE = 48'h8;
localparam NH_GROUP_MIN_REG_ENTRIES = 512;
localparam NH_GROUP_MIN_CR_ADDR = 48'h100000;
localparam NH_GROUP_MIN_SIZE = 64;
localparam NH_GROUP_MIN_MIN_3_LO = 48;
localparam NH_GROUP_MIN_MIN_3_HI = 63;
localparam NH_GROUP_MIN_MIN_3_RESET = 16'h0;
localparam NH_GROUP_MIN_MIN_2_LO = 32;
localparam NH_GROUP_MIN_MIN_2_HI = 47;
localparam NH_GROUP_MIN_MIN_2_RESET = 16'h0;
localparam NH_GROUP_MIN_MIN_1_LO = 16;
localparam NH_GROUP_MIN_MIN_1_HI = 31;
localparam NH_GROUP_MIN_MIN_1_RESET = 16'h0;
localparam NH_GROUP_MIN_MIN_0_LO = 0;
localparam NH_GROUP_MIN_MIN_0_HI = 15;
localparam NH_GROUP_MIN_MIN_0_RESET = 16'h0;
localparam NH_GROUP_MIN_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam NH_GROUP_MIN_RO_MASK = 64'h0;
localparam NH_GROUP_MIN_WO_MASK = 64'h0;
localparam NH_GROUP_MIN_RESET = 64'h0;

typedef struct packed {
    logic [49:0] reserved0;  // RSVD
    logic [13:0] MTU;  // RW
} MTU_TABLE_t;

localparam MTU_TABLE_REG_STRIDE = 48'h8;
localparam MTU_TABLE_REG_ENTRIES = 8;
localparam MTU_TABLE_CR_ADDR = 48'h101000;
localparam MTU_TABLE_SIZE = 64;
localparam MTU_TABLE_MTU_LO = 0;
localparam MTU_TABLE_MTU_HI = 13;
localparam MTU_TABLE_MTU_RESET = 14'h0;
localparam MTU_TABLE_USEMASK = 64'h3FFF;
localparam MTU_TABLE_RO_MASK = 64'h0;
localparam MTU_TABLE_WO_MASK = 64'h0;
localparam MTU_TABLE_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_NH_CONFIG_t;

typedef logic [7:0] we_NH_STATUS_t;

typedef logic [7:0] we_NH_NEIGHBORS_0_t;

typedef logic [7:0] we_NH_NEIGHBORS_1_t;

typedef logic [7:0] we_NH_GROUPS_0_t;

typedef logic [7:0] we_NH_GROUPS_1_t;

typedef logic [7:0] we_NH_ROUTES_t;

typedef logic [7:0] we_NH_WEIGHTS_t;

typedef logic [7:0] we_INGRESS_VID_TABLE_t;

typedef logic [7:0] we_FLOOD_GLORT_TABLE_t;

typedef logic [7:0] we_NH_USED_t;

typedef logic [7:0] we_NH_PATH_CTRS_t;

typedef logic [7:0] we_NH_GROUP_MIN_t;

typedef logic [7:0] we_MTU_TABLE_t;

typedef struct packed {
    we_NH_CONFIG_t NH_CONFIG;
    we_NH_STATUS_t NH_STATUS;
    we_NH_NEIGHBORS_0_t NH_NEIGHBORS_0;
    we_NH_NEIGHBORS_1_t NH_NEIGHBORS_1;
    we_NH_GROUPS_0_t NH_GROUPS_0;
    we_NH_GROUPS_1_t NH_GROUPS_1;
    we_NH_ROUTES_t NH_ROUTES;
    we_NH_WEIGHTS_t NH_WEIGHTS;
    we_INGRESS_VID_TABLE_t INGRESS_VID_TABLE;
    we_FLOOD_GLORT_TABLE_t FLOOD_GLORT_TABLE;
    we_NH_USED_t NH_USED;
    we_NH_PATH_CTRS_t NH_PATH_CTRS;
    we_NH_GROUP_MIN_t NH_GROUP_MIN;
    we_MTU_TABLE_t MTU_TABLE;
} mby_ppe_nexthop_map_handcoded_t;

typedef logic [7:0] re_NH_CONFIG_t;

typedef logic [7:0] re_NH_STATUS_t;

typedef logic [7:0] re_NH_NEIGHBORS_0_t;

typedef logic [7:0] re_NH_NEIGHBORS_1_t;

typedef logic [7:0] re_NH_GROUPS_0_t;

typedef logic [7:0] re_NH_GROUPS_1_t;

typedef logic [7:0] re_NH_ROUTES_t;

typedef logic [7:0] re_NH_WEIGHTS_t;

typedef logic [7:0] re_INGRESS_VID_TABLE_t;

typedef logic [7:0] re_FLOOD_GLORT_TABLE_t;

typedef logic [7:0] re_NH_USED_t;

typedef logic [7:0] re_NH_PATH_CTRS_t;

typedef logic [7:0] re_NH_GROUP_MIN_t;

typedef logic [7:0] re_MTU_TABLE_t;

typedef struct packed {
    re_NH_CONFIG_t NH_CONFIG;
    re_NH_STATUS_t NH_STATUS;
    re_NH_NEIGHBORS_0_t NH_NEIGHBORS_0;
    re_NH_NEIGHBORS_1_t NH_NEIGHBORS_1;
    re_NH_GROUPS_0_t NH_GROUPS_0;
    re_NH_GROUPS_1_t NH_GROUPS_1;
    re_NH_ROUTES_t NH_ROUTES;
    re_NH_WEIGHTS_t NH_WEIGHTS;
    re_INGRESS_VID_TABLE_t INGRESS_VID_TABLE;
    re_FLOOD_GLORT_TABLE_t FLOOD_GLORT_TABLE;
    re_NH_USED_t NH_USED;
    re_NH_PATH_CTRS_t NH_PATH_CTRS;
    re_NH_GROUP_MIN_t NH_GROUP_MIN;
    re_MTU_TABLE_t MTU_TABLE;
} mby_ppe_nexthop_map_hc_re_t;

typedef logic handcode_rvalid_NH_CONFIG_t;

typedef logic handcode_rvalid_NH_STATUS_t;

typedef logic handcode_rvalid_NH_NEIGHBORS_0_t;

typedef logic handcode_rvalid_NH_NEIGHBORS_1_t;

typedef logic handcode_rvalid_NH_GROUPS_0_t;

typedef logic handcode_rvalid_NH_GROUPS_1_t;

typedef logic handcode_rvalid_NH_ROUTES_t;

typedef logic handcode_rvalid_NH_WEIGHTS_t;

typedef logic handcode_rvalid_INGRESS_VID_TABLE_t;

typedef logic handcode_rvalid_FLOOD_GLORT_TABLE_t;

typedef logic handcode_rvalid_NH_USED_t;

typedef logic handcode_rvalid_NH_PATH_CTRS_t;

typedef logic handcode_rvalid_NH_GROUP_MIN_t;

typedef logic handcode_rvalid_MTU_TABLE_t;

typedef struct packed {
    handcode_rvalid_NH_CONFIG_t NH_CONFIG;
    handcode_rvalid_NH_STATUS_t NH_STATUS;
    handcode_rvalid_NH_NEIGHBORS_0_t NH_NEIGHBORS_0;
    handcode_rvalid_NH_NEIGHBORS_1_t NH_NEIGHBORS_1;
    handcode_rvalid_NH_GROUPS_0_t NH_GROUPS_0;
    handcode_rvalid_NH_GROUPS_1_t NH_GROUPS_1;
    handcode_rvalid_NH_ROUTES_t NH_ROUTES;
    handcode_rvalid_NH_WEIGHTS_t NH_WEIGHTS;
    handcode_rvalid_INGRESS_VID_TABLE_t INGRESS_VID_TABLE;
    handcode_rvalid_FLOOD_GLORT_TABLE_t FLOOD_GLORT_TABLE;
    handcode_rvalid_NH_USED_t NH_USED;
    handcode_rvalid_NH_PATH_CTRS_t NH_PATH_CTRS;
    handcode_rvalid_NH_GROUP_MIN_t NH_GROUP_MIN;
    handcode_rvalid_MTU_TABLE_t MTU_TABLE;
} mby_ppe_nexthop_map_hc_rvalid_t;

typedef logic handcode_wvalid_NH_CONFIG_t;

typedef logic handcode_wvalid_NH_STATUS_t;

typedef logic handcode_wvalid_NH_NEIGHBORS_0_t;

typedef logic handcode_wvalid_NH_NEIGHBORS_1_t;

typedef logic handcode_wvalid_NH_GROUPS_0_t;

typedef logic handcode_wvalid_NH_GROUPS_1_t;

typedef logic handcode_wvalid_NH_ROUTES_t;

typedef logic handcode_wvalid_NH_WEIGHTS_t;

typedef logic handcode_wvalid_INGRESS_VID_TABLE_t;

typedef logic handcode_wvalid_FLOOD_GLORT_TABLE_t;

typedef logic handcode_wvalid_NH_USED_t;

typedef logic handcode_wvalid_NH_PATH_CTRS_t;

typedef logic handcode_wvalid_NH_GROUP_MIN_t;

typedef logic handcode_wvalid_MTU_TABLE_t;

typedef struct packed {
    handcode_wvalid_NH_CONFIG_t NH_CONFIG;
    handcode_wvalid_NH_STATUS_t NH_STATUS;
    handcode_wvalid_NH_NEIGHBORS_0_t NH_NEIGHBORS_0;
    handcode_wvalid_NH_NEIGHBORS_1_t NH_NEIGHBORS_1;
    handcode_wvalid_NH_GROUPS_0_t NH_GROUPS_0;
    handcode_wvalid_NH_GROUPS_1_t NH_GROUPS_1;
    handcode_wvalid_NH_ROUTES_t NH_ROUTES;
    handcode_wvalid_NH_WEIGHTS_t NH_WEIGHTS;
    handcode_wvalid_INGRESS_VID_TABLE_t INGRESS_VID_TABLE;
    handcode_wvalid_FLOOD_GLORT_TABLE_t FLOOD_GLORT_TABLE;
    handcode_wvalid_NH_USED_t NH_USED;
    handcode_wvalid_NH_PATH_CTRS_t NH_PATH_CTRS;
    handcode_wvalid_NH_GROUP_MIN_t NH_GROUP_MIN;
    handcode_wvalid_MTU_TABLE_t MTU_TABLE;
} mby_ppe_nexthop_map_hc_wvalid_t;

typedef logic handcode_error_NH_CONFIG_t;

typedef logic handcode_error_NH_STATUS_t;

typedef logic handcode_error_NH_NEIGHBORS_0_t;

typedef logic handcode_error_NH_NEIGHBORS_1_t;

typedef logic handcode_error_NH_GROUPS_0_t;

typedef logic handcode_error_NH_GROUPS_1_t;

typedef logic handcode_error_NH_ROUTES_t;

typedef logic handcode_error_NH_WEIGHTS_t;

typedef logic handcode_error_INGRESS_VID_TABLE_t;

typedef logic handcode_error_FLOOD_GLORT_TABLE_t;

typedef logic handcode_error_NH_USED_t;

typedef logic handcode_error_NH_PATH_CTRS_t;

typedef logic handcode_error_NH_GROUP_MIN_t;

typedef logic handcode_error_MTU_TABLE_t;

typedef struct packed {
    handcode_error_NH_CONFIG_t NH_CONFIG;
    handcode_error_NH_STATUS_t NH_STATUS;
    handcode_error_NH_NEIGHBORS_0_t NH_NEIGHBORS_0;
    handcode_error_NH_NEIGHBORS_1_t NH_NEIGHBORS_1;
    handcode_error_NH_GROUPS_0_t NH_GROUPS_0;
    handcode_error_NH_GROUPS_1_t NH_GROUPS_1;
    handcode_error_NH_ROUTES_t NH_ROUTES;
    handcode_error_NH_WEIGHTS_t NH_WEIGHTS;
    handcode_error_INGRESS_VID_TABLE_t INGRESS_VID_TABLE;
    handcode_error_FLOOD_GLORT_TABLE_t FLOOD_GLORT_TABLE;
    handcode_error_NH_USED_t NH_USED;
    handcode_error_NH_PATH_CTRS_t NH_PATH_CTRS;
    handcode_error_NH_GROUP_MIN_t NH_GROUP_MIN;
    handcode_error_MTU_TABLE_t MTU_TABLE;
} mby_ppe_nexthop_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    NH_CONFIG_t NH_CONFIG;
    NH_STATUS_t NH_STATUS;
    NH_NEIGHBORS_0_t NH_NEIGHBORS_0;
    NH_NEIGHBORS_1_t NH_NEIGHBORS_1;
    NH_GROUPS_0_t NH_GROUPS_0;
    NH_GROUPS_1_t NH_GROUPS_1;
    NH_ROUTES_t NH_ROUTES;
    NH_WEIGHTS_t NH_WEIGHTS;
    INGRESS_VID_TABLE_t INGRESS_VID_TABLE;
    FLOOD_GLORT_TABLE_t FLOOD_GLORT_TABLE;
    NH_USED_t NH_USED;
    NH_PATH_CTRS_t NH_PATH_CTRS;
    NH_GROUP_MIN_t NH_GROUP_MIN;
    MTU_TABLE_t MTU_TABLE;
} mby_ppe_nexthop_map_hc_reg_read_t;

typedef struct packed {
    NH_CONFIG_t NH_CONFIG;
    NH_STATUS_t NH_STATUS;
    NH_NEIGHBORS_0_t NH_NEIGHBORS_0;
    NH_NEIGHBORS_1_t NH_NEIGHBORS_1;
    NH_GROUPS_0_t NH_GROUPS_0;
    NH_GROUPS_1_t NH_GROUPS_1;
    NH_ROUTES_t NH_ROUTES;
    NH_WEIGHTS_t NH_WEIGHTS;
    INGRESS_VID_TABLE_t INGRESS_VID_TABLE;
    FLOOD_GLORT_TABLE_t FLOOD_GLORT_TABLE;
    NH_USED_t NH_USED;
    NH_PATH_CTRS_t NH_PATH_CTRS;
    NH_GROUP_MIN_t NH_GROUP_MIN;
    MTU_TABLE_t MTU_TABLE;
} mby_ppe_nexthop_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_nexthop_map_pkg

`endif // MBY_PPE_NEXTHOP_MAP_PKG_VH
