magic
tech scmos
timestamp 970029517
<< ndiffusion >>
rect -35 44 -31 47
rect -16 37 -8 38
rect -35 33 -31 36
rect -16 33 -8 34
<< pdiffusion >>
rect 29 44 33 47
rect 8 37 16 38
rect 8 33 16 34
rect 29 33 33 40
rect 66 46 74 47
rect 66 42 74 43
<< ntransistor >>
rect -35 36 -31 44
rect -16 34 -8 37
<< ptransistor >>
rect 29 40 33 44
rect 8 34 16 37
rect 66 43 74 46
<< polysilicon >>
rect -28 44 -26 45
rect -39 36 -35 44
rect -31 42 -26 44
rect -31 36 -25 42
rect -2 37 2 46
rect 25 40 29 44
rect 33 40 37 44
rect -20 34 -16 37
rect -8 34 8 37
rect 16 34 20 37
rect 62 43 66 46
rect 74 43 78 46
<< ndcontact >>
rect -38 47 -30 55
rect -16 38 -8 46
rect -35 25 -27 33
rect -16 25 -8 33
<< pdcontact >>
rect 25 47 33 55
rect 66 47 74 55
rect 8 38 16 46
rect 8 25 16 33
rect 25 25 33 33
rect 66 34 74 42
<< psubstratepcontact >>
rect -52 29 -44 37
<< nsubstratencontact >>
rect 42 27 50 35
<< polycontact >>
rect -26 42 -18 50
rect -4 46 4 54
rect 37 39 45 47
rect 54 38 62 46
<< metal1 >>
rect -38 47 -30 49
rect -26 46 -18 50
rect -4 46 4 49
rect 25 47 33 49
rect 66 47 74 49
rect -26 42 -8 46
rect 8 43 16 46
rect 37 43 45 47
rect 8 42 45 43
rect -16 39 45 42
rect 54 43 62 46
rect -16 38 16 39
rect -52 33 -44 37
rect 42 33 50 35
rect 66 33 74 42
rect -52 31 -8 33
rect 8 31 74 33
rect -52 29 -19 31
rect -35 25 -19 29
rect 21 25 74 31
<< m2contact >>
rect -38 49 -30 55
rect -4 49 4 55
rect 25 49 33 55
rect 66 49 74 55
rect 54 37 62 43
rect -19 25 -3 31
rect 3 25 21 31
<< metal2 >>
rect -38 49 74 55
rect 0 37 62 43
<< m3contact >>
rect -21 25 -3 31
rect 3 25 21 31
<< metal3 >>
rect -21 22 -3 58
rect 3 22 21 58
<< labels >>
rlabel ndcontact -12 29 -12 29 1 GND!
rlabel pdcontact 12 29 12 29 1 Vdd!
rlabel metal2 0 37 0 43 3 a
rlabel metal2 0 49 0 55 1 x
rlabel metal1 -31 29 -31 29 1 GND!
rlabel metal1 -48 33 -48 33 3 GND!
rlabel pdcontact 29 29 29 29 1 Vdd!
rlabel metal1 46 31 46 31 1 Vdd!
rlabel metal1 70 38 70 38 1 Vdd!
rlabel polysilicon 65 44 65 44 1 a
rlabel space 74 25 79 55 3 ^p
rlabel metal2 -34 52 -34 52 1 x
rlabel metal2 29 52 29 52 1 x
rlabel metal2 70 52 70 52 1 x
rlabel metal2 58 40 58 40 1 a
<< end >>
