///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cm_usage_map.sv                                    
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_cm_usage_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_FF
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_FF

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_RSTD


module rtlgen_mby_ppe_cm_usage_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_cm_usage_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_PH2_FF
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CM_USAGE_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_cm_usage_map ( //lintra s-2096
    // Clocks
    gated_clk,
    rtl_clk,

    // Resets
    rst_n,


    // Register Inputs
    load_CM_GLOBAL_USAGE_MAX,

    new_CM_GLOBAL_USAGE,
    new_CM_GLOBAL_USAGE_MAX,

    handcode_reg_rdata_CM_AQM_DCTCP_CFG,
    handcode_reg_rdata_CM_AQM_EWMA_CFG,
    handcode_reg_rdata_CM_FORCE_PAUSE_CFG,
    handcode_reg_rdata_CM_MCAST_EPOCH_USAGE,
    handcode_reg_rdata_CM_PAUSE_GEN_STATE,
    handcode_reg_rdata_CM_PAUSE_PHYS_PORT_CFG,
    handcode_reg_rdata_CM_RX_SMP_HOG_WM,
    handcode_reg_rdata_CM_RX_SMP_PAUSE_WM,
    handcode_reg_rdata_CM_RX_SMP_PRIVATE_WM,
    handcode_reg_rdata_CM_RX_SMP_USAGE,
    handcode_reg_rdata_CM_RX_SMP_USAGE_MAX,
    handcode_reg_rdata_CM_RX_SMP_USAGE_MAX_CTRL,
    handcode_reg_rdata_CM_SHARED_SMP_PAUSE_CFG,
    handcode_reg_rdata_CM_SHARED_SMP_PAUSE_WM,
    handcode_reg_rdata_CM_SHARED_SMP_USAGE,
    handcode_reg_rdata_CM_SHARED_WM,
    handcode_reg_rdata_CM_SMP_USAGE,
    handcode_reg_rdata_CM_SOFTDROP_WM,
    handcode_reg_rdata_CM_TX_EWMA,
    handcode_reg_rdata_CM_TX_TC_HOG_WM,
    handcode_reg_rdata_CM_TX_TC_PRIVATE_WM,
    handcode_reg_rdata_CM_TX_TC_USAGE,

    handcode_rvalid_CM_AQM_DCTCP_CFG,
    handcode_rvalid_CM_AQM_EWMA_CFG,
    handcode_rvalid_CM_FORCE_PAUSE_CFG,
    handcode_rvalid_CM_MCAST_EPOCH_USAGE,
    handcode_rvalid_CM_PAUSE_GEN_STATE,
    handcode_rvalid_CM_PAUSE_PHYS_PORT_CFG,
    handcode_rvalid_CM_RX_SMP_HOG_WM,
    handcode_rvalid_CM_RX_SMP_PAUSE_WM,
    handcode_rvalid_CM_RX_SMP_PRIVATE_WM,
    handcode_rvalid_CM_RX_SMP_USAGE,
    handcode_rvalid_CM_RX_SMP_USAGE_MAX,
    handcode_rvalid_CM_RX_SMP_USAGE_MAX_CTRL,
    handcode_rvalid_CM_SHARED_SMP_PAUSE_CFG,
    handcode_rvalid_CM_SHARED_SMP_PAUSE_WM,
    handcode_rvalid_CM_SHARED_SMP_USAGE,
    handcode_rvalid_CM_SHARED_WM,
    handcode_rvalid_CM_SMP_USAGE,
    handcode_rvalid_CM_SOFTDROP_WM,
    handcode_rvalid_CM_TX_EWMA,
    handcode_rvalid_CM_TX_TC_HOG_WM,
    handcode_rvalid_CM_TX_TC_PRIVATE_WM,
    handcode_rvalid_CM_TX_TC_USAGE,

    handcode_wvalid_CM_AQM_DCTCP_CFG,
    handcode_wvalid_CM_AQM_EWMA_CFG,
    handcode_wvalid_CM_FORCE_PAUSE_CFG,
    handcode_wvalid_CM_MCAST_EPOCH_USAGE,
    handcode_wvalid_CM_PAUSE_GEN_STATE,
    handcode_wvalid_CM_PAUSE_PHYS_PORT_CFG,
    handcode_wvalid_CM_RX_SMP_HOG_WM,
    handcode_wvalid_CM_RX_SMP_PAUSE_WM,
    handcode_wvalid_CM_RX_SMP_PRIVATE_WM,
    handcode_wvalid_CM_RX_SMP_USAGE,
    handcode_wvalid_CM_RX_SMP_USAGE_MAX,
    handcode_wvalid_CM_RX_SMP_USAGE_MAX_CTRL,
    handcode_wvalid_CM_SHARED_SMP_PAUSE_CFG,
    handcode_wvalid_CM_SHARED_SMP_PAUSE_WM,
    handcode_wvalid_CM_SHARED_SMP_USAGE,
    handcode_wvalid_CM_SHARED_WM,
    handcode_wvalid_CM_SMP_USAGE,
    handcode_wvalid_CM_SOFTDROP_WM,
    handcode_wvalid_CM_TX_EWMA,
    handcode_wvalid_CM_TX_TC_HOG_WM,
    handcode_wvalid_CM_TX_TC_PRIVATE_WM,
    handcode_wvalid_CM_TX_TC_USAGE,

    handcode_error_CM_AQM_DCTCP_CFG,
    handcode_error_CM_AQM_EWMA_CFG,
    handcode_error_CM_FORCE_PAUSE_CFG,
    handcode_error_CM_MCAST_EPOCH_USAGE,
    handcode_error_CM_PAUSE_GEN_STATE,
    handcode_error_CM_PAUSE_PHYS_PORT_CFG,
    handcode_error_CM_RX_SMP_HOG_WM,
    handcode_error_CM_RX_SMP_PAUSE_WM,
    handcode_error_CM_RX_SMP_PRIVATE_WM,
    handcode_error_CM_RX_SMP_USAGE,
    handcode_error_CM_RX_SMP_USAGE_MAX,
    handcode_error_CM_RX_SMP_USAGE_MAX_CTRL,
    handcode_error_CM_SHARED_SMP_PAUSE_CFG,
    handcode_error_CM_SHARED_SMP_PAUSE_WM,
    handcode_error_CM_SHARED_SMP_USAGE,
    handcode_error_CM_SHARED_WM,
    handcode_error_CM_SMP_USAGE,
    handcode_error_CM_SOFTDROP_WM,
    handcode_error_CM_TX_EWMA,
    handcode_error_CM_TX_TC_HOG_WM,
    handcode_error_CM_TX_TC_PRIVATE_WM,
    handcode_error_CM_TX_TC_USAGE,


    // Register Outputs
    CM_GLOBAL_CFG,
    CM_GLOBAL_USAGE,
    CM_GLOBAL_USAGE_MAX,
    CM_GLOBAL_WM,
    CM_SWEEPER_TC_TO_SMP,


    // Register signals for HandCoded registers
    handcode_reg_wdata_CM_AQM_DCTCP_CFG,
    handcode_reg_wdata_CM_AQM_EWMA_CFG,
    handcode_reg_wdata_CM_FORCE_PAUSE_CFG,
    handcode_reg_wdata_CM_MCAST_EPOCH_USAGE,
    handcode_reg_wdata_CM_PAUSE_GEN_STATE,
    handcode_reg_wdata_CM_PAUSE_PHYS_PORT_CFG,
    handcode_reg_wdata_CM_RX_SMP_HOG_WM,
    handcode_reg_wdata_CM_RX_SMP_PAUSE_WM,
    handcode_reg_wdata_CM_RX_SMP_PRIVATE_WM,
    handcode_reg_wdata_CM_RX_SMP_USAGE,
    handcode_reg_wdata_CM_RX_SMP_USAGE_MAX,
    handcode_reg_wdata_CM_RX_SMP_USAGE_MAX_CTRL,
    handcode_reg_wdata_CM_SHARED_SMP_PAUSE_CFG,
    handcode_reg_wdata_CM_SHARED_SMP_PAUSE_WM,
    handcode_reg_wdata_CM_SHARED_SMP_USAGE,
    handcode_reg_wdata_CM_SHARED_WM,
    handcode_reg_wdata_CM_SMP_USAGE,
    handcode_reg_wdata_CM_SOFTDROP_WM,
    handcode_reg_wdata_CM_TX_EWMA,
    handcode_reg_wdata_CM_TX_TC_HOG_WM,
    handcode_reg_wdata_CM_TX_TC_PRIVATE_WM,
    handcode_reg_wdata_CM_TX_TC_USAGE,

    we_CM_AQM_DCTCP_CFG,
    we_CM_AQM_EWMA_CFG,
    we_CM_FORCE_PAUSE_CFG,
    we_CM_MCAST_EPOCH_USAGE,
    we_CM_PAUSE_GEN_STATE,
    we_CM_PAUSE_PHYS_PORT_CFG,
    we_CM_RX_SMP_HOG_WM,
    we_CM_RX_SMP_PAUSE_WM,
    we_CM_RX_SMP_PRIVATE_WM,
    we_CM_RX_SMP_USAGE,
    we_CM_RX_SMP_USAGE_MAX,
    we_CM_RX_SMP_USAGE_MAX_CTRL,
    we_CM_SHARED_SMP_PAUSE_CFG,
    we_CM_SHARED_SMP_PAUSE_WM,
    we_CM_SHARED_SMP_USAGE,
    we_CM_SHARED_WM,
    we_CM_SMP_USAGE,
    we_CM_SOFTDROP_WM,
    we_CM_TX_EWMA,
    we_CM_TX_TC_HOG_WM,
    we_CM_TX_TC_PRIVATE_WM,
    we_CM_TX_TC_USAGE,

    re_CM_AQM_DCTCP_CFG,
    re_CM_AQM_EWMA_CFG,
    re_CM_FORCE_PAUSE_CFG,
    re_CM_MCAST_EPOCH_USAGE,
    re_CM_PAUSE_GEN_STATE,
    re_CM_PAUSE_PHYS_PORT_CFG,
    re_CM_RX_SMP_HOG_WM,
    re_CM_RX_SMP_PAUSE_WM,
    re_CM_RX_SMP_PRIVATE_WM,
    re_CM_RX_SMP_USAGE,
    re_CM_RX_SMP_USAGE_MAX,
    re_CM_RX_SMP_USAGE_MAX_CTRL,
    re_CM_SHARED_SMP_PAUSE_CFG,
    re_CM_SHARED_SMP_PAUSE_WM,
    re_CM_SHARED_SMP_USAGE,
    re_CM_SHARED_WM,
    re_CM_SMP_USAGE,
    re_CM_SOFTDROP_WM,
    re_CM_TX_EWMA,
    re_CM_TX_TC_HOG_WM,
    re_CM_TX_TC_PRIVATE_WM,
    re_CM_TX_TC_USAGE,




    // Config Access
    req,
    ack
    

);

import mby_ppe_cm_usage_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:0] MBY_PPE_CM_USAGE_MAP_OFFSET = {MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] CM_USAGE_SB_BAR = 3'b0;
parameter [7:0] CM_USAGE_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
localparam [MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_GLOBAL_WM_DECODE_ADDR = CM_GLOBAL_WM_CR_ADDR[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_USAGE_MAP_OFFSET[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_GLOBAL_CFG_DECODE_ADDR = CM_GLOBAL_CFG_CR_ADDR[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_USAGE_MAP_OFFSET[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_SWEEPER_TC_TO_SMP_DECODE_ADDR = CM_SWEEPER_TC_TO_SMP_CR_ADDR[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_USAGE_MAP_OFFSET[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_GLOBAL_USAGE_DECODE_ADDR = CM_GLOBAL_USAGE_CR_ADDR[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_USAGE_MAP_OFFSET[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_GLOBAL_USAGE_MAX_DECODE_ADDR = CM_GLOBAL_USAGE_MAX_CR_ADDR[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_USAGE_MAP_OFFSET[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];

    // Clocks
input logic  gated_clk;
input logic  rtl_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input load_CM_GLOBAL_USAGE_MAX_t  load_CM_GLOBAL_USAGE_MAX;

input new_CM_GLOBAL_USAGE_t  new_CM_GLOBAL_USAGE;
input new_CM_GLOBAL_USAGE_MAX_t  new_CM_GLOBAL_USAGE_MAX;

input CM_AQM_DCTCP_CFG_t  handcode_reg_rdata_CM_AQM_DCTCP_CFG;
input CM_AQM_EWMA_CFG_t  handcode_reg_rdata_CM_AQM_EWMA_CFG;
input CM_FORCE_PAUSE_CFG_t  handcode_reg_rdata_CM_FORCE_PAUSE_CFG;
input CM_MCAST_EPOCH_USAGE_t  handcode_reg_rdata_CM_MCAST_EPOCH_USAGE;
input CM_PAUSE_GEN_STATE_t  handcode_reg_rdata_CM_PAUSE_GEN_STATE;
input CM_PAUSE_PHYS_PORT_CFG_t  handcode_reg_rdata_CM_PAUSE_PHYS_PORT_CFG;
input CM_RX_SMP_HOG_WM_t  handcode_reg_rdata_CM_RX_SMP_HOG_WM;
input CM_RX_SMP_PAUSE_WM_t  handcode_reg_rdata_CM_RX_SMP_PAUSE_WM;
input CM_RX_SMP_PRIVATE_WM_t  handcode_reg_rdata_CM_RX_SMP_PRIVATE_WM;
input CM_RX_SMP_USAGE_t  handcode_reg_rdata_CM_RX_SMP_USAGE;
input CM_RX_SMP_USAGE_MAX_t  handcode_reg_rdata_CM_RX_SMP_USAGE_MAX;
input CM_RX_SMP_USAGE_MAX_CTRL_t  handcode_reg_rdata_CM_RX_SMP_USAGE_MAX_CTRL;
input CM_SHARED_SMP_PAUSE_CFG_t  handcode_reg_rdata_CM_SHARED_SMP_PAUSE_CFG;
input CM_SHARED_SMP_PAUSE_WM_t  handcode_reg_rdata_CM_SHARED_SMP_PAUSE_WM;
input CM_SHARED_SMP_USAGE_t  handcode_reg_rdata_CM_SHARED_SMP_USAGE;
input CM_SHARED_WM_t  handcode_reg_rdata_CM_SHARED_WM;
input CM_SMP_USAGE_t  handcode_reg_rdata_CM_SMP_USAGE;
input CM_SOFTDROP_WM_t  handcode_reg_rdata_CM_SOFTDROP_WM;
input CM_TX_EWMA_t  handcode_reg_rdata_CM_TX_EWMA;
input CM_TX_TC_HOG_WM_t  handcode_reg_rdata_CM_TX_TC_HOG_WM;
input CM_TX_TC_PRIVATE_WM_t  handcode_reg_rdata_CM_TX_TC_PRIVATE_WM;
input CM_TX_TC_USAGE_t  handcode_reg_rdata_CM_TX_TC_USAGE;

input handcode_rvalid_CM_AQM_DCTCP_CFG_t  handcode_rvalid_CM_AQM_DCTCP_CFG;
input handcode_rvalid_CM_AQM_EWMA_CFG_t  handcode_rvalid_CM_AQM_EWMA_CFG;
input handcode_rvalid_CM_FORCE_PAUSE_CFG_t  handcode_rvalid_CM_FORCE_PAUSE_CFG;
input handcode_rvalid_CM_MCAST_EPOCH_USAGE_t  handcode_rvalid_CM_MCAST_EPOCH_USAGE;
input handcode_rvalid_CM_PAUSE_GEN_STATE_t  handcode_rvalid_CM_PAUSE_GEN_STATE;
input handcode_rvalid_CM_PAUSE_PHYS_PORT_CFG_t  handcode_rvalid_CM_PAUSE_PHYS_PORT_CFG;
input handcode_rvalid_CM_RX_SMP_HOG_WM_t  handcode_rvalid_CM_RX_SMP_HOG_WM;
input handcode_rvalid_CM_RX_SMP_PAUSE_WM_t  handcode_rvalid_CM_RX_SMP_PAUSE_WM;
input handcode_rvalid_CM_RX_SMP_PRIVATE_WM_t  handcode_rvalid_CM_RX_SMP_PRIVATE_WM;
input handcode_rvalid_CM_RX_SMP_USAGE_t  handcode_rvalid_CM_RX_SMP_USAGE;
input handcode_rvalid_CM_RX_SMP_USAGE_MAX_t  handcode_rvalid_CM_RX_SMP_USAGE_MAX;
input handcode_rvalid_CM_RX_SMP_USAGE_MAX_CTRL_t  handcode_rvalid_CM_RX_SMP_USAGE_MAX_CTRL;
input handcode_rvalid_CM_SHARED_SMP_PAUSE_CFG_t  handcode_rvalid_CM_SHARED_SMP_PAUSE_CFG;
input handcode_rvalid_CM_SHARED_SMP_PAUSE_WM_t  handcode_rvalid_CM_SHARED_SMP_PAUSE_WM;
input handcode_rvalid_CM_SHARED_SMP_USAGE_t  handcode_rvalid_CM_SHARED_SMP_USAGE;
input handcode_rvalid_CM_SHARED_WM_t  handcode_rvalid_CM_SHARED_WM;
input handcode_rvalid_CM_SMP_USAGE_t  handcode_rvalid_CM_SMP_USAGE;
input handcode_rvalid_CM_SOFTDROP_WM_t  handcode_rvalid_CM_SOFTDROP_WM;
input handcode_rvalid_CM_TX_EWMA_t  handcode_rvalid_CM_TX_EWMA;
input handcode_rvalid_CM_TX_TC_HOG_WM_t  handcode_rvalid_CM_TX_TC_HOG_WM;
input handcode_rvalid_CM_TX_TC_PRIVATE_WM_t  handcode_rvalid_CM_TX_TC_PRIVATE_WM;
input handcode_rvalid_CM_TX_TC_USAGE_t  handcode_rvalid_CM_TX_TC_USAGE;

input handcode_wvalid_CM_AQM_DCTCP_CFG_t  handcode_wvalid_CM_AQM_DCTCP_CFG;
input handcode_wvalid_CM_AQM_EWMA_CFG_t  handcode_wvalid_CM_AQM_EWMA_CFG;
input handcode_wvalid_CM_FORCE_PAUSE_CFG_t  handcode_wvalid_CM_FORCE_PAUSE_CFG;
input handcode_wvalid_CM_MCAST_EPOCH_USAGE_t  handcode_wvalid_CM_MCAST_EPOCH_USAGE;
input handcode_wvalid_CM_PAUSE_GEN_STATE_t  handcode_wvalid_CM_PAUSE_GEN_STATE;
input handcode_wvalid_CM_PAUSE_PHYS_PORT_CFG_t  handcode_wvalid_CM_PAUSE_PHYS_PORT_CFG;
input handcode_wvalid_CM_RX_SMP_HOG_WM_t  handcode_wvalid_CM_RX_SMP_HOG_WM;
input handcode_wvalid_CM_RX_SMP_PAUSE_WM_t  handcode_wvalid_CM_RX_SMP_PAUSE_WM;
input handcode_wvalid_CM_RX_SMP_PRIVATE_WM_t  handcode_wvalid_CM_RX_SMP_PRIVATE_WM;
input handcode_wvalid_CM_RX_SMP_USAGE_t  handcode_wvalid_CM_RX_SMP_USAGE;
input handcode_wvalid_CM_RX_SMP_USAGE_MAX_t  handcode_wvalid_CM_RX_SMP_USAGE_MAX;
input handcode_wvalid_CM_RX_SMP_USAGE_MAX_CTRL_t  handcode_wvalid_CM_RX_SMP_USAGE_MAX_CTRL;
input handcode_wvalid_CM_SHARED_SMP_PAUSE_CFG_t  handcode_wvalid_CM_SHARED_SMP_PAUSE_CFG;
input handcode_wvalid_CM_SHARED_SMP_PAUSE_WM_t  handcode_wvalid_CM_SHARED_SMP_PAUSE_WM;
input handcode_wvalid_CM_SHARED_SMP_USAGE_t  handcode_wvalid_CM_SHARED_SMP_USAGE;
input handcode_wvalid_CM_SHARED_WM_t  handcode_wvalid_CM_SHARED_WM;
input handcode_wvalid_CM_SMP_USAGE_t  handcode_wvalid_CM_SMP_USAGE;
input handcode_wvalid_CM_SOFTDROP_WM_t  handcode_wvalid_CM_SOFTDROP_WM;
input handcode_wvalid_CM_TX_EWMA_t  handcode_wvalid_CM_TX_EWMA;
input handcode_wvalid_CM_TX_TC_HOG_WM_t  handcode_wvalid_CM_TX_TC_HOG_WM;
input handcode_wvalid_CM_TX_TC_PRIVATE_WM_t  handcode_wvalid_CM_TX_TC_PRIVATE_WM;
input handcode_wvalid_CM_TX_TC_USAGE_t  handcode_wvalid_CM_TX_TC_USAGE;

input handcode_error_CM_AQM_DCTCP_CFG_t  handcode_error_CM_AQM_DCTCP_CFG;
input handcode_error_CM_AQM_EWMA_CFG_t  handcode_error_CM_AQM_EWMA_CFG;
input handcode_error_CM_FORCE_PAUSE_CFG_t  handcode_error_CM_FORCE_PAUSE_CFG;
input handcode_error_CM_MCAST_EPOCH_USAGE_t  handcode_error_CM_MCAST_EPOCH_USAGE;
input handcode_error_CM_PAUSE_GEN_STATE_t  handcode_error_CM_PAUSE_GEN_STATE;
input handcode_error_CM_PAUSE_PHYS_PORT_CFG_t  handcode_error_CM_PAUSE_PHYS_PORT_CFG;
input handcode_error_CM_RX_SMP_HOG_WM_t  handcode_error_CM_RX_SMP_HOG_WM;
input handcode_error_CM_RX_SMP_PAUSE_WM_t  handcode_error_CM_RX_SMP_PAUSE_WM;
input handcode_error_CM_RX_SMP_PRIVATE_WM_t  handcode_error_CM_RX_SMP_PRIVATE_WM;
input handcode_error_CM_RX_SMP_USAGE_t  handcode_error_CM_RX_SMP_USAGE;
input handcode_error_CM_RX_SMP_USAGE_MAX_t  handcode_error_CM_RX_SMP_USAGE_MAX;
input handcode_error_CM_RX_SMP_USAGE_MAX_CTRL_t  handcode_error_CM_RX_SMP_USAGE_MAX_CTRL;
input handcode_error_CM_SHARED_SMP_PAUSE_CFG_t  handcode_error_CM_SHARED_SMP_PAUSE_CFG;
input handcode_error_CM_SHARED_SMP_PAUSE_WM_t  handcode_error_CM_SHARED_SMP_PAUSE_WM;
input handcode_error_CM_SHARED_SMP_USAGE_t  handcode_error_CM_SHARED_SMP_USAGE;
input handcode_error_CM_SHARED_WM_t  handcode_error_CM_SHARED_WM;
input handcode_error_CM_SMP_USAGE_t  handcode_error_CM_SMP_USAGE;
input handcode_error_CM_SOFTDROP_WM_t  handcode_error_CM_SOFTDROP_WM;
input handcode_error_CM_TX_EWMA_t  handcode_error_CM_TX_EWMA;
input handcode_error_CM_TX_TC_HOG_WM_t  handcode_error_CM_TX_TC_HOG_WM;
input handcode_error_CM_TX_TC_PRIVATE_WM_t  handcode_error_CM_TX_TC_PRIVATE_WM;
input handcode_error_CM_TX_TC_USAGE_t  handcode_error_CM_TX_TC_USAGE;


    // Register Outputs
output CM_GLOBAL_CFG_t  CM_GLOBAL_CFG;
output CM_GLOBAL_USAGE_t  CM_GLOBAL_USAGE;
output CM_GLOBAL_USAGE_MAX_t  CM_GLOBAL_USAGE_MAX;
output CM_GLOBAL_WM_t  CM_GLOBAL_WM;
output CM_SWEEPER_TC_TO_SMP_t  CM_SWEEPER_TC_TO_SMP;


    // Register signals for HandCoded registers
output CM_AQM_DCTCP_CFG_t  handcode_reg_wdata_CM_AQM_DCTCP_CFG;
output CM_AQM_EWMA_CFG_t  handcode_reg_wdata_CM_AQM_EWMA_CFG;
output CM_FORCE_PAUSE_CFG_t  handcode_reg_wdata_CM_FORCE_PAUSE_CFG;
output CM_MCAST_EPOCH_USAGE_t  handcode_reg_wdata_CM_MCAST_EPOCH_USAGE;
output CM_PAUSE_GEN_STATE_t  handcode_reg_wdata_CM_PAUSE_GEN_STATE;
output CM_PAUSE_PHYS_PORT_CFG_t  handcode_reg_wdata_CM_PAUSE_PHYS_PORT_CFG;
output CM_RX_SMP_HOG_WM_t  handcode_reg_wdata_CM_RX_SMP_HOG_WM;
output CM_RX_SMP_PAUSE_WM_t  handcode_reg_wdata_CM_RX_SMP_PAUSE_WM;
output CM_RX_SMP_PRIVATE_WM_t  handcode_reg_wdata_CM_RX_SMP_PRIVATE_WM;
output CM_RX_SMP_USAGE_t  handcode_reg_wdata_CM_RX_SMP_USAGE;
output CM_RX_SMP_USAGE_MAX_t  handcode_reg_wdata_CM_RX_SMP_USAGE_MAX;
output CM_RX_SMP_USAGE_MAX_CTRL_t  handcode_reg_wdata_CM_RX_SMP_USAGE_MAX_CTRL;
output CM_SHARED_SMP_PAUSE_CFG_t  handcode_reg_wdata_CM_SHARED_SMP_PAUSE_CFG;
output CM_SHARED_SMP_PAUSE_WM_t  handcode_reg_wdata_CM_SHARED_SMP_PAUSE_WM;
output CM_SHARED_SMP_USAGE_t  handcode_reg_wdata_CM_SHARED_SMP_USAGE;
output CM_SHARED_WM_t  handcode_reg_wdata_CM_SHARED_WM;
output CM_SMP_USAGE_t  handcode_reg_wdata_CM_SMP_USAGE;
output CM_SOFTDROP_WM_t  handcode_reg_wdata_CM_SOFTDROP_WM;
output CM_TX_EWMA_t  handcode_reg_wdata_CM_TX_EWMA;
output CM_TX_TC_HOG_WM_t  handcode_reg_wdata_CM_TX_TC_HOG_WM;
output CM_TX_TC_PRIVATE_WM_t  handcode_reg_wdata_CM_TX_TC_PRIVATE_WM;
output CM_TX_TC_USAGE_t  handcode_reg_wdata_CM_TX_TC_USAGE;

output we_CM_AQM_DCTCP_CFG_t  we_CM_AQM_DCTCP_CFG;
output we_CM_AQM_EWMA_CFG_t  we_CM_AQM_EWMA_CFG;
output we_CM_FORCE_PAUSE_CFG_t  we_CM_FORCE_PAUSE_CFG;
output we_CM_MCAST_EPOCH_USAGE_t  we_CM_MCAST_EPOCH_USAGE;
output we_CM_PAUSE_GEN_STATE_t  we_CM_PAUSE_GEN_STATE;
output we_CM_PAUSE_PHYS_PORT_CFG_t  we_CM_PAUSE_PHYS_PORT_CFG;
output we_CM_RX_SMP_HOG_WM_t  we_CM_RX_SMP_HOG_WM;
output we_CM_RX_SMP_PAUSE_WM_t  we_CM_RX_SMP_PAUSE_WM;
output we_CM_RX_SMP_PRIVATE_WM_t  we_CM_RX_SMP_PRIVATE_WM;
output we_CM_RX_SMP_USAGE_t  we_CM_RX_SMP_USAGE;
output we_CM_RX_SMP_USAGE_MAX_t  we_CM_RX_SMP_USAGE_MAX;
output we_CM_RX_SMP_USAGE_MAX_CTRL_t  we_CM_RX_SMP_USAGE_MAX_CTRL;
output we_CM_SHARED_SMP_PAUSE_CFG_t  we_CM_SHARED_SMP_PAUSE_CFG;
output we_CM_SHARED_SMP_PAUSE_WM_t  we_CM_SHARED_SMP_PAUSE_WM;
output we_CM_SHARED_SMP_USAGE_t  we_CM_SHARED_SMP_USAGE;
output we_CM_SHARED_WM_t  we_CM_SHARED_WM;
output we_CM_SMP_USAGE_t  we_CM_SMP_USAGE;
output we_CM_SOFTDROP_WM_t  we_CM_SOFTDROP_WM;
output we_CM_TX_EWMA_t  we_CM_TX_EWMA;
output we_CM_TX_TC_HOG_WM_t  we_CM_TX_TC_HOG_WM;
output we_CM_TX_TC_PRIVATE_WM_t  we_CM_TX_TC_PRIVATE_WM;
output we_CM_TX_TC_USAGE_t  we_CM_TX_TC_USAGE;

output re_CM_AQM_DCTCP_CFG_t  re_CM_AQM_DCTCP_CFG;
output re_CM_AQM_EWMA_CFG_t  re_CM_AQM_EWMA_CFG;
output re_CM_FORCE_PAUSE_CFG_t  re_CM_FORCE_PAUSE_CFG;
output re_CM_MCAST_EPOCH_USAGE_t  re_CM_MCAST_EPOCH_USAGE;
output re_CM_PAUSE_GEN_STATE_t  re_CM_PAUSE_GEN_STATE;
output re_CM_PAUSE_PHYS_PORT_CFG_t  re_CM_PAUSE_PHYS_PORT_CFG;
output re_CM_RX_SMP_HOG_WM_t  re_CM_RX_SMP_HOG_WM;
output re_CM_RX_SMP_PAUSE_WM_t  re_CM_RX_SMP_PAUSE_WM;
output re_CM_RX_SMP_PRIVATE_WM_t  re_CM_RX_SMP_PRIVATE_WM;
output re_CM_RX_SMP_USAGE_t  re_CM_RX_SMP_USAGE;
output re_CM_RX_SMP_USAGE_MAX_t  re_CM_RX_SMP_USAGE_MAX;
output re_CM_RX_SMP_USAGE_MAX_CTRL_t  re_CM_RX_SMP_USAGE_MAX_CTRL;
output re_CM_SHARED_SMP_PAUSE_CFG_t  re_CM_SHARED_SMP_PAUSE_CFG;
output re_CM_SHARED_SMP_PAUSE_WM_t  re_CM_SHARED_SMP_PAUSE_WM;
output re_CM_SHARED_SMP_USAGE_t  re_CM_SHARED_SMP_USAGE;
output re_CM_SHARED_WM_t  re_CM_SHARED_WM;
output re_CM_SMP_USAGE_t  re_CM_SMP_USAGE;
output re_CM_SOFTDROP_WM_t  re_CM_SOFTDROP_WM;
output re_CM_TX_EWMA_t  re_CM_TX_EWMA;
output re_CM_TX_TC_HOG_WM_t  re_CM_TX_TC_HOG_WM;
output re_CM_TX_TC_PRIVATE_WM_t  re_CM_TX_TC_PRIVATE_WM;
output re_CM_TX_TC_USAGE_t  re_CM_TX_TC_USAGE;




    // Config Access
input mby_ppe_cm_usage_map_cr_req_t  req;
output mby_ppe_cm_usage_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_cm_usage_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_CM_USAGE_MAP_MEM;
assign case_req_addr_MBY_PPE_CM_USAGE_MAP_MEM = req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_cm_usage;
always_comb begin : sb_fid_cond_cm_usage_BLOCK
    unique casez (req_fid) 
		CM_USAGE_SB_FID: sb_fid_cond_cm_usage = 1;
		default: sb_fid_cond_cm_usage = 0;
    endcase 
end


logic sb_bar_cond_cm_usage;
always_comb begin : sb_bar_cond_cm_usage_BLOCK
    unique casez (req_bar) 
		CM_USAGE_SB_BAR: sb_bar_cond_cm_usage = 1;
		default: sb_bar_cond_cm_usage = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// CM_TX_TC_PRIVATE_WM using HANDCODED_REG template.
logic addr_decode_CM_TX_TC_PRIVATE_WM;
logic write_req_CM_TX_TC_PRIVATE_WM;
logic read_req_CM_TX_TC_PRIVATE_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h0??,1'b?}: 
         addr_decode_CM_TX_TC_PRIVATE_WM = req.valid;
      default: 
         addr_decode_CM_TX_TC_PRIVATE_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_TX_TC_PRIVATE_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_TX_TC_PRIVATE_WM ;
always_comb read_req_CM_TX_TC_PRIVATE_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_TX_TC_PRIVATE_WM ;

always_comb we_CM_TX_TC_PRIVATE_WM = {8{write_req_CM_TX_TC_PRIVATE_WM}} & be;
always_comb re_CM_TX_TC_PRIVATE_WM = {8{read_req_CM_TX_TC_PRIVATE_WM}} & be;
always_comb handcode_reg_wdata_CM_TX_TC_PRIVATE_WM = write_data;


// ----------------------------------------------------------------------
// CM_TX_TC_HOG_WM using HANDCODED_REG template.
logic addr_decode_CM_TX_TC_HOG_WM;
logic write_req_CM_TX_TC_HOG_WM;
logic read_req_CM_TX_TC_HOG_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h1??,1'b?}: 
         addr_decode_CM_TX_TC_HOG_WM = req.valid;
      default: 
         addr_decode_CM_TX_TC_HOG_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_TX_TC_HOG_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_TX_TC_HOG_WM ;
always_comb read_req_CM_TX_TC_HOG_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_TX_TC_HOG_WM ;

always_comb we_CM_TX_TC_HOG_WM = {8{write_req_CM_TX_TC_HOG_WM}} & be;
always_comb re_CM_TX_TC_HOG_WM = {8{read_req_CM_TX_TC_HOG_WM}} & be;
always_comb handcode_reg_wdata_CM_TX_TC_HOG_WM = write_data;


// ----------------------------------------------------------------------
// CM_RX_SMP_PRIVATE_WM using HANDCODED_REG template.
logic addr_decode_CM_RX_SMP_PRIVATE_WM;
logic write_req_CM_RX_SMP_PRIVATE_WM;
logic read_req_CM_RX_SMP_PRIVATE_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h2,4'b000?,4'h?,1'b?}: 
         addr_decode_CM_RX_SMP_PRIVATE_WM = req.valid;
      default: 
         addr_decode_CM_RX_SMP_PRIVATE_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_RX_SMP_PRIVATE_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_RX_SMP_PRIVATE_WM ;
always_comb read_req_CM_RX_SMP_PRIVATE_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_RX_SMP_PRIVATE_WM ;

always_comb we_CM_RX_SMP_PRIVATE_WM = {8{write_req_CM_RX_SMP_PRIVATE_WM}} & be;
always_comb re_CM_RX_SMP_PRIVATE_WM = {8{read_req_CM_RX_SMP_PRIVATE_WM}} & be;
always_comb handcode_reg_wdata_CM_RX_SMP_PRIVATE_WM = write_data;


// ----------------------------------------------------------------------
// CM_RX_SMP_HOG_WM using HANDCODED_REG template.
logic addr_decode_CM_RX_SMP_HOG_WM;
logic write_req_CM_RX_SMP_HOG_WM;
logic read_req_CM_RX_SMP_HOG_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h2,4'b001?,4'h?,1'b?}: 
         addr_decode_CM_RX_SMP_HOG_WM = req.valid;
      default: 
         addr_decode_CM_RX_SMP_HOG_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_RX_SMP_HOG_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_RX_SMP_HOG_WM ;
always_comb read_req_CM_RX_SMP_HOG_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_RX_SMP_HOG_WM ;

always_comb we_CM_RX_SMP_HOG_WM = {8{write_req_CM_RX_SMP_HOG_WM}} & be;
always_comb re_CM_RX_SMP_HOG_WM = {8{read_req_CM_RX_SMP_HOG_WM}} & be;
always_comb handcode_reg_wdata_CM_RX_SMP_HOG_WM = write_data;


// ----------------------------------------------------------------------
// CM_RX_SMP_PAUSE_WM using HANDCODED_REG template.
logic addr_decode_CM_RX_SMP_PAUSE_WM;
logic write_req_CM_RX_SMP_PAUSE_WM;
logic read_req_CM_RX_SMP_PAUSE_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h2,4'b010?,4'h?,1'b?}: 
         addr_decode_CM_RX_SMP_PAUSE_WM = req.valid;
      default: 
         addr_decode_CM_RX_SMP_PAUSE_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_RX_SMP_PAUSE_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_RX_SMP_PAUSE_WM ;
always_comb read_req_CM_RX_SMP_PAUSE_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_RX_SMP_PAUSE_WM ;

always_comb we_CM_RX_SMP_PAUSE_WM = {8{write_req_CM_RX_SMP_PAUSE_WM}} & be;
always_comb re_CM_RX_SMP_PAUSE_WM = {8{read_req_CM_RX_SMP_PAUSE_WM}} & be;
always_comb handcode_reg_wdata_CM_RX_SMP_PAUSE_WM = write_data;


// ----------------------------------------------------------------------
// CM_SHARED_WM using HANDCODED_REG template.
logic addr_decode_CM_SHARED_WM;
logic write_req_CM_SHARED_WM;
logic read_req_CM_SHARED_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h26,4'b00??,1'b?}: 
         addr_decode_CM_SHARED_WM = req.valid;
      default: 
         addr_decode_CM_SHARED_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_SHARED_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_SHARED_WM ;
always_comb read_req_CM_SHARED_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_SHARED_WM ;

always_comb we_CM_SHARED_WM = {8{write_req_CM_SHARED_WM}} & be;
always_comb re_CM_SHARED_WM = {8{read_req_CM_SHARED_WM}} & be;
always_comb handcode_reg_wdata_CM_SHARED_WM = write_data;


// ----------------------------------------------------------------------
// CM_SOFTDROP_WM using HANDCODED_REG template.
logic addr_decode_CM_SOFTDROP_WM;
logic write_req_CM_SOFTDROP_WM;
logic read_req_CM_SOFTDROP_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h26,4'b01??,1'b?}: 
         addr_decode_CM_SOFTDROP_WM = req.valid;
      default: 
         addr_decode_CM_SOFTDROP_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_SOFTDROP_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_SOFTDROP_WM ;
always_comb read_req_CM_SOFTDROP_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_SOFTDROP_WM ;

always_comb we_CM_SOFTDROP_WM = {8{write_req_CM_SOFTDROP_WM}} & be;
always_comb re_CM_SOFTDROP_WM = {8{read_req_CM_SOFTDROP_WM}} & be;
always_comb handcode_reg_wdata_CM_SOFTDROP_WM = write_data;


// ----------------------------------------------------------------------
// CM_SHARED_SMP_PAUSE_WM using HANDCODED_REG template.
logic addr_decode_CM_SHARED_SMP_PAUSE_WM;
logic write_req_CM_SHARED_SMP_PAUSE_WM;
logic read_req_CM_SHARED_SMP_PAUSE_WM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h268,1'b?}: 
         addr_decode_CM_SHARED_SMP_PAUSE_WM = req.valid;
      default: 
         addr_decode_CM_SHARED_SMP_PAUSE_WM = 1'b0; 
   endcase
end

always_comb write_req_CM_SHARED_SMP_PAUSE_WM = f_IsMEMWr(req_opcode) && addr_decode_CM_SHARED_SMP_PAUSE_WM ;
always_comb read_req_CM_SHARED_SMP_PAUSE_WM  = f_IsMEMRd(req_opcode) && addr_decode_CM_SHARED_SMP_PAUSE_WM ;

always_comb we_CM_SHARED_SMP_PAUSE_WM = {8{write_req_CM_SHARED_SMP_PAUSE_WM}} & be;
always_comb re_CM_SHARED_SMP_PAUSE_WM = {8{read_req_CM_SHARED_SMP_PAUSE_WM}} & be;
always_comb handcode_reg_wdata_CM_SHARED_SMP_PAUSE_WM = write_data;


//---------------------------------------------------------------------
// CM_GLOBAL_WM Address Decode
logic  addr_decode_CM_GLOBAL_WM;
logic  write_req_CM_GLOBAL_WM;
always_comb begin
   addr_decode_CM_GLOBAL_WM = (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_GLOBAL_WM_DECODE_ADDR) && req.valid ;
   write_req_CM_GLOBAL_WM = IsMEMWr && addr_decode_CM_GLOBAL_WM && sb_fid_cond_cm_usage && sb_bar_cond_cm_usage;
end

// ----------------------------------------------------------------------
// CM_GLOBAL_WM.WATERMARK x7 RW, using RW template.
logic [1:0] up_CM_GLOBAL_WM_WATERMARK;
always_comb begin
 up_CM_GLOBAL_WM_WATERMARK =
    ({2{write_req_CM_GLOBAL_WM }} &
    be[1:0]);
end

logic [14:0] nxt_CM_GLOBAL_WM_WATERMARK;
always_comb begin
 nxt_CM_GLOBAL_WM_WATERMARK = write_data[14:0];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 8'h20, up_CM_GLOBAL_WM_WATERMARK[0], nxt_CM_GLOBAL_WM_WATERMARK[7:0], CM_GLOBAL_WM.WATERMARK[7:0])
`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 7'h5E, up_CM_GLOBAL_WM_WATERMARK[1], nxt_CM_GLOBAL_WM_WATERMARK[14:8], CM_GLOBAL_WM.WATERMARK[14:8])

// ----------------------------------------------------------------------
// CM_PAUSE_PHYS_PORT_CFG using HANDCODED_REG template.
logic addr_decode_CM_PAUSE_PHYS_PORT_CFG;
logic write_req_CM_PAUSE_PHYS_PORT_CFG;
logic read_req_CM_PAUSE_PHYS_PORT_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h27?,1'b?}: 
         addr_decode_CM_PAUSE_PHYS_PORT_CFG = req.valid;
      default: 
         addr_decode_CM_PAUSE_PHYS_PORT_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_PAUSE_PHYS_PORT_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_PAUSE_PHYS_PORT_CFG ;
always_comb read_req_CM_PAUSE_PHYS_PORT_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_PAUSE_PHYS_PORT_CFG ;

always_comb we_CM_PAUSE_PHYS_PORT_CFG = {8{write_req_CM_PAUSE_PHYS_PORT_CFG}} & be;
always_comb re_CM_PAUSE_PHYS_PORT_CFG = {8{read_req_CM_PAUSE_PHYS_PORT_CFG}} & be;
always_comb handcode_reg_wdata_CM_PAUSE_PHYS_PORT_CFG = write_data;


// ----------------------------------------------------------------------
// CM_FORCE_PAUSE_CFG using HANDCODED_REG template.
logic addr_decode_CM_FORCE_PAUSE_CFG;
logic write_req_CM_FORCE_PAUSE_CFG;
logic read_req_CM_FORCE_PAUSE_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h280,1'b0}: 
         addr_decode_CM_FORCE_PAUSE_CFG = req.valid;
      default: 
         addr_decode_CM_FORCE_PAUSE_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_FORCE_PAUSE_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_FORCE_PAUSE_CFG ;
always_comb read_req_CM_FORCE_PAUSE_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_FORCE_PAUSE_CFG ;

always_comb we_CM_FORCE_PAUSE_CFG = {8{write_req_CM_FORCE_PAUSE_CFG}} & be;
always_comb re_CM_FORCE_PAUSE_CFG = {8{read_req_CM_FORCE_PAUSE_CFG}} & be;
always_comb handcode_reg_wdata_CM_FORCE_PAUSE_CFG = write_data;


// ----------------------------------------------------------------------
// CM_AQM_EWMA_CFG using HANDCODED_REG template.
logic addr_decode_CM_AQM_EWMA_CFG;
logic write_req_CM_AQM_EWMA_CFG;
logic read_req_CM_AQM_EWMA_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h2,4'b11??,4'h?,1'b?}: 
         addr_decode_CM_AQM_EWMA_CFG = req.valid;
      default: 
         addr_decode_CM_AQM_EWMA_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_AQM_EWMA_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_AQM_EWMA_CFG ;
always_comb read_req_CM_AQM_EWMA_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_AQM_EWMA_CFG ;

always_comb we_CM_AQM_EWMA_CFG = {8{write_req_CM_AQM_EWMA_CFG}} & be;
always_comb re_CM_AQM_EWMA_CFG = {8{read_req_CM_AQM_EWMA_CFG}} & be;
always_comb handcode_reg_wdata_CM_AQM_EWMA_CFG = write_data;


// ----------------------------------------------------------------------
// CM_AQM_DCTCP_CFG using HANDCODED_REG template.
logic addr_decode_CM_AQM_DCTCP_CFG;
logic write_req_CM_AQM_DCTCP_CFG;
logic read_req_CM_AQM_DCTCP_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h3,4'b00??,4'h?,1'b?}: 
         addr_decode_CM_AQM_DCTCP_CFG = req.valid;
      default: 
         addr_decode_CM_AQM_DCTCP_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_AQM_DCTCP_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_AQM_DCTCP_CFG ;
always_comb read_req_CM_AQM_DCTCP_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_AQM_DCTCP_CFG ;

always_comb we_CM_AQM_DCTCP_CFG = {8{write_req_CM_AQM_DCTCP_CFG}} & be;
always_comb re_CM_AQM_DCTCP_CFG = {8{read_req_CM_AQM_DCTCP_CFG}} & be;
always_comb handcode_reg_wdata_CM_AQM_DCTCP_CFG = write_data;


//---------------------------------------------------------------------
// CM_GLOBAL_CFG Address Decode
logic  addr_decode_CM_GLOBAL_CFG;
logic  write_req_CM_GLOBAL_CFG;
always_comb begin
   addr_decode_CM_GLOBAL_CFG = (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_GLOBAL_CFG_DECODE_ADDR) && req.valid ;
   write_req_CM_GLOBAL_CFG = IsMEMWr && addr_decode_CM_GLOBAL_CFG && sb_fid_cond_cm_usage && sb_bar_cond_cm_usage;
end

// ----------------------------------------------------------------------
// CM_GLOBAL_CFG.NUM_SWEEPER_PORTS x5 RW, using RW template.
logic [0:0] up_CM_GLOBAL_CFG_NUM_SWEEPER_PORTS;
always_comb begin
 up_CM_GLOBAL_CFG_NUM_SWEEPER_PORTS =
    ({1{write_req_CM_GLOBAL_CFG }} &
    be[0:0]);
end

logic [4:0] nxt_CM_GLOBAL_CFG_NUM_SWEEPER_PORTS;
always_comb begin
 nxt_CM_GLOBAL_CFG_NUM_SWEEPER_PORTS = write_data[4:0];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 5'h0, up_CM_GLOBAL_CFG_NUM_SWEEPER_PORTS[0], nxt_CM_GLOBAL_CFG_NUM_SWEEPER_PORTS[4:0], CM_GLOBAL_CFG.NUM_SWEEPER_PORTS[4:0])

// ----------------------------------------------------------------------
// CM_GLOBAL_CFG.SWEEPER_EN x1 RW, using RW template.
logic [0:0] up_CM_GLOBAL_CFG_SWEEPER_EN;
always_comb begin
 up_CM_GLOBAL_CFG_SWEEPER_EN =
    ({1{write_req_CM_GLOBAL_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_CM_GLOBAL_CFG_SWEEPER_EN;
always_comb begin
 nxt_CM_GLOBAL_CFG_SWEEPER_EN = write_data[5:5];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_GLOBAL_CFG_SWEEPER_EN[0], nxt_CM_GLOBAL_CFG_SWEEPER_EN[0:0], CM_GLOBAL_CFG.SWEEPER_EN[0:0])

// ----------------------------------------------------------------------
// CM_SHARED_SMP_PAUSE_CFG using HANDCODED_REG template.
logic addr_decode_CM_SHARED_SMP_PAUSE_CFG;
logic write_req_CM_SHARED_SMP_PAUSE_CFG;
logic read_req_CM_SHARED_SMP_PAUSE_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h341,1'b?}: 
         addr_decode_CM_SHARED_SMP_PAUSE_CFG = req.valid;
      default: 
         addr_decode_CM_SHARED_SMP_PAUSE_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_SHARED_SMP_PAUSE_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_SHARED_SMP_PAUSE_CFG ;
always_comb read_req_CM_SHARED_SMP_PAUSE_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_SHARED_SMP_PAUSE_CFG ;

always_comb we_CM_SHARED_SMP_PAUSE_CFG = {8{write_req_CM_SHARED_SMP_PAUSE_CFG}} & be;
always_comb re_CM_SHARED_SMP_PAUSE_CFG = {8{read_req_CM_SHARED_SMP_PAUSE_CFG}} & be;
always_comb handcode_reg_wdata_CM_SHARED_SMP_PAUSE_CFG = write_data;


//---------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP Address Decode
logic  addr_decode_CM_SWEEPER_TC_TO_SMP;
logic  write_req_CM_SWEEPER_TC_TO_SMP;
always_comb begin
   addr_decode_CM_SWEEPER_TC_TO_SMP = (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_SWEEPER_TC_TO_SMP_DECODE_ADDR) && req.valid ;
   write_req_CM_SWEEPER_TC_TO_SMP = IsMEMWr && addr_decode_CM_SWEEPER_TC_TO_SMP && sb_fid_cond_cm_usage && sb_bar_cond_cm_usage;
end

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_0 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_0;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_0 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_0;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_0 = write_data[0:0];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_0[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_0[0:0], CM_SWEEPER_TC_TO_SMP.SMP_0[0:0])

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_1 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_1;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_1 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_1;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_1 = write_data[1:1];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_1[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_1[0:0], CM_SWEEPER_TC_TO_SMP.SMP_1[0:0])

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_2 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_2;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_2 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_2;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_2 = write_data[2:2];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_2[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_2[0:0], CM_SWEEPER_TC_TO_SMP.SMP_2[0:0])

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_3 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_3;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_3 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_3;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_3 = write_data[3:3];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_3[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_3[0:0], CM_SWEEPER_TC_TO_SMP.SMP_3[0:0])

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_4 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_4;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_4 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_4;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_4 = write_data[4:4];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_4[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_4[0:0], CM_SWEEPER_TC_TO_SMP.SMP_4[0:0])

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_5 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_5;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_5 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_5;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_5 = write_data[5:5];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_5[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_5[0:0], CM_SWEEPER_TC_TO_SMP.SMP_5[0:0])

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_6 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_6;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_6 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_6;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_6 = write_data[6:6];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_6[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_6[0:0], CM_SWEEPER_TC_TO_SMP.SMP_6[0:0])

// ----------------------------------------------------------------------
// CM_SWEEPER_TC_TO_SMP.SMP_7 x1 RW, using RW template.
logic [0:0] up_CM_SWEEPER_TC_TO_SMP_SMP_7;
always_comb begin
 up_CM_SWEEPER_TC_TO_SMP_SMP_7 =
    ({1{write_req_CM_SWEEPER_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_SWEEPER_TC_TO_SMP_SMP_7;
always_comb begin
 nxt_CM_SWEEPER_TC_TO_SMP_SMP_7 = write_data[7:7];

end


`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_SWEEPER_TC_TO_SMP_SMP_7[0], nxt_CM_SWEEPER_TC_TO_SMP_SMP_7[0:0], CM_SWEEPER_TC_TO_SMP.SMP_7[0:0])

//---------------------------------------------------------------------
// CM_GLOBAL_USAGE Address Decode
// ----------------------------------------------------------------------
// CM_GLOBAL_USAGE.COUNT x8 RO/V, using RO/V template.
assign CM_GLOBAL_USAGE.COUNT = new_CM_GLOBAL_USAGE.COUNT;




//---------------------------------------------------------------------
// CM_GLOBAL_USAGE_MAX Address Decode
logic  addr_decode_CM_GLOBAL_USAGE_MAX;
logic  write_req_CM_GLOBAL_USAGE_MAX;
always_comb begin
   addr_decode_CM_GLOBAL_USAGE_MAX = (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_GLOBAL_USAGE_MAX_DECODE_ADDR) && req.valid ;
   write_req_CM_GLOBAL_USAGE_MAX = IsMEMWr && addr_decode_CM_GLOBAL_USAGE_MAX && sb_fid_cond_cm_usage && sb_bar_cond_cm_usage;
end

// ----------------------------------------------------------------------
// CM_GLOBAL_USAGE_MAX.COUNT x8 RW/V, using RW/V template.
logic [1:0] req_up_CM_GLOBAL_USAGE_MAX_COUNT;
always_comb begin
 req_up_CM_GLOBAL_USAGE_MAX_COUNT[0] = 
   {write_req_CM_GLOBAL_USAGE_MAX & be[0]}
;
 req_up_CM_GLOBAL_USAGE_MAX_COUNT[1] = 
   {write_req_CM_GLOBAL_USAGE_MAX & be[1]}
;
end

logic [1:0] swwr_CM_GLOBAL_USAGE_MAX_COUNT;
always_comb begin
 swwr_CM_GLOBAL_USAGE_MAX_COUNT = req_up_CM_GLOBAL_USAGE_MAX_COUNT;

end


logic [1:0] up_CM_GLOBAL_USAGE_MAX_COUNT;
logic [15:0] nxt_CM_GLOBAL_USAGE_MAX_COUNT;
always_comb begin
 up_CM_GLOBAL_USAGE_MAX_COUNT =
    swwr_CM_GLOBAL_USAGE_MAX_COUNT |
    {2{load_CM_GLOBAL_USAGE_MAX.COUNT}};
end
always_comb begin
 nxt_CM_GLOBAL_USAGE_MAX_COUNT[7:0] = 
    swwr_CM_GLOBAL_USAGE_MAX_COUNT[0] ?
    write_data[7:0] :
    new_CM_GLOBAL_USAGE_MAX.COUNT[7:0];
 nxt_CM_GLOBAL_USAGE_MAX_COUNT[15:8] = 
    swwr_CM_GLOBAL_USAGE_MAX_COUNT[1] ?
    write_data[15:8] :
    new_CM_GLOBAL_USAGE_MAX.COUNT[15:8];
end

`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(rtl_clk, rst_n, 8'h0, up_CM_GLOBAL_USAGE_MAX_COUNT[0], nxt_CM_GLOBAL_USAGE_MAX_COUNT[7:0], CM_GLOBAL_USAGE_MAX.COUNT[7:0])
`RTLGEN_MBY_PPE_CM_USAGE_MAP_EN_FF(rtl_clk, rst_n, 8'h0, up_CM_GLOBAL_USAGE_MAX_COUNT[1], nxt_CM_GLOBAL_USAGE_MAX_COUNT[15:8], CM_GLOBAL_USAGE_MAX.COUNT[15:8])

// ----------------------------------------------------------------------
// CM_MCAST_EPOCH_USAGE using HANDCODED_REG template.
logic addr_decode_CM_MCAST_EPOCH_USAGE;
logic write_req_CM_MCAST_EPOCH_USAGE;
logic read_req_CM_MCAST_EPOCH_USAGE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h344,1'b?}: 
         addr_decode_CM_MCAST_EPOCH_USAGE = req.valid;
      default: 
         addr_decode_CM_MCAST_EPOCH_USAGE = 1'b0; 
   endcase
end

always_comb write_req_CM_MCAST_EPOCH_USAGE = f_IsMEMWr(req_opcode) && addr_decode_CM_MCAST_EPOCH_USAGE ;
always_comb read_req_CM_MCAST_EPOCH_USAGE  = f_IsMEMRd(req_opcode) && addr_decode_CM_MCAST_EPOCH_USAGE ;

always_comb we_CM_MCAST_EPOCH_USAGE = {8{write_req_CM_MCAST_EPOCH_USAGE}} & be;
always_comb re_CM_MCAST_EPOCH_USAGE = {8{read_req_CM_MCAST_EPOCH_USAGE}} & be;
always_comb handcode_reg_wdata_CM_MCAST_EPOCH_USAGE = write_data;


// ----------------------------------------------------------------------
// CM_SHARED_SMP_USAGE using HANDCODED_REG template.
logic addr_decode_CM_SHARED_SMP_USAGE;
logic write_req_CM_SHARED_SMP_USAGE;
logic read_req_CM_SHARED_SMP_USAGE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h345,1'b?}: 
         addr_decode_CM_SHARED_SMP_USAGE = req.valid;
      default: 
         addr_decode_CM_SHARED_SMP_USAGE = 1'b0; 
   endcase
end

always_comb write_req_CM_SHARED_SMP_USAGE = f_IsMEMWr(req_opcode) && addr_decode_CM_SHARED_SMP_USAGE ;
always_comb read_req_CM_SHARED_SMP_USAGE  = f_IsMEMRd(req_opcode) && addr_decode_CM_SHARED_SMP_USAGE ;

always_comb we_CM_SHARED_SMP_USAGE = {8{write_req_CM_SHARED_SMP_USAGE}} & be;
always_comb re_CM_SHARED_SMP_USAGE = {8{read_req_CM_SHARED_SMP_USAGE}} & be;
always_comb handcode_reg_wdata_CM_SHARED_SMP_USAGE = write_data;


// ----------------------------------------------------------------------
// CM_SMP_USAGE using HANDCODED_REG template.
logic addr_decode_CM_SMP_USAGE;
logic write_req_CM_SMP_USAGE;
logic read_req_CM_SMP_USAGE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h346,1'b?}: 
         addr_decode_CM_SMP_USAGE = req.valid;
      default: 
         addr_decode_CM_SMP_USAGE = 1'b0; 
   endcase
end

always_comb write_req_CM_SMP_USAGE = f_IsMEMWr(req_opcode) && addr_decode_CM_SMP_USAGE ;
always_comb read_req_CM_SMP_USAGE  = f_IsMEMRd(req_opcode) && addr_decode_CM_SMP_USAGE ;

always_comb we_CM_SMP_USAGE = {8{write_req_CM_SMP_USAGE}} & be;
always_comb re_CM_SMP_USAGE = {8{read_req_CM_SMP_USAGE}} & be;
always_comb handcode_reg_wdata_CM_SMP_USAGE = write_data;


// ----------------------------------------------------------------------
// CM_RX_SMP_USAGE using HANDCODED_REG template.
logic addr_decode_CM_RX_SMP_USAGE;
logic write_req_CM_RX_SMP_USAGE;
logic read_req_CM_RX_SMP_USAGE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h3,4'b011?,4'h?,1'b?}: 
         addr_decode_CM_RX_SMP_USAGE = req.valid;
      default: 
         addr_decode_CM_RX_SMP_USAGE = 1'b0; 
   endcase
end

always_comb write_req_CM_RX_SMP_USAGE = f_IsMEMWr(req_opcode) && addr_decode_CM_RX_SMP_USAGE ;
always_comb read_req_CM_RX_SMP_USAGE  = f_IsMEMRd(req_opcode) && addr_decode_CM_RX_SMP_USAGE ;

always_comb we_CM_RX_SMP_USAGE = {8{write_req_CM_RX_SMP_USAGE}} & be;
always_comb re_CM_RX_SMP_USAGE = {8{read_req_CM_RX_SMP_USAGE}} & be;
always_comb handcode_reg_wdata_CM_RX_SMP_USAGE = write_data;


// ----------------------------------------------------------------------
// CM_RX_SMP_USAGE_MAX using HANDCODED_REG template.
logic addr_decode_CM_RX_SMP_USAGE_MAX;
logic write_req_CM_RX_SMP_USAGE_MAX;
logic read_req_CM_RX_SMP_USAGE_MAX;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h38,4'b00??,1'b?}: 
         addr_decode_CM_RX_SMP_USAGE_MAX = req.valid;
      default: 
         addr_decode_CM_RX_SMP_USAGE_MAX = 1'b0; 
   endcase
end

always_comb write_req_CM_RX_SMP_USAGE_MAX = f_IsMEMWr(req_opcode) && addr_decode_CM_RX_SMP_USAGE_MAX ;
always_comb read_req_CM_RX_SMP_USAGE_MAX  = f_IsMEMRd(req_opcode) && addr_decode_CM_RX_SMP_USAGE_MAX ;

always_comb we_CM_RX_SMP_USAGE_MAX = {8{write_req_CM_RX_SMP_USAGE_MAX}} & be;
always_comb re_CM_RX_SMP_USAGE_MAX = {8{read_req_CM_RX_SMP_USAGE_MAX}} & be;
always_comb handcode_reg_wdata_CM_RX_SMP_USAGE_MAX = write_data;


// ----------------------------------------------------------------------
// CM_RX_SMP_USAGE_MAX_CTRL using HANDCODED_REG template.
logic addr_decode_CM_RX_SMP_USAGE_MAX_CTRL;
logic write_req_CM_RX_SMP_USAGE_MAX_CTRL;
logic read_req_CM_RX_SMP_USAGE_MAX_CTRL;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h384,1'b0}: 
         addr_decode_CM_RX_SMP_USAGE_MAX_CTRL = req.valid;
      default: 
         addr_decode_CM_RX_SMP_USAGE_MAX_CTRL = 1'b0; 
   endcase
end

always_comb write_req_CM_RX_SMP_USAGE_MAX_CTRL = f_IsMEMWr(req_opcode) && addr_decode_CM_RX_SMP_USAGE_MAX_CTRL ;
always_comb read_req_CM_RX_SMP_USAGE_MAX_CTRL  = f_IsMEMRd(req_opcode) && addr_decode_CM_RX_SMP_USAGE_MAX_CTRL ;

always_comb we_CM_RX_SMP_USAGE_MAX_CTRL = {8{write_req_CM_RX_SMP_USAGE_MAX_CTRL}} & be;
always_comb re_CM_RX_SMP_USAGE_MAX_CTRL = {8{read_req_CM_RX_SMP_USAGE_MAX_CTRL}} & be;
always_comb handcode_reg_wdata_CM_RX_SMP_USAGE_MAX_CTRL = write_data;


// ----------------------------------------------------------------------
// CM_PAUSE_GEN_STATE using HANDCODED_REG template.
logic addr_decode_CM_PAUSE_GEN_STATE;
logic write_req_CM_PAUSE_GEN_STATE;
logic read_req_CM_PAUSE_GEN_STATE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h39?,1'b?}: 
         addr_decode_CM_PAUSE_GEN_STATE = req.valid;
      default: 
         addr_decode_CM_PAUSE_GEN_STATE = 1'b0; 
   endcase
end

always_comb write_req_CM_PAUSE_GEN_STATE = f_IsMEMWr(req_opcode) && addr_decode_CM_PAUSE_GEN_STATE ;
always_comb read_req_CM_PAUSE_GEN_STATE  = f_IsMEMRd(req_opcode) && addr_decode_CM_PAUSE_GEN_STATE ;

always_comb we_CM_PAUSE_GEN_STATE = {8{write_req_CM_PAUSE_GEN_STATE}} & be;
always_comb re_CM_PAUSE_GEN_STATE = {8{read_req_CM_PAUSE_GEN_STATE}} & be;
always_comb handcode_reg_wdata_CM_PAUSE_GEN_STATE = write_data;


// ----------------------------------------------------------------------
// CM_TX_TC_USAGE using HANDCODED_REG template.
logic addr_decode_CM_TX_TC_USAGE;
logic write_req_CM_TX_TC_USAGE;
logic read_req_CM_TX_TC_USAGE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h4??,1'b?}: 
         addr_decode_CM_TX_TC_USAGE = req.valid;
      default: 
         addr_decode_CM_TX_TC_USAGE = 1'b0; 
   endcase
end

always_comb write_req_CM_TX_TC_USAGE = f_IsMEMWr(req_opcode) && addr_decode_CM_TX_TC_USAGE ;
always_comb read_req_CM_TX_TC_USAGE  = f_IsMEMRd(req_opcode) && addr_decode_CM_TX_TC_USAGE ;

always_comb we_CM_TX_TC_USAGE = {8{write_req_CM_TX_TC_USAGE}} & be;
always_comb re_CM_TX_TC_USAGE = {8{read_req_CM_TX_TC_USAGE}} & be;
always_comb handcode_reg_wdata_CM_TX_TC_USAGE = write_data;


// ----------------------------------------------------------------------
// CM_TX_EWMA using HANDCODED_REG template.
logic addr_decode_CM_TX_EWMA;
logic write_req_CM_TX_EWMA;
logic read_req_CM_TX_EWMA;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_USAGE_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h5,4'b00??,4'h?,1'b?}: 
         addr_decode_CM_TX_EWMA = req.valid;
      default: 
         addr_decode_CM_TX_EWMA = 1'b0; 
   endcase
end

always_comb write_req_CM_TX_EWMA = f_IsMEMWr(req_opcode) && addr_decode_CM_TX_EWMA ;
always_comb read_req_CM_TX_EWMA  = f_IsMEMRd(req_opcode) && addr_decode_CM_TX_EWMA ;

always_comb we_CM_TX_EWMA = {8{write_req_CM_TX_EWMA}} & be;
always_comb re_CM_TX_EWMA = {8{read_req_CM_TX_EWMA}} & be;
always_comb handcode_reg_wdata_CM_TX_EWMA = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_CM_USAGE_MAP_MEM) 
           {44'h0??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_TX_TC_PRIVATE_WM;
                    ack.read_miss = handcode_error_CM_TX_TC_PRIVATE_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h1??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_TX_TC_HOG_WM;
                    ack.read_miss = handcode_error_CM_TX_TC_HOG_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h2,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_RX_SMP_PRIVATE_WM;
                    ack.read_miss = handcode_error_CM_RX_SMP_PRIVATE_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h2,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_RX_SMP_HOG_WM;
                    ack.read_miss = handcode_error_CM_RX_SMP_HOG_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h2,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_RX_SMP_PAUSE_WM;
                    ack.read_miss = handcode_error_CM_RX_SMP_PAUSE_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h26,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_SHARED_WM;
                    ack.read_miss = handcode_error_CM_SHARED_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h26,4'b01??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_SOFTDROP_WM;
                    ack.read_miss = handcode_error_CM_SOFTDROP_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h268,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_SHARED_SMP_PAUSE_WM;
                    ack.read_miss = handcode_error_CM_SHARED_SMP_PAUSE_WM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_GLOBAL_WM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h27?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_PAUSE_PHYS_PORT_CFG;
                    ack.read_miss = handcode_error_CM_PAUSE_PHYS_PORT_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h280,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_FORCE_PAUSE_CFG;
                    ack.read_miss = handcode_error_CM_FORCE_PAUSE_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h2,4'b11??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_AQM_EWMA_CFG;
                    ack.read_miss = handcode_error_CM_AQM_EWMA_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h3,4'b00??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_AQM_DCTCP_CFG;
                    ack.read_miss = handcode_error_CM_AQM_DCTCP_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_GLOBAL_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h341,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_SHARED_SMP_PAUSE_CFG;
                    ack.read_miss = handcode_error_CM_SHARED_SMP_PAUSE_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_SWEEPER_TC_TO_SMP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_GLOBAL_USAGE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_GLOBAL_USAGE_MAX_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h344,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_MCAST_EPOCH_USAGE;
                    ack.read_miss = handcode_error_CM_MCAST_EPOCH_USAGE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h345,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_SHARED_SMP_USAGE;
                    ack.read_miss = handcode_error_CM_SHARED_SMP_USAGE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h346,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_SMP_USAGE;
                    ack.read_miss = handcode_error_CM_SMP_USAGE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h3,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_RX_SMP_USAGE;
                    ack.read_miss = handcode_error_CM_RX_SMP_USAGE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h38,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_RX_SMP_USAGE_MAX;
                    ack.read_miss = handcode_error_CM_RX_SMP_USAGE_MAX;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h384,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_RX_SMP_USAGE_MAX_CTRL;
                    ack.read_miss = handcode_error_CM_RX_SMP_USAGE_MAX_CTRL;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h39?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_PAUSE_GEN_STATE;
                    ack.read_miss = handcode_error_CM_PAUSE_GEN_STATE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h4??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_TX_TC_USAGE;
                    ack.read_miss = handcode_error_CM_TX_TC_USAGE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h5,4'b00??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_TX_EWMA;
                    ack.read_miss = handcode_error_CM_TX_EWMA;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_CM_USAGE_MAP_MEM) 
           {44'h0??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_TX_TC_PRIVATE_WM;
                    ack.write_miss = handcode_error_CM_TX_TC_PRIVATE_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h1??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_TX_TC_HOG_WM;
                    ack.write_miss = handcode_error_CM_TX_TC_HOG_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h2,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_RX_SMP_PRIVATE_WM;
                    ack.write_miss = handcode_error_CM_RX_SMP_PRIVATE_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h2,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_RX_SMP_HOG_WM;
                    ack.write_miss = handcode_error_CM_RX_SMP_HOG_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h2,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_RX_SMP_PAUSE_WM;
                    ack.write_miss = handcode_error_CM_RX_SMP_PAUSE_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h26,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_SHARED_WM;
                    ack.write_miss = handcode_error_CM_SHARED_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h26,4'b01??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_SOFTDROP_WM;
                    ack.write_miss = handcode_error_CM_SOFTDROP_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h268,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_SHARED_SMP_PAUSE_WM;
                    ack.write_miss = handcode_error_CM_SHARED_SMP_PAUSE_WM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_GLOBAL_WM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h27?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_PAUSE_PHYS_PORT_CFG;
                    ack.write_miss = handcode_error_CM_PAUSE_PHYS_PORT_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h280,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_FORCE_PAUSE_CFG;
                    ack.write_miss = handcode_error_CM_FORCE_PAUSE_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h2,4'b11??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_AQM_EWMA_CFG;
                    ack.write_miss = handcode_error_CM_AQM_EWMA_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h3,4'b00??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_AQM_DCTCP_CFG;
                    ack.write_miss = handcode_error_CM_AQM_DCTCP_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_GLOBAL_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h341,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_SHARED_SMP_PAUSE_CFG;
                    ack.write_miss = handcode_error_CM_SHARED_SMP_PAUSE_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_SWEEPER_TC_TO_SMP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_GLOBAL_USAGE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_GLOBAL_USAGE_MAX_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h344,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_MCAST_EPOCH_USAGE;
                    ack.write_miss = handcode_error_CM_MCAST_EPOCH_USAGE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h345,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_SHARED_SMP_USAGE;
                    ack.write_miss = handcode_error_CM_SHARED_SMP_USAGE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h346,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_SMP_USAGE;
                    ack.write_miss = handcode_error_CM_SMP_USAGE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h3,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_RX_SMP_USAGE;
                    ack.write_miss = handcode_error_CM_RX_SMP_USAGE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h38,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_RX_SMP_USAGE_MAX;
                    ack.write_miss = handcode_error_CM_RX_SMP_USAGE_MAX;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h384,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_RX_SMP_USAGE_MAX_CTRL;
                    ack.write_miss = handcode_error_CM_RX_SMP_USAGE_MAX_CTRL;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h39?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_PAUSE_GEN_STATE;
                    ack.write_miss = handcode_error_CM_PAUSE_GEN_STATE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h4??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_TX_TC_USAGE;
                    ack.write_miss = handcode_error_CM_TX_TC_USAGE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h5,4'b00??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_TX_EWMA;
                    ack.write_miss = handcode_error_CM_TX_EWMA;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_CM_USAGE_MAP_MEM) 
           {44'h0??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_TX_TC_PRIVATE_WM;
                 default: read_data = '0;
              endcase
           end
           {44'h1??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_TX_TC_HOG_WM;
                 default: read_data = '0;
              endcase
           end
           {36'h2,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_RX_SMP_PRIVATE_WM;
                 default: read_data = '0;
              endcase
           end
           {36'h2,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_RX_SMP_HOG_WM;
                 default: read_data = '0;
              endcase
           end
           {36'h2,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_RX_SMP_PAUSE_WM;
                 default: read_data = '0;
              endcase
           end
           {40'h26,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_SHARED_WM;
                 default: read_data = '0;
              endcase
           end
           {40'h26,4'b01??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_SOFTDROP_WM;
                 default: read_data = '0;
              endcase
           end
           {44'h268,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_SHARED_SMP_PAUSE_WM;
                 default: read_data = '0;
              endcase
           end
           CM_GLOBAL_WM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = {CM_GLOBAL_WM};
                 default: read_data = '0;
              endcase
           end
           {44'h27?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_PAUSE_PHYS_PORT_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'h280,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_FORCE_PAUSE_CFG;
                 default: read_data = '0;
              endcase
           end
           {36'h2,4'b11??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_AQM_EWMA_CFG;
                 default: read_data = '0;
              endcase
           end
           {36'h3,4'b00??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_AQM_DCTCP_CFG;
                 default: read_data = '0;
              endcase
           end
           CM_GLOBAL_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = {CM_GLOBAL_CFG};
                 default: read_data = '0;
              endcase
           end
           {44'h341,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_SHARED_SMP_PAUSE_CFG;
                 default: read_data = '0;
              endcase
           end
           CM_SWEEPER_TC_TO_SMP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = {CM_SWEEPER_TC_TO_SMP};
                 default: read_data = '0;
              endcase
           end
           CM_GLOBAL_USAGE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = {CM_GLOBAL_USAGE};
                 default: read_data = '0;
              endcase
           end
           CM_GLOBAL_USAGE_MAX_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = {CM_GLOBAL_USAGE_MAX};
                 default: read_data = '0;
              endcase
           end
           {44'h344,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_MCAST_EPOCH_USAGE;
                 default: read_data = '0;
              endcase
           end
           {44'h345,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_SHARED_SMP_USAGE;
                 default: read_data = '0;
              endcase
           end
           {44'h346,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_SMP_USAGE;
                 default: read_data = '0;
              endcase
           end
           {36'h3,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_RX_SMP_USAGE;
                 default: read_data = '0;
              endcase
           end
           {40'h38,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_RX_SMP_USAGE_MAX;
                 default: read_data = '0;
              endcase
           end
           {44'h384,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_RX_SMP_USAGE_MAX_CTRL;
                 default: read_data = '0;
              endcase
           end
           {44'h39?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_PAUSE_GEN_STATE;
                 default: read_data = '0;
              endcase
           end
           {44'h4??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_TX_TC_USAGE;
                 default: read_data = '0;
              endcase
           end
           {36'h5,4'b00??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_USAGE_SB_FID,CM_USAGE_SB_BAR}: read_data = handcode_reg_rdata_CM_TX_EWMA;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    CM_GLOBAL_WM.reserved0 = '0;
    CM_GLOBAL_CFG.reserved0 = '0;
    CM_SWEEPER_TC_TO_SMP.reserved0 = '0;
    CM_GLOBAL_USAGE.reserved0 = '0;
    CM_GLOBAL_USAGE_MAX.reserved0 = '0;
end

// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
