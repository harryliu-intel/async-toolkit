// vim: noai : ts=3 : sw=3 : expandtab : ft=systemverilog

//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors.  The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//   Author        : Kaleem Sheriff
//   Project       : Madison Bay
//------------------------------------------------------------------------------

//   Class:    mby_rx_ppe_env_shutdown_seq
//
//   This is the rx_ppe env Shutdown sequence file.

`ifndef __MBY_RX_PPE_ENV_SHUTDOWN_SEQ_GUARD
`define __MBY_RX_PPE_ENV_SHUTDOWN_SEQ_GUARD

`ifndef __INSIDE_MBY_RX_PPE_SEQ_LIB
`error "Attempt to include file outside of mby_rx_ppe_seq_lib."
`endif

class mby_rx_ppe_env_shutdown_seq extends mby_rx_ppe_env_base_seq;

   `uvm_object_utils(mby_rx_ppe_env_shutdown_seq)

   // Variable: rx_ppe_eot_seq
   // rx_ppe_eot_seq
   mby_rx_ppe_seq_lib::mby_rx_ppe_eot_seq        rx_ppe_eot_seq;

   //------------------------------------------------------------------------------
   //  Constructor: new
   //  
   //  Arguments:
   //  string name  - rx_ppe env shutdown sequence object name.
   //------------------------------------------------------------------------------
   function new(input string name = "mby_rx_ppe_env_shutdown_seq");
      super.new(name);
   endfunction: new

   //------------------------------------------------------------------------------
   //  Task: body
   //  Check rx_ppe DUT.
   //------------------------------------------------------------------------------
   virtual task     body();

      `uvm_info(this.get_name(), ("Phase::shutdown_phase:mby_rx_ppe_env_shutdown_seq::Starting"), UVM_LOW)

//    rx_ppe_eot_seq = mby_rx_ppe_seq_lib::mby_rx_ppe_eot_seq::type_id::create("rx_ppe_eot_seq");
//    rx_ppe_eot_seq.env       = env;
//    rx_ppe_eot_seq.ral_env   = env.tp_env.get_tb_ral();
//    rx_ppe_eot_seq.dut_cfg       = env.tb_cfg.dut_cfg;
//    rx_ppe_eot_seq.access_type  = "FRONTDOOR";
	
      `uvm_info(get_name(), "********** Starting rx_ppe_eot_seq **********", UVM_MEDIUM);
//    rx_ppe_eot_seq.start(sla_sequencer::pick_sequencer("ral_sequencer"));
       
   endtask : body

endclass : mby_rx_ppe_env_shutdown_seq

`endif // __MBY_RX_PPE_ENV_SHUTDOWN_SEQ_GUARD
