magic
tech scmos
timestamp 982685175
<< nselect >>
rect -34 24 0 95
<< pselect >>
rect 0 10 46 103
<< ndiffusion >>
rect -28 81 -8 82
rect -28 73 -8 78
rect -28 65 -8 70
rect -28 57 -8 62
rect -28 49 -8 54
rect -28 41 -8 46
rect -28 37 -8 38
<< pdiffusion >>
rect 14 91 40 92
rect 14 87 40 88
rect 28 79 40 87
rect 14 78 40 79
rect 14 74 40 75
rect 14 65 40 66
rect 14 61 40 62
rect 28 53 40 61
rect 14 52 40 53
rect 14 48 40 49
rect 14 39 40 40
rect 14 35 40 36
rect 14 24 30 27
rect 14 20 30 21
<< ntransistor >>
rect -28 78 -8 81
rect -28 70 -8 73
rect -28 62 -8 65
rect -28 54 -8 57
rect -28 46 -8 49
rect -28 38 -8 41
<< ptransistor >>
rect 14 88 40 91
rect 14 75 40 78
rect 14 62 40 65
rect 14 49 40 52
rect 14 36 40 39
rect 14 21 30 24
<< polysilicon >>
rect -2 88 14 91
rect 40 88 44 91
rect -2 81 1 88
rect -32 78 -28 81
rect -8 78 1 81
rect 9 75 14 78
rect 40 75 44 78
rect 9 73 12 75
rect -32 70 -28 73
rect -8 70 12 73
rect -32 62 -28 65
rect -8 62 14 65
rect 40 62 44 65
rect -32 54 -28 57
rect -8 54 12 57
rect 9 52 12 54
rect 9 49 14 52
rect 40 49 44 52
rect -32 46 -28 49
rect -8 46 4 49
rect -32 38 -28 41
rect -8 38 -4 41
rect 1 39 4 46
rect 1 36 14 39
rect 40 36 44 39
rect 10 21 14 24
rect 30 21 34 24
<< ndcontact >>
rect -28 82 -8 90
rect -28 29 -8 37
<< pdcontact >>
rect 14 92 40 100
rect 14 79 28 87
rect 14 66 40 74
rect 14 53 28 61
rect 14 40 40 48
rect 14 27 40 35
rect 14 12 30 20
<< metal1 >>
rect 14 99 40 100
rect 27 93 40 99
rect 14 92 40 93
rect -28 87 5 90
rect -28 82 28 87
rect -3 79 28 82
rect -3 61 5 79
rect 32 74 40 92
rect 14 66 40 74
rect -3 53 28 61
rect -28 29 -8 37
rect -3 35 5 53
rect 32 48 40 66
rect 27 42 40 48
rect 14 40 40 42
rect -27 18 -9 29
rect -3 27 40 35
rect 14 18 30 20
rect 27 12 30 18
<< m2contact >>
rect 9 93 27 99
rect 9 42 27 48
rect -27 12 -9 18
rect 9 12 27 18
<< m3contact >>
rect 9 93 27 99
rect 9 42 27 48
rect -27 12 -9 18
rect 9 12 27 18
<< metal3 >>
rect -27 10 -9 103
rect 9 10 27 103
<< labels >>
rlabel space -35 23 -28 96 7 ^n
rlabel space 28 31 47 103 3 ^p
rlabel metal3 -27 10 -9 103 1 GND!|pin|s|0
rlabel metal1 -28 29 -8 37 1 GND!|pin|s|0
rlabel metal1 -27 12 -9 37 1 GND!|pin|s|0
rlabel metal3 9 10 27 103 1 Vdd!|pin|s|1
rlabel metal1 14 92 40 100 1 Vdd!|pin|s|1
rlabel metal1 14 66 40 74 1 Vdd!|pin|s|1
rlabel metal1 14 40 40 48 1 Vdd!|pin|s|1
rlabel metal1 32 40 40 100 1 Vdd!|pin|s|1
rlabel metal1 -3 27 5 90 1 x|pin|s|2
rlabel metal1 -28 82 5 90 1 x|pin|s|2
rlabel metal1 -3 79 28 87 1 x|pin|s|2
rlabel metal1 -3 53 28 61 1 x|pin|s|2
rlabel metal1 -3 27 40 35 1 x|pin|s|2
rlabel polysilicon 40 36 44 39 1 a|pin|w|3|poly
rlabel polysilicon 1 36 5 39 1 a|pin|w|3|poly
rlabel polysilicon -32 46 -28 49 1 a|pin|w|3|poly
rlabel polysilicon 40 49 44 52 1 b|pin|w|4|poly
rlabel polysilicon -32 54 -28 57 1 b|pin|w|4|poly
rlabel polysilicon 40 62 44 65 1 c|pin|w|5|poly
rlabel polysilicon -32 62 -28 65 1 c|pin|w|5|poly
rlabel polysilicon 40 75 44 78 1 d|pin|w|6|poly
rlabel polysilicon -32 70 -28 73 1 d|pin|w|6|poly
rlabel polysilicon 40 88 44 91 1 e|pin|w|7|poly
rlabel polysilicon -2 88 2 91 1 e|pin|w|7|poly
rlabel polysilicon -32 78 -28 81 1 e|pin|w|7|poly
rlabel polysilicon -32 38 -28 41 1 _SReset!|pin|w|8|poly
rlabel polysilicon -8 38 -4 41 1 _SReset!|pin|w|8|poly
rlabel polysilicon 10 21 14 24 1 _PReset!|pin|w|9|poly
rlabel polysilicon 30 21 34 24 1 _PReset!|pin|w|9|poly
rlabel metal1 14 12 30 20 1 Vdd!|pin|s|1
<< end >>
