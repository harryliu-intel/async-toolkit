///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_entropy_map.sv                                     
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_entropy_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_FF
`define RTLGEN_MBY_PPE_ENTROPY_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_FF

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF
`define RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_ENTROPY_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_FF_RSTD


module rtlgen_mby_ppe_entropy_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_entropy_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_ENTROPY_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_ENTROPY_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_ENTROPY_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_PH2_FF
`define RTLGEN_MBY_PPE_ENTROPY_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_ENTROPY_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_ENTROPY_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH
`define RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_ENTROPY_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_ENTROPY_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_entropy_map ( //lintra s-2096
    // Clocks
    gated_clk,

    // Resets
    rst_n,


    // Register Inputs
    handcode_reg_rdata_ENTROPY_HASH_CFG0,
    handcode_reg_rdata_ENTROPY_HASH_CFG1,
    handcode_reg_rdata_ENTROPY_HASH_KEY_MASK,
    handcode_reg_rdata_ENTROPY_HASH_SYM16,
    handcode_reg_rdata_ENTROPY_HASH_SYM32,
    handcode_reg_rdata_ENTROPY_HASH_SYM8,
    handcode_reg_rdata_ENTROPY_META_CFG,

    handcode_rvalid_ENTROPY_HASH_CFG0,
    handcode_rvalid_ENTROPY_HASH_CFG1,
    handcode_rvalid_ENTROPY_HASH_KEY_MASK,
    handcode_rvalid_ENTROPY_HASH_SYM16,
    handcode_rvalid_ENTROPY_HASH_SYM32,
    handcode_rvalid_ENTROPY_HASH_SYM8,
    handcode_rvalid_ENTROPY_META_CFG,

    handcode_wvalid_ENTROPY_HASH_CFG0,
    handcode_wvalid_ENTROPY_HASH_CFG1,
    handcode_wvalid_ENTROPY_HASH_KEY_MASK,
    handcode_wvalid_ENTROPY_HASH_SYM16,
    handcode_wvalid_ENTROPY_HASH_SYM32,
    handcode_wvalid_ENTROPY_HASH_SYM8,
    handcode_wvalid_ENTROPY_META_CFG,

    handcode_error_ENTROPY_HASH_CFG0,
    handcode_error_ENTROPY_HASH_CFG1,
    handcode_error_ENTROPY_HASH_KEY_MASK,
    handcode_error_ENTROPY_HASH_SYM16,
    handcode_error_ENTROPY_HASH_SYM32,
    handcode_error_ENTROPY_HASH_SYM8,
    handcode_error_ENTROPY_META_CFG,


    // Register Outputs
    ENTROPY_FWD_HASHING_CFG,


    // Register signals for HandCoded registers
    handcode_reg_wdata_ENTROPY_HASH_CFG0,
    handcode_reg_wdata_ENTROPY_HASH_CFG1,
    handcode_reg_wdata_ENTROPY_HASH_KEY_MASK,
    handcode_reg_wdata_ENTROPY_HASH_SYM16,
    handcode_reg_wdata_ENTROPY_HASH_SYM32,
    handcode_reg_wdata_ENTROPY_HASH_SYM8,
    handcode_reg_wdata_ENTROPY_META_CFG,

    we_ENTROPY_HASH_CFG0,
    we_ENTROPY_HASH_CFG1,
    we_ENTROPY_HASH_KEY_MASK,
    we_ENTROPY_HASH_SYM16,
    we_ENTROPY_HASH_SYM32,
    we_ENTROPY_HASH_SYM8,
    we_ENTROPY_META_CFG,

    re_ENTROPY_HASH_CFG0,
    re_ENTROPY_HASH_CFG1,
    re_ENTROPY_HASH_KEY_MASK,
    re_ENTROPY_HASH_SYM16,
    re_ENTROPY_HASH_SYM32,
    re_ENTROPY_HASH_SYM8,
    re_ENTROPY_META_CFG,




    // Config Access
    req,
    ack
    

);

import mby_ppe_entropy_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:0] MBY_PPE_ENTROPY_MAP_OFFSET = {MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] ENTROPY_SB_BAR = 3'b0;
parameter [7:0] ENTROPY_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
`define ENTROPY_FWD_HASHING_CFG_CR_ADDR_def(INDEX) ENTROPY_FWD_HASHING_CFG_CR_ADDR``INDEX``[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_ENTROPY_MAP_OFFSET[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
localparam [63:0][MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] ENTROPY_FWD_HASHING_CFG_DECODE_ADDR = {`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([63]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([62]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([61]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([60]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([59]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([58]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([57]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([56]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([55]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([54]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([53]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([52]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([51]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([50]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([49]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([48]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([47]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([46]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([45]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([44]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([43]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([42]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([41]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([40]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([39]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([38]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([37]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([36]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([35]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([34]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([33]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([32]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([31]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([30]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([29]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([28]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([27]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([26]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([25]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([24]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([23]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([22]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([21]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([20]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([19]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([18]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([17]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([16]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([15]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([14]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([13]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([12]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([11]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([10]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([9]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([8]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([7]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([6]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([5]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([4]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([3]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([2]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([1]),`ENTROPY_FWD_HASHING_CFG_CR_ADDR_def([0])};

    // Clocks
input logic  gated_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input ENTROPY_HASH_CFG0_t  handcode_reg_rdata_ENTROPY_HASH_CFG0;
input ENTROPY_HASH_CFG1_t  handcode_reg_rdata_ENTROPY_HASH_CFG1;
input ENTROPY_HASH_KEY_MASK_t  handcode_reg_rdata_ENTROPY_HASH_KEY_MASK;
input ENTROPY_HASH_SYM16_t  handcode_reg_rdata_ENTROPY_HASH_SYM16;
input ENTROPY_HASH_SYM32_t  handcode_reg_rdata_ENTROPY_HASH_SYM32;
input ENTROPY_HASH_SYM8_t  handcode_reg_rdata_ENTROPY_HASH_SYM8;
input ENTROPY_META_CFG_t  handcode_reg_rdata_ENTROPY_META_CFG;

input handcode_rvalid_ENTROPY_HASH_CFG0_t  handcode_rvalid_ENTROPY_HASH_CFG0;
input handcode_rvalid_ENTROPY_HASH_CFG1_t  handcode_rvalid_ENTROPY_HASH_CFG1;
input handcode_rvalid_ENTROPY_HASH_KEY_MASK_t  handcode_rvalid_ENTROPY_HASH_KEY_MASK;
input handcode_rvalid_ENTROPY_HASH_SYM16_t  handcode_rvalid_ENTROPY_HASH_SYM16;
input handcode_rvalid_ENTROPY_HASH_SYM32_t  handcode_rvalid_ENTROPY_HASH_SYM32;
input handcode_rvalid_ENTROPY_HASH_SYM8_t  handcode_rvalid_ENTROPY_HASH_SYM8;
input handcode_rvalid_ENTROPY_META_CFG_t  handcode_rvalid_ENTROPY_META_CFG;

input handcode_wvalid_ENTROPY_HASH_CFG0_t  handcode_wvalid_ENTROPY_HASH_CFG0;
input handcode_wvalid_ENTROPY_HASH_CFG1_t  handcode_wvalid_ENTROPY_HASH_CFG1;
input handcode_wvalid_ENTROPY_HASH_KEY_MASK_t  handcode_wvalid_ENTROPY_HASH_KEY_MASK;
input handcode_wvalid_ENTROPY_HASH_SYM16_t  handcode_wvalid_ENTROPY_HASH_SYM16;
input handcode_wvalid_ENTROPY_HASH_SYM32_t  handcode_wvalid_ENTROPY_HASH_SYM32;
input handcode_wvalid_ENTROPY_HASH_SYM8_t  handcode_wvalid_ENTROPY_HASH_SYM8;
input handcode_wvalid_ENTROPY_META_CFG_t  handcode_wvalid_ENTROPY_META_CFG;

input handcode_error_ENTROPY_HASH_CFG0_t  handcode_error_ENTROPY_HASH_CFG0;
input handcode_error_ENTROPY_HASH_CFG1_t  handcode_error_ENTROPY_HASH_CFG1;
input handcode_error_ENTROPY_HASH_KEY_MASK_t  handcode_error_ENTROPY_HASH_KEY_MASK;
input handcode_error_ENTROPY_HASH_SYM16_t  handcode_error_ENTROPY_HASH_SYM16;
input handcode_error_ENTROPY_HASH_SYM32_t  handcode_error_ENTROPY_HASH_SYM32;
input handcode_error_ENTROPY_HASH_SYM8_t  handcode_error_ENTROPY_HASH_SYM8;
input handcode_error_ENTROPY_META_CFG_t  handcode_error_ENTROPY_META_CFG;


    // Register Outputs
output ENTROPY_FWD_HASHING_CFG_t [63:0] ENTROPY_FWD_HASHING_CFG;


    // Register signals for HandCoded registers
output ENTROPY_HASH_CFG0_t  handcode_reg_wdata_ENTROPY_HASH_CFG0;
output ENTROPY_HASH_CFG1_t  handcode_reg_wdata_ENTROPY_HASH_CFG1;
output ENTROPY_HASH_KEY_MASK_t  handcode_reg_wdata_ENTROPY_HASH_KEY_MASK;
output ENTROPY_HASH_SYM16_t  handcode_reg_wdata_ENTROPY_HASH_SYM16;
output ENTROPY_HASH_SYM32_t  handcode_reg_wdata_ENTROPY_HASH_SYM32;
output ENTROPY_HASH_SYM8_t  handcode_reg_wdata_ENTROPY_HASH_SYM8;
output ENTROPY_META_CFG_t  handcode_reg_wdata_ENTROPY_META_CFG;

output we_ENTROPY_HASH_CFG0_t  we_ENTROPY_HASH_CFG0;
output we_ENTROPY_HASH_CFG1_t  we_ENTROPY_HASH_CFG1;
output we_ENTROPY_HASH_KEY_MASK_t  we_ENTROPY_HASH_KEY_MASK;
output we_ENTROPY_HASH_SYM16_t  we_ENTROPY_HASH_SYM16;
output we_ENTROPY_HASH_SYM32_t  we_ENTROPY_HASH_SYM32;
output we_ENTROPY_HASH_SYM8_t  we_ENTROPY_HASH_SYM8;
output we_ENTROPY_META_CFG_t  we_ENTROPY_META_CFG;

output re_ENTROPY_HASH_CFG0_t  re_ENTROPY_HASH_CFG0;
output re_ENTROPY_HASH_CFG1_t  re_ENTROPY_HASH_CFG1;
output re_ENTROPY_HASH_KEY_MASK_t  re_ENTROPY_HASH_KEY_MASK;
output re_ENTROPY_HASH_SYM16_t  re_ENTROPY_HASH_SYM16;
output re_ENTROPY_HASH_SYM32_t  re_ENTROPY_HASH_SYM32;
output re_ENTROPY_HASH_SYM8_t  re_ENTROPY_HASH_SYM8;
output re_ENTROPY_META_CFG_t  re_ENTROPY_META_CFG;




    // Config Access
input mby_ppe_entropy_map_cr_req_t  req;
output mby_ppe_entropy_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_entropy_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_ENTROPY_MAP_MEM;
assign case_req_addr_MBY_PPE_ENTROPY_MAP_MEM = req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_entropy;
always_comb begin : sb_fid_cond_entropy_BLOCK
    unique casez (req_fid) 
		ENTROPY_SB_FID: sb_fid_cond_entropy = 1;
		default: sb_fid_cond_entropy = 0;
    endcase 
end


logic sb_bar_cond_entropy;
always_comb begin : sb_bar_cond_entropy_BLOCK
    unique casez (req_bar) 
		ENTROPY_SB_BAR: sb_bar_cond_entropy = 1;
		default: sb_bar_cond_entropy = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// ENTROPY_HASH_CFG0 using HANDCODED_REG template.
logic addr_decode_ENTROPY_HASH_CFG0;
logic write_req_ENTROPY_HASH_CFG0;
logic read_req_ENTROPY_HASH_CFG0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b0??,4'h?,1'b?},
      {40'b10?,4'h?,1'b?}:
          addr_decode_ENTROPY_HASH_CFG0 = req.valid;
      default: 
         addr_decode_ENTROPY_HASH_CFG0 = 1'b0; 
   endcase
end

always_comb write_req_ENTROPY_HASH_CFG0 = f_IsMEMWr(req_opcode) && addr_decode_ENTROPY_HASH_CFG0 ;
always_comb read_req_ENTROPY_HASH_CFG0  = f_IsMEMRd(req_opcode) && addr_decode_ENTROPY_HASH_CFG0 ;

always_comb we_ENTROPY_HASH_CFG0 = {8{write_req_ENTROPY_HASH_CFG0}} & be;
always_comb re_ENTROPY_HASH_CFG0 = {8{read_req_ENTROPY_HASH_CFG0}} & be;
always_comb handcode_reg_wdata_ENTROPY_HASH_CFG0 = write_data;


// ----------------------------------------------------------------------
// ENTROPY_HASH_CFG1 using HANDCODED_REG template.
logic addr_decode_ENTROPY_HASH_CFG1;
logic write_req_ENTROPY_HASH_CFG1;
logic read_req_ENTROPY_HASH_CFG1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b10??,4'h?,1'b?},
      {40'b110?,4'h?,1'b?}:
          addr_decode_ENTROPY_HASH_CFG1 = req.valid;
      default: 
         addr_decode_ENTROPY_HASH_CFG1 = 1'b0; 
   endcase
end

always_comb write_req_ENTROPY_HASH_CFG1 = f_IsMEMWr(req_opcode) && addr_decode_ENTROPY_HASH_CFG1 ;
always_comb read_req_ENTROPY_HASH_CFG1  = f_IsMEMRd(req_opcode) && addr_decode_ENTROPY_HASH_CFG1 ;

always_comb we_ENTROPY_HASH_CFG1 = {8{write_req_ENTROPY_HASH_CFG1}} & be;
always_comb re_ENTROPY_HASH_CFG1 = {8{read_req_ENTROPY_HASH_CFG1}} & be;
always_comb handcode_reg_wdata_ENTROPY_HASH_CFG1 = write_data;


// ----------------------------------------------------------------------
// ENTROPY_META_CFG using HANDCODED_REG template.
logic addr_decode_ENTROPY_META_CFG;
logic write_req_ENTROPY_META_CFG;
logic read_req_ENTROPY_META_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b111?,4'h?,1'b?}: 
         addr_decode_ENTROPY_META_CFG = req.valid;
      default: 
         addr_decode_ENTROPY_META_CFG = 1'b0; 
   endcase
end

always_comb write_req_ENTROPY_META_CFG = f_IsMEMWr(req_opcode) && addr_decode_ENTROPY_META_CFG ;
always_comb read_req_ENTROPY_META_CFG  = f_IsMEMRd(req_opcode) && addr_decode_ENTROPY_META_CFG ;

always_comb we_ENTROPY_META_CFG = {8{write_req_ENTROPY_META_CFG}} & be;
always_comb re_ENTROPY_META_CFG = {8{read_req_ENTROPY_META_CFG}} & be;
always_comb handcode_reg_wdata_ENTROPY_META_CFG = write_data;


// ----------------------------------------------------------------------
// ENTROPY_HASH_SYM8 using HANDCODED_REG template.
logic addr_decode_ENTROPY_HASH_SYM8;
logic write_req_ENTROPY_HASH_SYM8;
logic read_req_ENTROPY_HASH_SYM8;

always_comb begin 
   unique casez (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h10,4'b00??,1'b?},
      {40'h10,4'b010?,1'b?}:
          addr_decode_ENTROPY_HASH_SYM8 = req.valid;
      default: 
         addr_decode_ENTROPY_HASH_SYM8 = 1'b0; 
   endcase
end

always_comb write_req_ENTROPY_HASH_SYM8 = f_IsMEMWr(req_opcode) && addr_decode_ENTROPY_HASH_SYM8 ;
always_comb read_req_ENTROPY_HASH_SYM8  = f_IsMEMRd(req_opcode) && addr_decode_ENTROPY_HASH_SYM8 ;

always_comb we_ENTROPY_HASH_SYM8 = {8{write_req_ENTROPY_HASH_SYM8}} & be;
always_comb re_ENTROPY_HASH_SYM8 = {8{read_req_ENTROPY_HASH_SYM8}} & be;
always_comb handcode_reg_wdata_ENTROPY_HASH_SYM8 = write_data;


// ----------------------------------------------------------------------
// ENTROPY_HASH_SYM16 using HANDCODED_REG template.
logic addr_decode_ENTROPY_HASH_SYM16;
logic write_req_ENTROPY_HASH_SYM16;
logic read_req_ENTROPY_HASH_SYM16;

always_comb begin 
   unique casez (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h10,4'b10??,1'b?},
      {40'h10,4'b110?,1'b?}:
          addr_decode_ENTROPY_HASH_SYM16 = req.valid;
      default: 
         addr_decode_ENTROPY_HASH_SYM16 = 1'b0; 
   endcase
end

always_comb write_req_ENTROPY_HASH_SYM16 = f_IsMEMWr(req_opcode) && addr_decode_ENTROPY_HASH_SYM16 ;
always_comb read_req_ENTROPY_HASH_SYM16  = f_IsMEMRd(req_opcode) && addr_decode_ENTROPY_HASH_SYM16 ;

always_comb we_ENTROPY_HASH_SYM16 = {8{write_req_ENTROPY_HASH_SYM16}} & be;
always_comb re_ENTROPY_HASH_SYM16 = {8{read_req_ENTROPY_HASH_SYM16}} & be;
always_comb handcode_reg_wdata_ENTROPY_HASH_SYM16 = write_data;


// ----------------------------------------------------------------------
// ENTROPY_HASH_SYM32 using HANDCODED_REG template.
logic addr_decode_ENTROPY_HASH_SYM32;
logic write_req_ENTROPY_HASH_SYM32;
logic read_req_ENTROPY_HASH_SYM32;

always_comb begin 
   unique casez (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h11,4'b00??,1'b?},
      {40'h11,4'b010?,1'b?}:
          addr_decode_ENTROPY_HASH_SYM32 = req.valid;
      default: 
         addr_decode_ENTROPY_HASH_SYM32 = 1'b0; 
   endcase
end

always_comb write_req_ENTROPY_HASH_SYM32 = f_IsMEMWr(req_opcode) && addr_decode_ENTROPY_HASH_SYM32 ;
always_comb read_req_ENTROPY_HASH_SYM32  = f_IsMEMRd(req_opcode) && addr_decode_ENTROPY_HASH_SYM32 ;

always_comb we_ENTROPY_HASH_SYM32 = {8{write_req_ENTROPY_HASH_SYM32}} & be;
always_comb re_ENTROPY_HASH_SYM32 = {8{read_req_ENTROPY_HASH_SYM32}} & be;
always_comb handcode_reg_wdata_ENTROPY_HASH_SYM32 = write_data;


// ----------------------------------------------------------------------
// ENTROPY_HASH_KEY_MASK using HANDCODED_REG template.
logic addr_decode_ENTROPY_HASH_KEY_MASK;
logic write_req_ENTROPY_HASH_KEY_MASK;
logic read_req_ENTROPY_HASH_KEY_MASK;

always_comb begin 
   unique casez (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h2,4'b0???,4'h?,1'b?},
      {36'h2,4'b10??,4'h?,1'b?}:
          addr_decode_ENTROPY_HASH_KEY_MASK = req.valid;
      default: 
         addr_decode_ENTROPY_HASH_KEY_MASK = 1'b0; 
   endcase
end

always_comb write_req_ENTROPY_HASH_KEY_MASK = f_IsMEMWr(req_opcode) && addr_decode_ENTROPY_HASH_KEY_MASK ;
always_comb read_req_ENTROPY_HASH_KEY_MASK  = f_IsMEMRd(req_opcode) && addr_decode_ENTROPY_HASH_KEY_MASK ;

always_comb we_ENTROPY_HASH_KEY_MASK = {8{write_req_ENTROPY_HASH_KEY_MASK}} & be;
always_comb re_ENTROPY_HASH_KEY_MASK = {8{read_req_ENTROPY_HASH_KEY_MASK}} & be;
always_comb handcode_reg_wdata_ENTROPY_HASH_KEY_MASK = write_data;


//---------------------------------------------------------------------
// ENTROPY_FWD_HASHING_CFG Address Decode
logic [63:0] addr_decode_ENTROPY_FWD_HASHING_CFG;
logic [63:0] write_req_ENTROPY_FWD_HASHING_CFG;
always_comb begin
   addr_decode_ENTROPY_FWD_HASHING_CFG[0] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[0]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[1] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[1]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[2] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[2]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[3] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[3]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[4] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[4]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[5] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[5]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[6] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[6]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[7] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[7]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[8] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[8]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[9] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[9]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[10] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[10]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[11] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[11]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[12] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[12]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[13] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[13]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[14] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[14]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[15] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[15]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[16] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[16]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[17] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[17]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[18] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[18]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[19] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[19]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[20] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[20]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[21] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[21]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[22] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[22]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[23] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[23]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[24] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[24]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[25] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[25]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[26] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[26]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[27] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[27]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[28] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[28]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[29] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[29]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[30] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[30]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[31] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[31]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[32] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[32]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[33] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[33]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[34] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[34]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[35] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[35]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[36] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[36]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[37] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[37]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[38] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[38]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[39] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[39]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[40] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[40]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[41] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[41]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[42] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[42]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[43] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[43]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[44] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[44]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[45] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[45]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[46] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[46]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[47] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[47]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[48] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[48]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[49] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[49]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[50] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[50]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[51] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[51]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[52] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[52]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[53] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[53]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[54] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[54]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[55] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[55]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[56] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[56]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[57] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[57]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[58] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[58]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[59] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[59]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[60] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[60]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[61] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[61]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[62] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[62]) && req.valid ;
   addr_decode_ENTROPY_FWD_HASHING_CFG[63] = (req_addr[MBY_PPE_ENTROPY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[63]) && req.valid ;
   write_req_ENTROPY_FWD_HASHING_CFG[0] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[0] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[1] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[1] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[2] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[2] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[3] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[3] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[4] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[4] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[5] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[5] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[6] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[6] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[7] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[7] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[8] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[8] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[9] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[9] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[10] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[10] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[11] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[11] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[12] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[12] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[13] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[13] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[14] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[14] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[15] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[15] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[16] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[16] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[17] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[17] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[18] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[18] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[19] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[19] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[20] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[20] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[21] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[21] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[22] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[22] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[23] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[23] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[24] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[24] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[25] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[25] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[26] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[26] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[27] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[27] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[28] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[28] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[29] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[29] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[30] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[30] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[31] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[31] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[32] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[32] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[33] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[33] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[34] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[34] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[35] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[35] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[36] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[36] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[37] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[37] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[38] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[38] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[39] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[39] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[40] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[40] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[41] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[41] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[42] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[42] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[43] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[43] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[44] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[44] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[45] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[45] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[46] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[46] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[47] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[47] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[48] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[48] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[49] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[49] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[50] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[50] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[51] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[51] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[52] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[52] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[53] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[53] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[54] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[54] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[55] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[55] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[56] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[56] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[57] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[57] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[58] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[58] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[59] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[59] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[60] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[60] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[61] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[61] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[62] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[62] && sb_fid_cond_entropy && sb_bar_cond_entropy;
   write_req_ENTROPY_FWD_HASHING_CFG[63] = IsMEMWr && addr_decode_ENTROPY_FWD_HASHING_CFG[63] && sb_fid_cond_entropy && sb_bar_cond_entropy;
end


// ----------------------------------------------------------------------
// ENTROPY_FWD_HASHING_CFG.ROTATION_A x2 RW, using RW template.
logic [63:0][0:0] up_ENTROPY_FWD_HASHING_CFG_ROTATION_A;
always_comb begin
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[0] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[0] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[1] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[1] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[2] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[2] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[3] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[3] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[4] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[4] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[5] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[5] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[6] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[6] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[7] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[7] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[8] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[8] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[9] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[9] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[10] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[10] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[11] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[11] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[12] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[12] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[13] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[13] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[14] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[14] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[15] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[15] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[16] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[16] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[17] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[17] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[18] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[18] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[19] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[19] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[20] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[20] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[21] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[21] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[22] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[22] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[23] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[23] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[24] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[24] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[25] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[25] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[26] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[26] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[27] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[27] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[28] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[28] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[29] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[29] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[30] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[30] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[31] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[31] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[32] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[32] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[33] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[33] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[34] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[34] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[35] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[35] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[36] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[36] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[37] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[37] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[38] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[38] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[39] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[39] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[40] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[40] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[41] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[41] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[42] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[42] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[43] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[43] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[44] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[44] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[45] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[45] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[46] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[46] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[47] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[47] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[48] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[48] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[49] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[49] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[50] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[50] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[51] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[51] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[52] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[52] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[53] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[53] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[54] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[54] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[55] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[55] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[56] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[56] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[57] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[57] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[58] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[58] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[59] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[59] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[60] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[60] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[61] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[61] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[62] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[62] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[63] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[63] }} &
    be[1:1]);
end

logic [63:0][1:0] nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A;
always_comb begin
 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[0] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[1] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[2] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[3] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[4] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[5] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[6] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[7] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[8] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[9] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[10] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[11] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[12] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[13] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[14] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[15] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[16] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[17] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[18] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[19] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[20] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[21] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[22] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[23] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[24] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[25] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[26] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[27] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[28] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[29] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[30] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[31] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[32] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[33] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[34] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[35] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[36] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[37] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[38] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[39] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[40] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[41] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[42] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[43] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[44] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[45] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[46] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[47] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[48] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[49] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[50] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[51] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[52] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[53] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[54] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[55] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[56] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[57] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[58] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[59] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[60] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[61] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[62] = write_data[9:8];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[63] = write_data[9:8];

end


`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[0][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[0][1:0], ENTROPY_FWD_HASHING_CFG[0].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[1][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[1][1:0], ENTROPY_FWD_HASHING_CFG[1].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[2][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[2][1:0], ENTROPY_FWD_HASHING_CFG[2].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[3][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[3][1:0], ENTROPY_FWD_HASHING_CFG[3].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[4][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[4][1:0], ENTROPY_FWD_HASHING_CFG[4].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[5][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[5][1:0], ENTROPY_FWD_HASHING_CFG[5].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[6][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[6][1:0], ENTROPY_FWD_HASHING_CFG[6].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[7][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[7][1:0], ENTROPY_FWD_HASHING_CFG[7].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[8][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[8][1:0], ENTROPY_FWD_HASHING_CFG[8].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[9][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[9][1:0], ENTROPY_FWD_HASHING_CFG[9].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[10][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[10][1:0], ENTROPY_FWD_HASHING_CFG[10].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[11][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[11][1:0], ENTROPY_FWD_HASHING_CFG[11].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[12][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[12][1:0], ENTROPY_FWD_HASHING_CFG[12].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[13][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[13][1:0], ENTROPY_FWD_HASHING_CFG[13].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[14][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[14][1:0], ENTROPY_FWD_HASHING_CFG[14].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[15][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[15][1:0], ENTROPY_FWD_HASHING_CFG[15].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[16][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[16][1:0], ENTROPY_FWD_HASHING_CFG[16].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[17][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[17][1:0], ENTROPY_FWD_HASHING_CFG[17].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[18][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[18][1:0], ENTROPY_FWD_HASHING_CFG[18].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[19][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[19][1:0], ENTROPY_FWD_HASHING_CFG[19].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[20][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[20][1:0], ENTROPY_FWD_HASHING_CFG[20].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[21][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[21][1:0], ENTROPY_FWD_HASHING_CFG[21].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[22][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[22][1:0], ENTROPY_FWD_HASHING_CFG[22].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[23][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[23][1:0], ENTROPY_FWD_HASHING_CFG[23].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[24][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[24][1:0], ENTROPY_FWD_HASHING_CFG[24].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[25][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[25][1:0], ENTROPY_FWD_HASHING_CFG[25].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[26][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[26][1:0], ENTROPY_FWD_HASHING_CFG[26].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[27][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[27][1:0], ENTROPY_FWD_HASHING_CFG[27].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[28][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[28][1:0], ENTROPY_FWD_HASHING_CFG[28].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[29][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[29][1:0], ENTROPY_FWD_HASHING_CFG[29].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[30][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[30][1:0], ENTROPY_FWD_HASHING_CFG[30].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[31][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[31][1:0], ENTROPY_FWD_HASHING_CFG[31].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[32][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[32][1:0], ENTROPY_FWD_HASHING_CFG[32].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[33][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[33][1:0], ENTROPY_FWD_HASHING_CFG[33].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[34][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[34][1:0], ENTROPY_FWD_HASHING_CFG[34].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[35][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[35][1:0], ENTROPY_FWD_HASHING_CFG[35].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[36][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[36][1:0], ENTROPY_FWD_HASHING_CFG[36].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[37][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[37][1:0], ENTROPY_FWD_HASHING_CFG[37].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[38][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[38][1:0], ENTROPY_FWD_HASHING_CFG[38].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[39][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[39][1:0], ENTROPY_FWD_HASHING_CFG[39].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[40][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[40][1:0], ENTROPY_FWD_HASHING_CFG[40].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[41][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[41][1:0], ENTROPY_FWD_HASHING_CFG[41].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[42][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[42][1:0], ENTROPY_FWD_HASHING_CFG[42].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[43][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[43][1:0], ENTROPY_FWD_HASHING_CFG[43].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[44][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[44][1:0], ENTROPY_FWD_HASHING_CFG[44].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[45][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[45][1:0], ENTROPY_FWD_HASHING_CFG[45].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[46][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[46][1:0], ENTROPY_FWD_HASHING_CFG[46].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[47][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[47][1:0], ENTROPY_FWD_HASHING_CFG[47].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[48][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[48][1:0], ENTROPY_FWD_HASHING_CFG[48].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[49][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[49][1:0], ENTROPY_FWD_HASHING_CFG[49].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[50][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[50][1:0], ENTROPY_FWD_HASHING_CFG[50].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[51][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[51][1:0], ENTROPY_FWD_HASHING_CFG[51].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[52][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[52][1:0], ENTROPY_FWD_HASHING_CFG[52].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[53][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[53][1:0], ENTROPY_FWD_HASHING_CFG[53].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[54][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[54][1:0], ENTROPY_FWD_HASHING_CFG[54].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[55][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[55][1:0], ENTROPY_FWD_HASHING_CFG[55].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[56][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[56][1:0], ENTROPY_FWD_HASHING_CFG[56].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[57][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[57][1:0], ENTROPY_FWD_HASHING_CFG[57].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[58][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[58][1:0], ENTROPY_FWD_HASHING_CFG[58].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[59][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[59][1:0], ENTROPY_FWD_HASHING_CFG[59].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[60][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[60][1:0], ENTROPY_FWD_HASHING_CFG[60].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[61][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[61][1:0], ENTROPY_FWD_HASHING_CFG[61].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[62][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[62][1:0], ENTROPY_FWD_HASHING_CFG[62].ROTATION_A[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_ENTROPY_FWD_HASHING_CFG_ROTATION_A[63][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_A[63][1:0], ENTROPY_FWD_HASHING_CFG[63].ROTATION_A[1:0])

// ----------------------------------------------------------------------
// ENTROPY_FWD_HASHING_CFG.ROTATION_B x2 RW, using RW template.
logic [63:0][0:0] up_ENTROPY_FWD_HASHING_CFG_ROTATION_B;
always_comb begin
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[0] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[0] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[1] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[1] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[2] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[2] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[3] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[3] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[4] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[4] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[5] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[5] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[6] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[6] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[7] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[7] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[8] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[8] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[9] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[9] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[10] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[10] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[11] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[11] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[12] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[12] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[13] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[13] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[14] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[14] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[15] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[15] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[16] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[16] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[17] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[17] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[18] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[18] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[19] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[19] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[20] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[20] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[21] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[21] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[22] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[22] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[23] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[23] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[24] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[24] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[25] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[25] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[26] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[26] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[27] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[27] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[28] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[28] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[29] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[29] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[30] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[30] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[31] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[31] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[32] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[32] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[33] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[33] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[34] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[34] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[35] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[35] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[36] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[36] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[37] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[37] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[38] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[38] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[39] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[39] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[40] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[40] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[41] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[41] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[42] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[42] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[43] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[43] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[44] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[44] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[45] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[45] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[46] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[46] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[47] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[47] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[48] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[48] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[49] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[49] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[50] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[50] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[51] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[51] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[52] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[52] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[53] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[53] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[54] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[54] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[55] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[55] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[56] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[56] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[57] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[57] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[58] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[58] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[59] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[59] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[60] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[60] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[61] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[61] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[62] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[62] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[63] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[63] }} &
    be[1:1]);
end

logic [63:0][1:0] nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B;
always_comb begin
 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[0] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[1] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[2] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[3] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[4] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[5] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[6] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[7] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[8] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[9] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[10] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[11] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[12] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[13] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[14] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[15] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[16] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[17] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[18] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[19] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[20] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[21] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[22] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[23] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[24] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[25] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[26] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[27] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[28] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[29] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[30] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[31] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[32] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[33] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[34] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[35] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[36] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[37] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[38] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[39] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[40] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[41] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[42] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[43] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[44] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[45] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[46] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[47] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[48] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[49] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[50] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[51] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[52] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[53] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[54] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[55] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[56] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[57] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[58] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[59] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[60] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[61] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[62] = write_data[11:10];

 nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[63] = write_data[11:10];

end


`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[0][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[0][1:0], ENTROPY_FWD_HASHING_CFG[0].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[1][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[1][1:0], ENTROPY_FWD_HASHING_CFG[1].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[2][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[2][1:0], ENTROPY_FWD_HASHING_CFG[2].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[3][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[3][1:0], ENTROPY_FWD_HASHING_CFG[3].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[4][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[4][1:0], ENTROPY_FWD_HASHING_CFG[4].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[5][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[5][1:0], ENTROPY_FWD_HASHING_CFG[5].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[6][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[6][1:0], ENTROPY_FWD_HASHING_CFG[6].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[7][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[7][1:0], ENTROPY_FWD_HASHING_CFG[7].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[8][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[8][1:0], ENTROPY_FWD_HASHING_CFG[8].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[9][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[9][1:0], ENTROPY_FWD_HASHING_CFG[9].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[10][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[10][1:0], ENTROPY_FWD_HASHING_CFG[10].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[11][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[11][1:0], ENTROPY_FWD_HASHING_CFG[11].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[12][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[12][1:0], ENTROPY_FWD_HASHING_CFG[12].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[13][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[13][1:0], ENTROPY_FWD_HASHING_CFG[13].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[14][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[14][1:0], ENTROPY_FWD_HASHING_CFG[14].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[15][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[15][1:0], ENTROPY_FWD_HASHING_CFG[15].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[16][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[16][1:0], ENTROPY_FWD_HASHING_CFG[16].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[17][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[17][1:0], ENTROPY_FWD_HASHING_CFG[17].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[18][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[18][1:0], ENTROPY_FWD_HASHING_CFG[18].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[19][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[19][1:0], ENTROPY_FWD_HASHING_CFG[19].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[20][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[20][1:0], ENTROPY_FWD_HASHING_CFG[20].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[21][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[21][1:0], ENTROPY_FWD_HASHING_CFG[21].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[22][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[22][1:0], ENTROPY_FWD_HASHING_CFG[22].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[23][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[23][1:0], ENTROPY_FWD_HASHING_CFG[23].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[24][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[24][1:0], ENTROPY_FWD_HASHING_CFG[24].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[25][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[25][1:0], ENTROPY_FWD_HASHING_CFG[25].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[26][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[26][1:0], ENTROPY_FWD_HASHING_CFG[26].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[27][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[27][1:0], ENTROPY_FWD_HASHING_CFG[27].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[28][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[28][1:0], ENTROPY_FWD_HASHING_CFG[28].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[29][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[29][1:0], ENTROPY_FWD_HASHING_CFG[29].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[30][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[30][1:0], ENTROPY_FWD_HASHING_CFG[30].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[31][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[31][1:0], ENTROPY_FWD_HASHING_CFG[31].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[32][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[32][1:0], ENTROPY_FWD_HASHING_CFG[32].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[33][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[33][1:0], ENTROPY_FWD_HASHING_CFG[33].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[34][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[34][1:0], ENTROPY_FWD_HASHING_CFG[34].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[35][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[35][1:0], ENTROPY_FWD_HASHING_CFG[35].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[36][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[36][1:0], ENTROPY_FWD_HASHING_CFG[36].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[37][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[37][1:0], ENTROPY_FWD_HASHING_CFG[37].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[38][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[38][1:0], ENTROPY_FWD_HASHING_CFG[38].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[39][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[39][1:0], ENTROPY_FWD_HASHING_CFG[39].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[40][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[40][1:0], ENTROPY_FWD_HASHING_CFG[40].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[41][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[41][1:0], ENTROPY_FWD_HASHING_CFG[41].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[42][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[42][1:0], ENTROPY_FWD_HASHING_CFG[42].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[43][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[43][1:0], ENTROPY_FWD_HASHING_CFG[43].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[44][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[44][1:0], ENTROPY_FWD_HASHING_CFG[44].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[45][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[45][1:0], ENTROPY_FWD_HASHING_CFG[45].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[46][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[46][1:0], ENTROPY_FWD_HASHING_CFG[46].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[47][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[47][1:0], ENTROPY_FWD_HASHING_CFG[47].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[48][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[48][1:0], ENTROPY_FWD_HASHING_CFG[48].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[49][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[49][1:0], ENTROPY_FWD_HASHING_CFG[49].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[50][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[50][1:0], ENTROPY_FWD_HASHING_CFG[50].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[51][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[51][1:0], ENTROPY_FWD_HASHING_CFG[51].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[52][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[52][1:0], ENTROPY_FWD_HASHING_CFG[52].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[53][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[53][1:0], ENTROPY_FWD_HASHING_CFG[53].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[54][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[54][1:0], ENTROPY_FWD_HASHING_CFG[54].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[55][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[55][1:0], ENTROPY_FWD_HASHING_CFG[55].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[56][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[56][1:0], ENTROPY_FWD_HASHING_CFG[56].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[57][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[57][1:0], ENTROPY_FWD_HASHING_CFG[57].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[58][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[58][1:0], ENTROPY_FWD_HASHING_CFG[58].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[59][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[59][1:0], ENTROPY_FWD_HASHING_CFG[59].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[60][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[60][1:0], ENTROPY_FWD_HASHING_CFG[60].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[61][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[61][1:0], ENTROPY_FWD_HASHING_CFG[61].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[62][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[62][1:0], ENTROPY_FWD_HASHING_CFG[62].ROTATION_B[1:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 2'h1, up_ENTROPY_FWD_HASHING_CFG_ROTATION_B[63][0], nxt_ENTROPY_FWD_HASHING_CFG_ROTATION_B[63][1:0], ENTROPY_FWD_HASHING_CFG[63].ROTATION_B[1:0])

// ----------------------------------------------------------------------
// ENTROPY_FWD_HASHING_CFG.ECMP_ROTATION x1 RW, using RW template.
logic [63:0][0:0] up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION;
always_comb begin
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[0] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[0] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[1] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[1] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[2] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[2] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[3] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[3] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[4] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[4] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[5] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[5] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[6] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[6] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[7] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[7] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[8] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[8] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[9] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[9] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[10] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[10] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[11] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[11] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[12] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[12] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[13] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[13] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[14] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[14] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[15] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[15] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[16] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[16] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[17] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[17] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[18] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[18] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[19] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[19] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[20] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[20] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[21] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[21] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[22] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[22] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[23] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[23] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[24] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[24] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[25] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[25] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[26] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[26] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[27] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[27] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[28] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[28] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[29] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[29] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[30] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[30] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[31] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[31] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[32] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[32] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[33] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[33] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[34] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[34] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[35] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[35] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[36] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[36] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[37] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[37] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[38] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[38] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[39] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[39] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[40] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[40] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[41] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[41] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[42] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[42] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[43] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[43] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[44] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[44] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[45] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[45] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[46] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[46] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[47] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[47] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[48] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[48] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[49] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[49] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[50] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[50] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[51] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[51] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[52] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[52] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[53] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[53] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[54] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[54] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[55] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[55] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[56] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[56] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[57] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[57] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[58] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[58] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[59] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[59] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[60] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[60] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[61] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[61] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[62] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[62] }} &
    be[1:1]);
 up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[63] =
    ({1{write_req_ENTROPY_FWD_HASHING_CFG[63] }} &
    be[1:1]);
end

logic [63:0][0:0] nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION;
always_comb begin
 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[0] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[1] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[2] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[3] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[4] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[5] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[6] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[7] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[8] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[9] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[10] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[11] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[12] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[13] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[14] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[15] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[16] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[17] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[18] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[19] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[20] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[21] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[22] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[23] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[24] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[25] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[26] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[27] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[28] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[29] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[30] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[31] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[32] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[33] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[34] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[35] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[36] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[37] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[38] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[39] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[40] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[41] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[42] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[43] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[44] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[45] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[46] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[47] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[48] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[49] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[50] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[51] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[52] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[53] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[54] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[55] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[56] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[57] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[58] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[59] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[60] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[61] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[62] = write_data[12:12];

 nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[63] = write_data[12:12];

end


`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[0][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[0][0:0], ENTROPY_FWD_HASHING_CFG[0].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[1][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[1][0:0], ENTROPY_FWD_HASHING_CFG[1].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[2][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[2][0:0], ENTROPY_FWD_HASHING_CFG[2].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[3][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[3][0:0], ENTROPY_FWD_HASHING_CFG[3].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[4][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[4][0:0], ENTROPY_FWD_HASHING_CFG[4].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[5][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[5][0:0], ENTROPY_FWD_HASHING_CFG[5].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[6][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[6][0:0], ENTROPY_FWD_HASHING_CFG[6].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[7][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[7][0:0], ENTROPY_FWD_HASHING_CFG[7].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[8][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[8][0:0], ENTROPY_FWD_HASHING_CFG[8].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[9][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[9][0:0], ENTROPY_FWD_HASHING_CFG[9].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[10][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[10][0:0], ENTROPY_FWD_HASHING_CFG[10].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[11][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[11][0:0], ENTROPY_FWD_HASHING_CFG[11].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[12][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[12][0:0], ENTROPY_FWD_HASHING_CFG[12].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[13][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[13][0:0], ENTROPY_FWD_HASHING_CFG[13].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[14][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[14][0:0], ENTROPY_FWD_HASHING_CFG[14].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[15][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[15][0:0], ENTROPY_FWD_HASHING_CFG[15].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[16][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[16][0:0], ENTROPY_FWD_HASHING_CFG[16].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[17][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[17][0:0], ENTROPY_FWD_HASHING_CFG[17].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[18][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[18][0:0], ENTROPY_FWD_HASHING_CFG[18].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[19][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[19][0:0], ENTROPY_FWD_HASHING_CFG[19].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[20][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[20][0:0], ENTROPY_FWD_HASHING_CFG[20].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[21][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[21][0:0], ENTROPY_FWD_HASHING_CFG[21].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[22][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[22][0:0], ENTROPY_FWD_HASHING_CFG[22].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[23][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[23][0:0], ENTROPY_FWD_HASHING_CFG[23].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[24][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[24][0:0], ENTROPY_FWD_HASHING_CFG[24].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[25][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[25][0:0], ENTROPY_FWD_HASHING_CFG[25].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[26][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[26][0:0], ENTROPY_FWD_HASHING_CFG[26].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[27][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[27][0:0], ENTROPY_FWD_HASHING_CFG[27].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[28][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[28][0:0], ENTROPY_FWD_HASHING_CFG[28].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[29][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[29][0:0], ENTROPY_FWD_HASHING_CFG[29].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[30][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[30][0:0], ENTROPY_FWD_HASHING_CFG[30].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[31][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[31][0:0], ENTROPY_FWD_HASHING_CFG[31].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[32][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[32][0:0], ENTROPY_FWD_HASHING_CFG[32].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[33][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[33][0:0], ENTROPY_FWD_HASHING_CFG[33].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[34][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[34][0:0], ENTROPY_FWD_HASHING_CFG[34].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[35][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[35][0:0], ENTROPY_FWD_HASHING_CFG[35].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[36][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[36][0:0], ENTROPY_FWD_HASHING_CFG[36].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[37][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[37][0:0], ENTROPY_FWD_HASHING_CFG[37].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[38][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[38][0:0], ENTROPY_FWD_HASHING_CFG[38].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[39][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[39][0:0], ENTROPY_FWD_HASHING_CFG[39].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[40][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[40][0:0], ENTROPY_FWD_HASHING_CFG[40].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[41][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[41][0:0], ENTROPY_FWD_HASHING_CFG[41].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[42][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[42][0:0], ENTROPY_FWD_HASHING_CFG[42].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[43][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[43][0:0], ENTROPY_FWD_HASHING_CFG[43].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[44][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[44][0:0], ENTROPY_FWD_HASHING_CFG[44].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[45][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[45][0:0], ENTROPY_FWD_HASHING_CFG[45].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[46][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[46][0:0], ENTROPY_FWD_HASHING_CFG[46].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[47][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[47][0:0], ENTROPY_FWD_HASHING_CFG[47].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[48][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[48][0:0], ENTROPY_FWD_HASHING_CFG[48].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[49][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[49][0:0], ENTROPY_FWD_HASHING_CFG[49].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[50][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[50][0:0], ENTROPY_FWD_HASHING_CFG[50].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[51][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[51][0:0], ENTROPY_FWD_HASHING_CFG[51].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[52][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[52][0:0], ENTROPY_FWD_HASHING_CFG[52].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[53][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[53][0:0], ENTROPY_FWD_HASHING_CFG[53].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[54][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[54][0:0], ENTROPY_FWD_HASHING_CFG[54].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[55][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[55][0:0], ENTROPY_FWD_HASHING_CFG[55].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[56][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[56][0:0], ENTROPY_FWD_HASHING_CFG[56].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[57][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[57][0:0], ENTROPY_FWD_HASHING_CFG[57].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[58][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[58][0:0], ENTROPY_FWD_HASHING_CFG[58].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[59][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[59][0:0], ENTROPY_FWD_HASHING_CFG[59].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[60][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[60][0:0], ENTROPY_FWD_HASHING_CFG[60].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[61][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[61][0:0], ENTROPY_FWD_HASHING_CFG[61].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[62][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[62][0:0], ENTROPY_FWD_HASHING_CFG[62].ECMP_ROTATION[0:0])
`RTLGEN_MBY_PPE_ENTROPY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[63][0], nxt_ENTROPY_FWD_HASHING_CFG_ECMP_ROTATION[63][0:0], ENTROPY_FWD_HASHING_CFG[63].ECMP_ROTATION[0:0])


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_ENTROPY_MAP_MEM) 
           {40'b0??,4'h?,1'b?},
           {40'b10?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_ENTROPY_HASH_CFG0;
                    ack.read_miss = handcode_error_ENTROPY_HASH_CFG0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'b10??,4'h?,1'b?},
           {40'b110?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_ENTROPY_HASH_CFG1;
                    ack.read_miss = handcode_error_ENTROPY_HASH_CFG1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'b111?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_ENTROPY_META_CFG;
                    ack.read_miss = handcode_error_ENTROPY_META_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h10,4'b00??,1'b?},
           {40'h10,4'b010?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_ENTROPY_HASH_SYM8;
                    ack.read_miss = handcode_error_ENTROPY_HASH_SYM8;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h10,4'b10??,1'b?},
           {40'h10,4'b110?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_ENTROPY_HASH_SYM16;
                    ack.read_miss = handcode_error_ENTROPY_HASH_SYM16;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h11,4'b00??,1'b?},
           {40'h11,4'b010?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_ENTROPY_HASH_SYM32;
                    ack.read_miss = handcode_error_ENTROPY_HASH_SYM32;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h2,4'b0???,4'h?,1'b?},
           {36'h2,4'b10??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_ENTROPY_HASH_KEY_MASK;
                    ack.read_miss = handcode_error_ENTROPY_HASH_KEY_MASK;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[17]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[18]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[19]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[20]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[21]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[22]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[23]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[24]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[25]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[26]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[27]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[28]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[29]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[30]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[31]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[32]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[33]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[34]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[35]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[36]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[37]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[38]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[39]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[40]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[41]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[42]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[43]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[44]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[45]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[46]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[47]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[48]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[49]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[50]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[51]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[52]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[53]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[54]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[55]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[56]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[57]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[58]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[59]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[60]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[61]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[62]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[63]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_ENTROPY_MAP_MEM) 
           {40'b0??,4'h?,1'b?},
           {40'b10?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_ENTROPY_HASH_CFG0;
                    ack.write_miss = handcode_error_ENTROPY_HASH_CFG0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'b10??,4'h?,1'b?},
           {40'b110?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_ENTROPY_HASH_CFG1;
                    ack.write_miss = handcode_error_ENTROPY_HASH_CFG1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'b111?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_ENTROPY_META_CFG;
                    ack.write_miss = handcode_error_ENTROPY_META_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h10,4'b00??,1'b?},
           {40'h10,4'b010?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_ENTROPY_HASH_SYM8;
                    ack.write_miss = handcode_error_ENTROPY_HASH_SYM8;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h10,4'b10??,1'b?},
           {40'h10,4'b110?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_ENTROPY_HASH_SYM16;
                    ack.write_miss = handcode_error_ENTROPY_HASH_SYM16;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h11,4'b00??,1'b?},
           {40'h11,4'b010?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_ENTROPY_HASH_SYM32;
                    ack.write_miss = handcode_error_ENTROPY_HASH_SYM32;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h2,4'b0???,4'h?,1'b?},
           {36'h2,4'b10??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_ENTROPY_HASH_KEY_MASK;
                    ack.write_miss = handcode_error_ENTROPY_HASH_KEY_MASK;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[17]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[18]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[19]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[20]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[21]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[22]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[23]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[24]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[25]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[26]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[27]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[28]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[29]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[30]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[31]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[32]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[33]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[34]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[35]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[36]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[37]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[38]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[39]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[40]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[41]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[42]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[43]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[44]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[45]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[46]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[47]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[48]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[49]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[50]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[51]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[52]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[53]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[54]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[55]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[56]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[57]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[58]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[59]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[60]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[61]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[62]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[63]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_ENTROPY_MAP_MEM) 
           {40'b0??,4'h?,1'b?},
           {40'b10?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = handcode_reg_rdata_ENTROPY_HASH_CFG0;
                 default: read_data = '0;
              endcase
           end
           {40'b10??,4'h?,1'b?},
           {40'b110?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = handcode_reg_rdata_ENTROPY_HASH_CFG1;
                 default: read_data = '0;
              endcase
           end
           {40'b111?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = handcode_reg_rdata_ENTROPY_META_CFG;
                 default: read_data = '0;
              endcase
           end
           {40'h10,4'b00??,1'b?},
           {40'h10,4'b010?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = handcode_reg_rdata_ENTROPY_HASH_SYM8;
                 default: read_data = '0;
              endcase
           end
           {40'h10,4'b10??,1'b?},
           {40'h10,4'b110?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = handcode_reg_rdata_ENTROPY_HASH_SYM16;
                 default: read_data = '0;
              endcase
           end
           {40'h11,4'b00??,1'b?},
           {40'h11,4'b010?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = handcode_reg_rdata_ENTROPY_HASH_SYM32;
                 default: read_data = '0;
              endcase
           end
           {36'h2,4'b0???,4'h?,1'b?},
           {36'h2,4'b10??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = handcode_reg_rdata_ENTROPY_HASH_KEY_MASK;
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[0]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[1]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[2]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[3]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[4]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[5]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[6]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[7]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[8]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[9]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[10]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[11]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[12]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[13]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[14]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[15]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[16]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[17]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[17]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[18]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[18]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[19]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[19]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[20]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[20]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[21]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[21]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[22]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[22]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[23]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[23]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[24]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[24]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[25]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[25]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[26]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[26]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[27]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[27]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[28]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[28]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[29]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[29]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[30]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[30]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[31]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[31]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[32]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[32]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[33]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[33]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[34]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[34]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[35]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[35]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[36]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[36]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[37]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[37]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[38]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[38]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[39]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[39]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[40]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[40]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[41]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[41]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[42]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[42]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[43]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[43]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[44]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[44]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[45]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[45]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[46]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[46]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[47]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[47]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[48]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[48]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[49]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[49]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[50]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[50]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[51]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[51]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[52]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[52]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[53]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[53]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[54]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[54]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[55]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[55]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[56]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[56]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[57]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[57]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[58]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[58]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[59]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[59]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[60]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[60]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[61]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[61]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[62]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[62]};
                 default: read_data = '0;
              endcase
           end
           ENTROPY_FWD_HASHING_CFG_DECODE_ADDR[63]: begin
              unique casez ({req_fid,req_bar})
                 {ENTROPY_SB_FID,ENTROPY_SB_BAR}: read_data = {ENTROPY_FWD_HASHING_CFG[63]};
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {


// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
