magic
tech scmos
timestamp 962519208
<< ndiffusion >>
rect 0 37 6 38
rect 0 34 6 35
rect 0 30 2 34
rect 0 29 6 30
rect 0 26 6 27
rect 0 13 6 14
rect 0 7 6 11
rect 0 4 6 5
rect 0 -1 6 0
rect 0 -4 6 -3
rect 0 -8 2 -4
rect 0 -9 6 -8
rect 0 -12 6 -11
<< pdiffusion >>
rect 18 35 24 36
rect 18 29 24 33
rect 18 23 24 27
rect 18 15 24 19
rect 18 12 24 13
rect 22 8 24 12
rect 18 7 24 8
rect 18 4 24 5
rect 18 -1 24 0
rect 18 -7 24 -3
rect 18 -10 24 -9
<< ntransistor >>
rect 0 35 6 37
rect 0 27 6 29
rect 0 11 6 13
rect 0 5 6 7
rect 0 -3 6 -1
rect 0 -11 6 -9
<< ptransistor >>
rect 18 33 24 35
rect 18 27 24 29
rect 18 13 24 15
rect 18 5 24 7
rect 18 -3 24 -1
rect 18 -9 24 -7
<< polysilicon >>
rect -3 35 0 37
rect 6 35 10 37
rect 8 33 18 35
rect 24 33 27 35
rect -3 27 0 29
rect 6 27 18 29
rect 24 27 27 29
rect 12 15 14 17
rect 12 13 18 15
rect 24 13 27 15
rect -3 11 0 13
rect 6 11 14 13
rect -3 5 0 7
rect 6 5 10 7
rect 14 5 18 7
rect 24 5 27 7
rect -3 -3 0 -1
rect 6 -3 18 -1
rect 24 -3 27 -1
rect 8 -9 18 -7
rect 24 -9 27 -7
rect -3 -11 0 -9
rect 6 -11 10 -9
<< ndcontact >>
rect 0 38 6 42
rect 2 30 6 34
rect 0 22 6 26
rect 0 14 6 18
rect 0 0 6 4
rect 2 -8 6 -4
rect 0 -16 6 -12
<< pdcontact >>
rect 18 36 24 40
rect 18 19 24 23
rect 18 8 22 12
rect 18 0 24 4
rect 18 -14 24 -10
<< polycontact >>
rect 10 17 14 21
rect 10 3 14 7
<< metal1 >>
rect 0 38 6 42
rect 18 36 24 40
rect 2 33 6 34
rect 18 33 21 36
rect 2 30 21 33
rect 0 22 6 26
rect 10 21 13 30
rect 0 14 6 18
rect 10 17 14 21
rect 18 19 24 23
rect 3 13 6 14
rect 3 12 21 13
rect 3 10 22 12
rect 18 8 22 10
rect 0 0 6 4
rect 10 3 14 7
rect 10 -4 13 3
rect 18 0 24 4
rect 2 -7 21 -4
rect 2 -8 6 -7
rect 18 -10 21 -7
rect 0 -16 6 -12
rect 18 -14 24 -10
<< labels >>
rlabel polysilicon 25 6 25 6 1 _a_01
rlabel polysilicon 25 14 25 14 1 _a_23
rlabel polysilicon -1 28 -1 28 1 a2
rlabel polysilicon -1 36 -1 36 1 a3
rlabel polysilicon -1 -2 -1 -2 1 a1
rlabel polysilicon -1 -10 -1 -10 1 a0
rlabel polysilicon 25 28 25 28 1 a2
rlabel polysilicon 25 34 25 34 1 a3
rlabel polysilicon 25 -2 25 -2 1 a1
rlabel polysilicon 25 -8 25 -8 1 a0
rlabel polysilicon -1 6 -1 6 1 _a_01
rlabel polysilicon -1 12 -1 12 1 _a_23
rlabel space -3 25 3 43 7 ^n1
rlabel space -3 3 1 19 7 ^n2
rlabel space 22 3 27 20 3 ^p2
rlabel space 23 22 27 41 3 ^p1
rlabel space 23 -15 27 1 3 ^p3
rlabel space -3 -17 3 1 7 ^n3
rlabel pdcontact 20 10 20 10 1 av
rlabel ndcontact 4 16 4 16 1 av
rlabel ndcontact 4 -6 4 -6 5 _a_01
rlabel pdcontact 20 -12 20 -12 5 _a_01
rlabel pdcontact 20 38 20 38 1 _a_23
rlabel ndcontact 4 32 4 32 1 _a_23
rlabel ndcontact 4 -14 4 -14 5 GND!
rlabel ndcontact 4 2 4 2 5 GND!
rlabel ndcontact 4 24 4 24 1 GND!
rlabel ndcontact 4 40 4 40 1 GND!
rlabel pdcontact 20 2 20 2 1 Vdd!
rlabel metal1 21 21 21 21 1 Vdd!
<< end >>
