// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

module read_ecc
  (
input  logic [1013-1:0] i_data,
input  logic [11-1:0] i_chk,

output logic          o_err_detect,
output logic          o_err_multpl,
output logic [1013-1:0] o_data
  );
logic  xor0000;
logic  xor0001;
logic  xor0002;
logic  xor0003;
logic  xor0004;
logic  xor0005;
logic  xor0006;
logic  xor0007;
logic  xor0008;
logic  xor0009;
logic  xor0010;
logic  xor0011;
logic  xor0012;
logic  xor0013;
logic  xor0014;
logic  xor0015;
logic  xor0016;
logic  xor0017;
logic  xor0018;
logic  xor0019;
logic  xor0020;
logic  xor0021;
logic  xor0022;
logic  xor0023;
logic  xor0024;
logic  xor0025;
logic  xor0026;
logic  xor0027;
logic  xor0028;
logic  xor0029;
logic  xor0030;
logic  xor0031;
logic  xor0032;
logic  xor0033;
logic  xor0034;
logic  xor0035;
logic  xor0036;
logic  xor0037;
logic  xor0038;
logic  xor0039;
logic  xor0040;
logic  xor0041;
logic  xor0042;
logic  xor0043;
logic  xor0044;
logic  xor0045;
logic  xor0046;
logic  xor0047;
logic  xor0048;
logic  xor0049;
logic  xor0050;
logic  xor0051;
logic  xor0052;
logic  xor0053;
logic  xor0054;
logic  xor0055;
logic  xor0056;
logic  xor0057;
logic  xor0058;
logic  xor0059;
logic  xor0060;
logic  xor0061;
logic  xor0062;
logic  xor0063;
logic  xor0064;
logic  xor0065;
logic  xor0066;
logic  xor0067;
logic  xor0068;
logic  xor0069;
logic  xor0070;
logic  xor0071;
logic  xor0072;
logic  xor0073;
logic  xor0074;
logic  xor0075;
logic  xor0076;
logic  xor0077;
logic  xor0078;
logic  xor0079;
logic  xor0080;
logic  xor0081;
logic  xor0082;
logic  xor0083;
logic  xor0084;
logic  xor0085;
logic  xor0086;
logic  xor0087;
logic  xor0088;
logic  xor0089;
logic  xor0090;
logic  xor0091;
logic  xor0092;
logic  xor0093;
logic  xor0094;
logic  xor0095;
logic  xor0096;
logic  xor0097;
logic  xor0098;
logic  xor0099;
logic  xor0100;
logic  xor0101;
logic  xor0102;
logic  xor0103;
logic  xor0104;
logic  xor0105;
logic  xor0106;
logic  xor0107;
logic  xor0108;
logic  xor0109;
logic  xor0110;
logic  xor0111;
logic  xor0112;
logic  xor0113;
logic  xor0114;
logic  xor0115;
logic  xor0116;
logic  xor0117;
logic  xor0118;
logic  xor0119;
logic  xor0120;
logic  xor0121;
logic  xor0122;
logic  xor0123;
logic  xor0124;
logic  xor0125;
logic  xor0126;
logic  xor0127;
logic  xor0128;
logic  xor0129;
logic  xor0130;
logic  xor0131;
logic  xor0132;
logic  xor0133;
logic  xor0134;
logic  xor0135;
logic  xor0136;
logic  xor0137;
logic  xor0138;
logic  xor0139;
logic  xor0140;
logic  xor0141;
logic  xor0142;
logic  xor0143;
logic  xor0144;
logic  xor0145;
logic  xor0146;
logic  xor0147;
logic  xor0148;
logic  xor0149;
logic  xor0150;
logic  xor0151;
logic  xor0152;
logic  xor0153;
logic  xor0154;
logic  xor0155;
logic  xor0156;
logic  xor0157;
logic  xor0158;
logic  xor0159;
logic  xor0160;
logic  xor0161;
logic  xor0162;
logic  xor0163;
logic  xor0164;
logic  xor0165;
logic  xor0166;
logic  xor0167;
logic  xor0168;
logic  xor0169;
logic  xor0170;
logic  xor0171;
logic  xor0172;
logic  xor0173;
logic  xor0174;
logic  xor0175;
logic  xor0176;
logic  xor0177;
logic  xor0178;
logic  xor0179;
logic  xor0180;
logic  xor0181;
logic  xor0182;
logic  xor0183;
logic  xor0184;
logic  xor0185;
logic  xor0186;
logic  xor0187;
logic  xor0188;
logic  xor0189;
logic  xor0190;
logic  xor0191;
logic  xor0192;
logic  xor0193;
logic  xor0194;
logic  xor0195;
logic  xor0196;
logic  xor0197;
logic  xor0198;
logic  xor0199;
logic  xor0200;
logic  xor0201;
logic  xor0202;
logic  xor0203;
logic  xor0204;
logic  xor0205;
logic  xor0206;
logic  xor0207;
logic  xor0208;
logic  xor0209;
logic  xor0210;
logic  xor0211;
logic  xor0212;
logic  xor0213;
logic  xor0214;
logic  xor0215;
logic  xor0216;
logic  xor0217;
logic  xor0218;
logic  xor0219;
logic  xor0220;
logic  xor0221;
logic  xor0222;
logic  xor0223;
logic  xor0224;
logic  xor0225;
logic  xor0226;
logic  xor0227;
logic  xor0228;
logic  xor0229;
logic  xor0230;
logic  xor0231;
logic  xor0232;
logic  xor0233;
logic  xor0234;
logic  xor0235;
logic  xor0236;
logic  xor0237;
logic  xor0238;
logic  xor0239;
logic  xor0240;
logic  xor0241;
logic  xor0242;
logic  xor0243;
logic  xor0244;
logic  xor0245;
logic  xor0246;
logic  xor0247;
logic  xor0248;
logic  xor0249;
logic  xor0250;
logic  xor0251;
logic  xor0252;
logic  xor0253;
logic  xor0254;
logic  xor0255;
logic  xor0256;
logic  xor0257;
logic  xor0258;
logic  xor0259;
logic  xor0260;
logic  xor0261;
logic  xor0262;
logic  xor0263;
logic  xor0264;
logic  xor0265;
logic  xor0266;
logic  xor0267;
logic  xor0268;
logic  xor0269;
logic  xor0270;
logic  xor0271;
logic  xor0272;
logic  xor0273;
logic  xor0274;
logic  xor0275;
logic  xor0276;
logic  xor0277;
logic  xor0278;
logic  xor0279;
logic  xor0280;
logic  xor0281;
logic  xor0282;
logic  xor0283;
logic  xor0284;
logic  xor0285;
logic  xor0286;
logic  xor0287;
logic  xor0288;
logic  xor0289;
logic  xor0290;
logic  xor0291;
logic  xor0292;
logic  xor0293;
logic  xor0294;
logic  xor0295;
logic  xor0296;
logic  xor0297;
logic  xor0298;
logic  xor0299;
logic  xor0300;
logic  xor0301;
logic  xor0302;
logic  xor0303;
logic  xor0304;
logic  xor0305;
logic  xor0306;
logic  xor0307;
logic  xor0308;
logic  xor0309;
logic  xor0310;
logic  xor0311;
logic  xor0312;
logic  xor0313;
logic  xor0314;
logic  xor0315;
logic  xor0316;
logic  xor0317;
logic  xor0318;
logic  xor0319;
logic  xor0320;
logic  xor0321;
logic  xor0322;
logic  xor0323;
logic  xor0324;
logic  xor0325;
logic  xor0326;
logic  xor0327;
logic  xor0328;
logic  xor0329;
logic  xor0330;
logic  xor0331;
logic  xor0332;
logic  xor0333;
logic  xor0334;
logic  xor0335;
logic  xor0336;
logic  xor0337;
logic  xor0338;
logic  xor0339;
logic  xor0340;
logic  xor0341;
logic  xor0342;
logic  xor0343;
logic  xor0344;
logic  xor0345;
logic  xor0346;
logic  xor0347;
logic  xor0348;
logic  xor0349;
logic  xor0350;
logic  xor0351;
logic  xor0352;
logic  xor0353;
logic  xor0354;
logic  xor0355;
logic  xor0356;
logic  xor0357;
logic  xor0358;
logic  xor0359;
logic  xor0360;
logic  xor0361;
logic  xor0362;
logic  xor0363;
logic  xor0364;
logic  xor0365;
logic  xor0366;
logic  xor0367;
logic  xor0368;
logic  xor0369;
logic  xor0370;
logic  xor0371;
logic  xor0372;
logic  xor0373;
logic  xor0374;
logic  xor0375;
logic  xor0376;
logic  xor0377;
logic  xor0378;
logic  xor0379;
logic  xor0380;
logic  xor0381;
logic  xor0382;
logic  xor0383;
logic  xor0384;
logic  xor0385;
logic  xor0386;
logic  xor0387;
logic  xor0388;
logic  xor0389;
logic  xor0390;
logic  xor0391;
logic  xor0392;
logic  xor0393;
logic  xor0394;
logic  xor0395;
logic  xor0396;
logic  xor0397;
logic  xor0398;
logic  xor0399;
logic  xor0400;
logic  xor0401;
logic  xor0402;
logic  xor0403;
logic  xor0404;
logic  xor0405;
logic  xor0406;
logic  xor0407;
logic  xor0408;
logic  xor0409;
logic  xor0410;
logic  xor0411;
logic  xor0412;
logic  xor0413;
logic  xor0414;
logic  xor0415;
logic  xor0416;
logic  xor0417;
logic  xor0418;
logic  xor0419;
logic  xor0420;
logic  xor0421;
logic  xor0422;
logic  xor0423;
logic  xor0424;
logic  xor0425;
logic  xor0426;
logic  xor0427;
logic  xor0428;
logic  xor0429;
logic  xor0430;
logic  xor0431;
logic  xor0432;
logic  xor0433;
logic  xor0434;
logic  xor0435;
logic  xor0436;
logic  xor0437;
logic  xor0438;
logic  xor0439;
logic  xor0440;
logic  xor0441;
logic  xor0442;
logic  xor0443;
logic  xor0444;
logic  xor0445;
logic  xor0446;
logic  xor0447;
logic  xor0448;
logic  xor0449;
logic  xor0450;
logic  xor0451;
logic  xor0452;
logic  xor0453;
logic  xor0454;
logic  xor0455;
logic  xor0456;
logic  xor0457;
logic  xor0458;
logic  xor0459;
logic  xor0460;
logic  xor0461;
logic  xor0462;
logic  xor0463;
logic  xor0464;
logic  xor0465;
logic  xor0466;
logic  xor0467;
logic  xor0468;
logic  xor0469;
logic  xor0470;
logic  xor0471;
logic  xor0472;
logic  xor0473;
logic  xor0474;
logic  xor0475;
logic  xor0476;
logic  xor0477;
logic  xor0478;
logic  xor0479;
logic  xor0480;
logic  xor0481;
logic  xor0482;
logic  xor0483;
logic  xor0484;
logic  xor0485;
logic  xor0486;
logic  xor0487;
logic  xor0488;
logic  xor0489;
logic  xor0490;
logic  xor0491;
logic  xor0492;
logic  xor0493;
logic  xor0494;
logic  xor0495;
logic  xor0496;
logic  xor0497;
logic  xor0498;
logic  xor0499;
logic  xor0500;
logic  xor0501;
logic  xor0502;
logic  xor0503;
logic  xor0504;
logic  xor0505;
logic  xor0506;
logic  xor0507;
logic  xor0508;
logic  xor0509;
logic  xor0510;
logic  xor0511;
logic  xor0512;
logic  xor0513;
logic  xor0514;
logic  xor0515;
logic  xor0516;
logic  xor0517;
logic  xor0518;
logic  xor0519;
logic  xor0520;
logic  xor0521;
logic  xor0522;
logic  xor0523;
logic  xor0524;
logic  xor0525;
logic  xor0526;
logic  xor0527;
logic  xor0528;
logic  xor0529;
logic  xor0530;
logic  xor0531;
logic  xor0532;
logic  xor0533;
logic  xor0534;
logic  xor0535;
logic  xor0536;
logic  xor0537;
logic  xor0538;
logic  xor0539;
logic  xor0540;
logic  xor0541;
logic  xor0542;
logic  xor0543;
logic  xor0544;
logic  xor0545;
logic  xor0546;
logic  xor0547;
logic  xor0548;
logic  xor0549;
logic  xor0550;
logic  xor0551;
logic  xor0552;
logic  xor0553;
logic  xor0554;
logic  xor0555;
logic  xor0556;
logic  xor0557;
logic  xor0558;
logic  xor0559;
logic  xor0560;
logic  xor0561;
logic  xor0562;
logic  xor0563;
logic  xor0564;
logic  xor0565;
logic  xor0566;
logic  xor0567;
logic  xor0568;
logic  xor0569;
logic  xor0570;
logic  xor0571;
logic  xor0572;
logic  xor0573;
logic  xor0574;
logic  xor0575;
logic  xor0576;
logic  xor0577;
logic  xor0578;
logic  xor0579;
logic  xor0580;
logic  xor0581;
logic  xor0582;
logic  xor0583;
logic  xor0584;
logic  xor0585;
logic  xor0586;
logic  xor0587;
logic  xor0588;
logic  xor0589;
logic  xor0590;
logic  xor0591;
logic  xor0592;
logic  xor0593;
logic  xor0594;
logic  xor0595;
logic  xor0596;
logic  xor0597;
logic  xor0598;
logic  xor0599;
logic  xor0600;
logic  xor0601;
logic  xor0602;
logic  xor0603;
logic  xor0604;
logic  xor0605;
logic  xor0606;
logic  xor0607;
logic  xor0608;
logic  xor0609;
logic  xor0610;
logic  xor0611;
logic  xor0612;
logic  xor0613;
logic  xor0614;
logic  xor0615;
logic  xor0616;
logic  xor0617;
logic  xor0618;
logic  xor0619;
logic  xor0620;
logic  xor0621;
logic  xor0622;
logic  xor0623;
logic  xor0624;
logic  xor0625;
logic  xor0626;
logic  xor0627;
logic  xor0628;
logic  xor0629;
logic  xor0630;
logic  xor0631;
logic  xor0632;
logic  xor0633;
logic  xor0634;
logic  xor0635;
logic  xor0636;
logic  xor0637;
logic  xor0638;
logic  xor0639;
logic  xor0640;
logic  xor0641;
logic  xor0642;
logic  xor0643;
logic  xor0644;
logic  xor0645;
logic  xor0646;
logic  xor0647;
logic  xor0648;
logic  xor0649;
logic  xor0650;
logic  xor0651;
logic  xor0652;
logic  xor0653;
logic  xor0654;
logic  xor0655;
logic  xor0656;
logic  xor0657;
logic  xor0658;
logic  xor0659;
logic  xor0660;
logic  xor0661;
logic  xor0662;
logic  xor0663;
logic  xor0664;
logic  xor0665;
logic  xor0666;
logic  xor0667;
logic  xor0668;
logic  xor0669;
logic  xor0670;
logic  xor0671;
logic  xor0672;
logic  xor0673;
logic  xor0674;
logic  xor0675;
logic  xor0676;
logic  xor0677;
logic  xor0678;
logic  xor0679;
logic  xor0680;
logic  xor0681;
logic  xor0682;
logic  xor0683;
logic  xor0684;
logic  xor0685;
logic  xor0686;
logic  xor0687;
logic  xor0688;
logic  xor0689;
logic  xor0690;
logic  xor0691;
logic  xor0692;
logic  xor0693;
logic  xor0694;
logic  xor0695;
logic  xor0696;
logic  xor0697;
logic  xor0698;
logic  xor0699;
logic  xor0700;
logic  xor0701;
logic  xor0702;
logic  xor0703;
logic  xor0704;
logic  xor0705;
logic  xor0706;
logic  xor0707;
logic  xor0708;
logic  xor0709;
logic  xor0710;
logic  xor0711;
logic  xor0712;
logic  xor0713;
logic  xor0714;
logic  xor0715;
logic  xor0716;
logic  xor0717;
logic  xor0718;
logic  xor0719;
logic  xor0720;
logic  xor0721;
logic  xor0722;
logic  xor0723;
logic  xor0724;
logic  xor0725;
logic  xor0726;
logic  xor0727;
logic  xor0728;
logic  xor0729;
logic  xor0730;
logic  xor0731;
logic  xor0732;
logic  xor0733;
logic  xor0734;
logic  xor0735;
logic  xor0736;
logic  xor0737;
logic  xor0738;
logic  xor0739;
logic  xor0740;
logic  xor0741;
logic  xor0742;
logic  xor0743;
logic  xor0744;
logic  xor0745;
logic  xor0746;
logic  xor0747;
logic  xor0748;
logic  xor0749;
logic  xor0750;
logic  xor0751;
logic  xor0752;
logic  xor0753;
logic  xor0754;
logic  xor0755;
logic  xor0756;
logic  xor0757;
logic  xor0758;
logic  xor0759;
logic  xor0760;
logic  xor0761;
logic  xor0762;
logic  xor0763;
logic  xor0764;
logic  xor0765;
logic  xor0766;
logic  xor0767;
logic  xor0768;
logic  xor0769;
logic  xor0770;
logic  xor0771;
logic  xor0772;
logic  xor0773;
logic  xor0774;
logic  xor0775;
logic  xor0776;
logic  xor0777;
logic  xor0778;
logic  xor0779;
logic  xor0780;
logic  xor0781;
logic  xor0782;
logic  xor0783;
logic  xor0784;
logic  xor0785;
logic  xor0786;
logic  xor0787;
logic  xor0788;
logic  xor0789;
logic  xor0790;
logic  xor0791;
logic  xor0792;
logic  xor0793;
logic  xor0794;
logic  xor0795;
logic  xor0796;
logic  xor0797;
logic  xor0798;
logic  xor0799;
logic  xor0800;
logic  xor0801;
logic  xor0802;
logic  xor0803;
logic  xor0804;
logic  xor0805;
logic  xor0806;
logic  xor0807;
logic  xor0808;
logic  xor0809;
logic  xor0810;
logic  xor0811;
logic  xor0812;
logic  xor0813;
logic  xor0814;
logic  xor0815;
logic  xor0816;
logic  xor0817;
logic  xor0818;
logic  xor0819;
logic  xor0820;
logic  xor0821;
logic  xor0822;
logic  xor0823;
logic  xor0824;
logic  xor0825;
logic  xor0826;
logic  xor0827;
logic  xor0828;
logic  xor0829;
logic  xor0830;
logic  xor0831;
logic  xor0832;
logic  xor0833;
logic  xor0834;
logic  xor0835;
logic  xor0836;
logic  xor0837;
logic  xor0838;
logic  xor0839;
logic  xor0840;
logic  xor0841;
logic  xor0842;
logic  xor0843;
logic  xor0844;
logic  xor0845;
logic  xor0846;
logic  xor0847;
logic  xor0848;
logic  xor0849;
logic  xor0850;
logic  xor0851;
logic  xor0852;
logic  xor0853;
logic  xor0854;
logic  xor0855;
logic  xor0856;
logic  xor0857;
logic  xor0858;
logic  xor0859;
logic  xor0860;
logic  xor0861;
logic  xor0862;
logic  xor0863;
logic  xor0864;
logic  xor0865;
logic  xor0866;
logic  xor0867;
logic  xor0868;
logic  xor0869;
logic  xor0870;
logic  xor0871;
logic  xor0872;
logic  xor0873;
logic  xor0874;
logic  xor0875;
logic  xor0876;
logic  xor0877;
logic  xor0878;
logic  xor0879;
logic  xor0880;
logic  xor0881;
logic  xor0882;
logic  xor0883;
logic  xor0884;
logic  xor0885;
logic  xor0886;
logic  xor0887;
logic  xor0888;
logic  xor0889;
logic  xor0890;
logic  xor0891;
logic  xor0892;
logic  xor0893;
logic  xor0894;
logic  xor0895;
logic  xor0896;
logic  xor0897;
logic  xor0898;
logic  xor0899;
logic  xor0900;
logic  xor0901;
logic  xor0902;
logic  xor0903;
logic  xor0904;
logic  xor0905;
logic  xor0906;
logic  xor0907;
logic  xor0908;
logic  xor0909;
logic  xor0910;
logic  xor0911;
logic  xor0912;
logic  xor0913;
logic  xor0914;
logic  xor0915;
logic  xor0916;
logic  xor0917;
logic  xor0918;
logic  xor0919;
logic  xor0920;
logic  xor0921;
logic  xor0922;
logic  xor0923;
logic  xor0924;
logic  xor0925;
logic  xor0926;
logic  xor0927;
logic  xor0928;
logic  xor0929;
logic  xor0930;
logic  xor0931;
logic  xor0932;
logic  xor0933;
logic  xor0934;
logic  xor0935;
logic  xor0936;
logic  xor0937;
logic  xor0938;
logic  xor0939;
logic  xor0940;
logic  xor0941;
logic  xor0942;
logic  xor0943;
logic  xor0944;
logic  xor0945;
logic  xor0946;
logic  xor0947;
logic  xor0948;
logic  xor0949;
logic  xor0950;
logic  xor0951;
logic  xor0952;
logic  xor0953;
logic  xor0954;
logic  xor0955;
logic  xor0956;
logic  xor0957;
logic  xor0958;
logic  xor0959;
logic  xor0960;
logic  xor0961;
logic[9:-1] ecc_parity;
logic[1023:0] input_data;
logic[1023:0] corrected;
logic  syn_0000_n;
logic  syn_0000;
logic  syn_0001_n;
logic  syn_0001;
logic  syn_0002_n;
logic  syn_0002;
logic  syn_0003_n;
logic  syn_0003;
logic  syn_0004_n;
logic  syn_0004;
logic  syn_0005_n;
logic  syn_0005;
logic  syn_0006_n;
logic  syn_0006;
logic  syn_0007_n;
logic  syn_0007;
logic  syn_0008_n;
logic  syn_0008;
logic  syn_0009_n;
logic  syn_0009;
logic  nand0972;
logic  nand0973;
logic  nand0974;
logic  nand0975;
logic  nand0976;
logic  nand0977;
logic  nand0978;
logic  nand0979;
logic  nand0980;
logic  nand0981;
logic  nand0982;
logic  nand0983;
logic  nand0984;
logic  nand0985;
logic  nand0986;
logic  nand0987;
logic  nand0988;
logic  nand0989;
logic  nand0990;
logic  nand0991;
logic  nand0992;
logic  nand0993;
logic  nand0994;
logic  nand0995;
logic  nand0996;
logic  nand0997;
logic  nor0998;
logic  invert0000;
logic  nor0999;
logic  invert0001;
logic  nor1000;
logic  invert0002;
logic  nor1001;
logic  invert0003;
logic  nor1002;
logic  invert0004;
logic  nor1003;
logic  invert0005;
logic  nor1004;
logic  invert0006;
logic  nor1005;
logic  invert0007;
logic  nor1006;
logic  invert0008;
logic  nor1007;
logic  invert0009;
logic  nor1008;
logic  invert0010;
logic  nor1009;
logic  invert0011;
logic  nor1010;
logic  invert0012;
logic  nor1011;
logic  invert0013;
logic  nor1012;
logic  invert0014;
logic  nor1013;
logic  invert0015;
logic  nor1014;
logic  invert0016;
logic  nor1015;
logic  invert0017;
logic  nor1016;
logic  invert0018;
logic  nor1017;
logic  invert0019;
logic  nor1018;
logic  invert0020;
logic  nor1019;
logic  invert0021;
logic  nor1020;
logic  invert0022;
logic  nor1021;
logic  invert0023;
logic  nor1022;
logic  invert0024;
logic  nor1023;
logic  invert0025;
logic  nor1024;
logic  invert0026;
logic  nor1025;
logic  invert0027;
logic  nor1026;
logic  invert0028;
logic  nor1027;
logic  invert0029;
logic  nor1028;
logic  invert0030;
logic  nor1029;
logic  invert0031;
logic  nor1030;
logic  invert0032;
logic  nor1031;
logic  invert0033;
logic  nor1032;
logic  invert0034;
logic  nor1033;
logic  invert0035;
logic  nor1034;
logic  invert0036;
logic  nor1035;
logic  invert0037;
logic  nor1036;
logic  invert0038;
logic  nor1037;
logic  invert0039;
logic  nor1038;
logic  invert0040;
logic  nor1039;
logic  invert0041;
logic  nor1040;
logic  invert0042;
logic  nor1041;
logic  invert0043;
logic  nor1042;
logic  invert0044;
logic  nor1043;
logic  invert0045;
logic  nor1044;
logic  invert0046;
logic  nor1045;
logic  invert0047;
logic  nor1046;
logic  invert0048;
logic  nor1047;
logic  invert0049;
logic  nor1048;
logic  invert0050;
logic  nor1049;
logic  invert0051;
logic  nor1050;
logic  invert0052;
logic  nor1051;
logic  invert0053;
logic  nor1052;
logic  invert0054;
logic  nor1053;
logic  invert0055;
logic  nor1054;
logic  invert0056;
logic  nor1055;
logic  invert0057;
logic  nor1056;
logic  invert0058;
logic  nor1057;
logic  invert0059;
logic  nor1058;
logic  invert0060;
logic  nor1059;
logic  invert0061;
logic  nor1060;
logic  invert0062;
logic  nor1061;
logic  invert0063;
logic  nor1062;
logic  invert0064;
logic  nor1063;
logic  invert0065;
logic  nor1064;
logic  invert0066;
logic  nor1065;
logic  invert0067;
logic  nor1066;
logic  invert0068;
logic  nor1067;
logic  invert0069;
logic  nor1068;
logic  invert0070;
logic  nor1069;
logic  invert0071;
logic  nor1070;
logic  invert0072;
logic  nor1071;
logic  invert0073;
logic  nor1072;
logic  invert0074;
logic  nor1073;
logic  invert0075;
logic  nor1074;
logic  invert0076;
logic  nor1075;
logic  invert0077;
logic  nor1076;
logic  invert0078;
logic  nor1077;
logic  invert0079;
logic  nor1078;
logic  invert0080;
logic  nor1079;
logic  invert0081;
logic  nor1080;
logic  invert0082;
logic  nor1081;
logic  invert0083;
logic  nor1082;
logic  invert0084;
logic  nor1083;
logic  invert0085;
logic  nor1084;
logic  invert0086;
logic  nor1085;
logic  invert0087;
logic  nor1086;
logic  invert0088;
logic  nor1087;
logic  invert0089;
logic  nor1088;
logic  invert0090;
logic  nor1089;
logic  invert0091;
logic  nor1090;
logic  invert0092;
logic  nor1091;
logic  invert0093;
logic  nor1092;
logic  invert0094;
logic  nor1093;
logic  invert0095;
logic  nor1094;
logic  invert0096;
logic  nor1095;
logic  invert0097;
logic  nor1096;
logic  invert0098;
logic  nor1097;
logic  invert0099;
logic  nor1098;
logic  invert0100;
logic  nor1099;
logic  invert0101;
logic  nor1100;
logic  invert0102;
logic  nor1101;
logic  invert0103;
logic  nor1102;
logic  invert0104;
logic  nor1103;
logic  invert0105;
logic  nor1104;
logic  invert0106;
logic  nor1105;
logic  invert0107;
logic  nor1106;
logic  invert0108;
logic  nor1107;
logic  invert0109;
logic  nor1108;
logic  invert0110;
logic  nor1109;
logic  invert0111;
logic  nor1110;
logic  invert0112;
logic  nor1111;
logic  invert0113;
logic  nor1112;
logic  invert0114;
logic  nor1113;
logic  invert0115;
logic  nor1114;
logic  invert0116;
logic  nor1115;
logic  invert0117;
logic  nor1116;
logic  invert0118;
logic  nor1117;
logic  invert0119;
logic  nor1118;
logic  invert0120;
logic  nor1119;
logic  invert0121;
logic  nor1120;
logic  invert0122;
logic  nor1121;
logic  invert0123;
logic  nor1122;
logic  invert0124;
logic  nor1123;
logic  invert0125;
logic  nor1124;
logic  invert0126;
logic  nor1125;
logic  invert0127;
logic  nor1126;
logic  invert0128;
logic  nor1127;
logic  invert0129;
logic  nor1128;
logic  invert0130;
logic  nor1129;
logic  invert0131;
logic  nor1130;
logic  invert0132;
logic  nor1131;
logic  invert0133;
logic  nor1132;
logic  invert0134;
logic  nor1133;
logic  invert0135;
logic  nor1134;
logic  invert0136;
logic  nor1135;
logic  invert0137;
logic  nor1136;
logic  invert0138;
logic  nor1137;
logic  invert0139;
logic  nor1138;
logic  invert0140;
logic  nor1139;
logic  invert0141;
logic  nor1140;
logic  invert0142;
logic  nor1141;
logic  invert0143;
logic  nor1142;
logic  invert0144;
logic  nor1143;
logic  invert0145;
logic  nor1144;
logic  invert0146;
logic  nor1145;
logic  invert0147;
logic  nor1146;
logic  invert0148;
logic  nor1147;
logic  invert0149;
logic  nor1148;
logic  invert0150;
logic  nor1149;
logic  invert0151;
logic  nor1150;
logic  invert0152;
logic  nor1151;
logic  invert0153;
logic  nor1152;
logic  invert0154;
logic  nor1153;
logic  invert0155;
logic  nor1154;
logic  invert0156;
logic  nor1155;
logic  invert0157;
logic  nor1156;
logic  invert0158;
logic  nor1157;
logic  invert0159;
logic  nor1158;
logic  invert0160;
logic  nor1159;
logic  invert0161;
logic  nor1160;
logic  invert0162;
logic  nor1161;
logic  invert0163;
logic  nor1162;
logic  invert0164;
logic  nor1163;
logic  invert0165;
logic  nor1164;
logic  invert0166;
logic  nor1165;
logic  invert0167;
logic  nor1166;
logic  invert0168;
logic  nor1167;
logic  invert0169;
logic  nor1168;
logic  invert0170;
logic  nor1169;
logic  invert0171;
logic  nor1170;
logic  invert0172;
logic  nor1171;
logic  invert0173;
logic  nor1172;
logic  invert0174;
logic  nor1173;
logic  invert0175;
logic  nor1174;
logic  invert0176;
logic  nor1175;
logic  invert0177;
logic  nor1176;
logic  invert0178;
logic  nor1177;
logic  invert0179;
logic  nor1178;
logic  invert0180;
logic  nor1179;
logic  invert0181;
logic  nor1180;
logic  invert0182;
logic  nor1181;
logic  invert0183;
logic  nor1182;
logic  invert0184;
logic  nor1183;
logic  invert0185;
logic  nor1184;
logic  invert0186;
logic  nor1185;
logic  invert0187;
logic  nor1186;
logic  invert0188;
logic  nor1187;
logic  invert0189;
logic  nor1188;
logic  invert0190;
logic  nor1189;
logic  invert0191;
logic  nor1190;
logic  invert0192;
logic  nor1191;
logic  invert0193;
logic  nor1192;
logic  invert0194;
logic  nor1193;
logic  invert0195;
logic  nor1194;
logic  invert0196;
logic  nor1195;
logic  invert0197;
logic  nor1196;
logic  invert0198;
logic  nor1197;
logic  invert0199;
logic  nor1198;
logic  invert0200;
logic  nor1199;
logic  invert0201;
logic  nor1200;
logic  invert0202;
logic  nor1201;
logic  invert0203;
logic  nor1202;
logic  invert0204;
logic  nor1203;
logic  invert0205;
logic  nor1204;
logic  invert0206;
logic  nor1205;
logic  invert0207;
logic  nor1206;
logic  invert0208;
logic  nor1207;
logic  invert0209;
logic  nor1208;
logic  invert0210;
logic  nor1209;
logic  invert0211;
logic  nor1210;
logic  invert0212;
logic  nor1211;
logic  invert0213;
logic  nor1212;
logic  invert0214;
logic  nor1213;
logic  invert0215;
logic  nor1214;
logic  invert0216;
logic  nor1215;
logic  invert0217;
logic  nor1216;
logic  invert0218;
logic  nor1217;
logic  invert0219;
logic  nor1218;
logic  invert0220;
logic  nor1219;
logic  invert0221;
logic  nor1220;
logic  invert0222;
logic  nor1221;
logic  invert0223;
logic  nor1222;
logic  invert0224;
logic  nor1223;
logic  invert0225;
logic  nor1224;
logic  invert0226;
logic  nor1225;
logic  invert0227;
logic  nor1226;
logic  invert0228;
logic  nor1227;
logic  invert0229;
logic  nor1228;
logic  invert0230;
logic  nor1229;
logic  invert0231;
logic  nor1230;
logic  invert0232;
logic  nor1231;
logic  invert0233;
logic  nor1232;
logic  invert0234;
logic  nor1233;
logic  invert0235;
logic  nor1234;
logic  invert0236;
logic  nor1235;
logic  invert0237;
logic  nor1236;
logic  invert0238;
logic  nor1237;
logic  invert0239;
logic  nor1238;
logic  invert0240;
logic  nor1239;
logic  invert0241;
logic  nor1240;
logic  invert0242;
logic  nor1241;
logic  invert0243;
logic  nor1242;
logic  invert0244;
logic  nor1243;
logic  invert0245;
logic  nor1244;
logic  invert0246;
logic  nor1245;
logic  invert0247;
logic  nor1246;
logic  invert0248;
logic  nor1247;
logic  invert0249;
logic  nor1248;
logic  invert0250;
logic  nor1249;
logic  invert0251;
logic  nor1250;
logic  invert0252;
logic  nor1251;
logic  invert0253;
logic  nor1252;
logic  invert0254;
logic  nor1253;
logic  invert0255;
logic  nor1254;
logic  invert0256;
logic  nor1255;
logic  invert0257;
logic  nor1256;
logic  invert0258;
logic  nor1257;
logic  invert0259;
logic  nor1258;
logic  invert0260;
logic  nor1259;
logic  invert0261;
logic  nor1260;
logic  invert0262;
logic  nor1261;
logic  invert0263;
logic  nor1262;
logic  invert0264;
logic  nor1263;
logic  invert0265;
logic  nor1264;
logic  invert0266;
logic  nor1265;
logic  invert0267;
logic  nor1266;
logic  invert0268;
logic  nor1267;
logic  invert0269;
logic  nor1268;
logic  invert0270;
logic  nor1269;
logic  invert0271;
logic  nor1270;
logic  invert0272;
logic  nor1271;
logic  invert0273;
logic  nor1272;
logic  invert0274;
logic  nor1273;
logic  invert0275;
logic  nor1274;
logic  invert0276;
logic  nor1275;
logic  invert0277;
logic  nor1276;
logic  invert0278;
logic  nor1277;
logic  invert0279;
logic  nor1278;
logic  invert0280;
logic  nor1279;
logic  invert0281;
logic  nor1280;
logic  invert0282;
logic  nor1281;
logic  invert0283;
logic  nor1282;
logic  invert0284;
logic  nor1283;
logic  invert0285;
logic  nor1284;
logic  invert0286;
logic  nor1285;
logic  invert0287;
logic  nor1286;
logic  invert0288;
logic  nor1287;
logic  invert0289;
logic  nor1288;
logic  invert0290;
logic  nor1289;
logic  invert0291;
logic  nor1290;
logic  invert0292;
logic  nor1291;
logic  invert0293;
logic  nor1292;
logic  invert0294;
logic  nor1293;
logic  invert0295;
logic  nor1294;
logic  invert0296;
logic  nor1295;
logic  invert0297;
logic  nor1296;
logic  invert0298;
logic  nor1297;
logic  invert0299;
logic  nor1298;
logic  invert0300;
logic  nor1299;
logic  invert0301;
logic  nor1300;
logic  invert0302;
logic  nor1301;
logic  invert0303;
logic  nor1302;
logic  invert0304;
logic  nor1303;
logic  invert0305;
logic  nor1304;
logic  invert0306;
logic  nor1305;
logic  invert0307;
logic  nor1306;
logic  invert0308;
logic  nor1307;
logic  invert0309;
logic  nor1308;
logic  invert0310;
logic  nor1309;
logic  invert0311;
logic  nor1310;
logic  invert0312;
logic  nor1311;
logic  invert0313;
logic  nor1312;
logic  invert0314;
logic  nor1313;
logic  invert0315;
logic  nor1314;
logic  invert0316;
logic  nor1315;
logic  invert0317;
logic  nor1316;
logic  invert0318;
logic  nor1317;
logic  invert0319;
logic  nor1318;
logic  invert0320;
logic  nor1319;
logic  invert0321;
logic  nor1320;
logic  invert0322;
logic  nor1321;
logic  invert0323;
logic  nor1322;
logic  invert0324;
logic  nor1323;
logic  invert0325;
logic  nor1324;
logic  invert0326;
logic  nor1325;
logic  invert0327;
logic  nor1326;
logic  invert0328;
logic  nor1327;
logic  invert0329;
logic  nor1328;
logic  invert0330;
logic  nor1329;
logic  invert0331;
logic  nor1330;
logic  invert0332;
logic  nor1331;
logic  invert0333;
logic  nor1332;
logic  invert0334;
logic  nor1333;
logic  invert0335;
logic  nor1334;
logic  invert0336;
logic  nor1335;
logic  invert0337;
logic  nor1336;
logic  invert0338;
logic  nor1337;
logic  invert0339;
logic  nor1338;
logic  invert0340;
logic  nor1339;
logic  invert0341;
logic  nor1340;
logic  invert0342;
logic  nor1341;
logic  invert0343;
logic  nor1342;
logic  invert0344;
logic  nor1343;
logic  invert0345;
logic  nor1344;
logic  invert0346;
logic  nor1345;
logic  invert0347;
logic  nor1346;
logic  invert0348;
logic  nor1347;
logic  invert0349;
logic  nor1348;
logic  invert0350;
logic  nor1349;
logic  invert0351;
logic  nor1350;
logic  invert0352;
logic  nor1351;
logic  invert0353;
logic  nor1352;
logic  invert0354;
logic  nor1353;
logic  invert0355;
logic  nor1354;
logic  invert0356;
logic  nor1355;
logic  invert0357;
logic  nor1356;
logic  invert0358;
logic  nor1357;
logic  invert0359;
logic  nor1358;
logic  invert0360;
logic  nor1359;
logic  invert0361;
logic  nor1360;
logic  invert0362;
logic  nor1361;
logic  invert0363;
logic  nor1362;
logic  invert0364;
logic  nor1363;
logic  invert0365;
logic  nor1364;
logic  invert0366;
logic  nor1365;
logic  invert0367;
logic  nor1366;
logic  invert0368;
logic  nor1367;
logic  invert0369;
logic  nor1368;
logic  invert0370;
logic  nor1369;
logic  invert0371;
logic  nor1370;
logic  invert0372;
logic  nor1371;
logic  invert0373;
logic  nor1372;
logic  invert0374;
logic  nor1373;
logic  invert0375;
logic  nor1374;
logic  invert0376;
logic  nor1375;
logic  invert0377;
logic  nor1376;
logic  invert0378;
logic  nor1377;
logic  invert0379;
logic  nor1378;
logic  invert0380;
logic  nor1379;
logic  invert0381;
logic  nor1380;
logic  invert0382;
logic  nor1381;
logic  invert0383;
logic  nor1382;
logic  invert0384;
logic  nor1383;
logic  invert0385;
logic  nor1384;
logic  invert0386;
logic  nor1385;
logic  invert0387;
logic  nor1386;
logic  invert0388;
logic  nor1387;
logic  invert0389;
logic  nor1388;
logic  invert0390;
logic  nor1389;
logic  invert0391;
logic  nor1390;
logic  invert0392;
logic  nor1391;
logic  invert0393;
logic  nor1392;
logic  invert0394;
logic  nor1393;
logic  invert0395;
logic  nor1394;
logic  invert0396;
logic  nor1395;
logic  invert0397;
logic  nor1396;
logic  invert0398;
logic  nor1397;
logic  invert0399;
logic  nor1398;
logic  invert0400;
logic  nor1399;
logic  invert0401;
logic  nor1400;
logic  invert0402;
logic  nor1401;
logic  invert0403;
logic  nor1402;
logic  invert0404;
logic  nor1403;
logic  invert0405;
logic  nor1404;
logic  invert0406;
logic  nor1405;
logic  invert0407;
logic  nor1406;
logic  invert0408;
logic  nor1407;
logic  invert0409;
logic  nor1408;
logic  invert0410;
logic  nor1409;
logic  invert0411;
logic  nor1410;
logic  invert0412;
logic  nor1411;
logic  invert0413;
logic  nor1412;
logic  invert0414;
logic  nor1413;
logic  invert0415;
logic  nor1414;
logic  invert0416;
logic  nor1415;
logic  invert0417;
logic  nor1416;
logic  invert0418;
logic  nor1417;
logic  invert0419;
logic  nor1418;
logic  invert0420;
logic  nor1419;
logic  invert0421;
logic  nor1420;
logic  invert0422;
logic  nor1421;
logic  invert0423;
logic  nor1422;
logic  invert0424;
logic  nor1423;
logic  invert0425;
logic  nor1424;
logic  invert0426;
logic  nor1425;
logic  invert0427;
logic  nor1426;
logic  invert0428;
logic  nor1427;
logic  invert0429;
logic  nor1428;
logic  invert0430;
logic  nor1429;
logic  invert0431;
logic  nor1430;
logic  invert0432;
logic  nor1431;
logic  invert0433;
logic  nor1432;
logic  invert0434;
logic  nor1433;
logic  invert0435;
logic  nor1434;
logic  invert0436;
logic  nor1435;
logic  invert0437;
logic  nor1436;
logic  invert0438;
logic  nor1437;
logic  invert0439;
logic  nor1438;
logic  invert0440;
logic  nor1439;
logic  invert0441;
logic  nor1440;
logic  invert0442;
logic  nor1441;
logic  invert0443;
logic  nor1442;
logic  invert0444;
logic  nor1443;
logic  invert0445;
logic  nor1444;
logic  invert0446;
logic  nor1445;
logic  invert0447;
logic  nor1446;
logic  invert0448;
logic  nor1447;
logic  invert0449;
logic  nor1448;
logic  invert0450;
logic  nor1449;
logic  invert0451;
logic  nor1450;
logic  invert0452;
logic  nor1451;
logic  invert0453;
logic  nor1452;
logic  invert0454;
logic  nor1453;
logic  invert0455;
logic  nor1454;
logic  invert0456;
logic  nor1455;
logic  invert0457;
logic  nor1456;
logic  invert0458;
logic  nor1457;
logic  invert0459;
logic  nor1458;
logic  invert0460;
logic  nor1459;
logic  invert0461;
logic  nor1460;
logic  invert0462;
logic  nor1461;
logic  invert0463;
logic  nor1462;
logic  invert0464;
logic  nor1463;
logic  invert0465;
logic  nor1464;
logic  invert0466;
logic  nor1465;
logic  invert0467;
logic  nor1466;
logic  invert0468;
logic  nor1467;
logic  invert0469;
logic  nor1468;
logic  invert0470;
logic  nor1469;
logic  invert0471;
logic  nor1470;
logic  invert0472;
logic  nor1471;
logic  invert0473;
logic  nor1472;
logic  invert0474;
logic  nor1473;
logic  invert0475;
logic  nor1474;
logic  invert0476;
logic  nor1475;
logic  invert0477;
logic  nor1476;
logic  invert0478;
logic  nor1477;
logic  invert0479;
logic  nor1478;
logic  invert0480;
logic  nor1479;
logic  invert0481;
logic  nor1480;
logic  invert0482;
logic  nor1481;
logic  invert0483;
logic  nor1482;
logic  invert0484;
logic  nor1483;
logic  invert0485;
logic  nor1484;
logic  invert0486;
logic  nor1485;
logic  invert0487;
logic  nor1486;
logic  invert0488;
logic  nor1487;
logic  invert0489;
logic  nor1488;
logic  invert0490;
logic  nor1489;
logic  invert0491;
logic  nor1490;
logic  invert0492;
logic  nor1491;
logic  invert0493;
logic  nor1492;
logic  invert0494;
logic  nor1493;
logic  invert0495;
logic  nor1494;
logic  invert0496;
logic  nor1495;
logic  invert0497;
logic  nor1496;
logic  invert0498;
logic  nor1497;
logic  invert0499;
logic  nor1498;
logic  invert0500;
logic  nor1499;
logic  invert0501;
logic  nor1500;
logic  invert0502;
logic  nor1501;
logic  invert0503;
logic  nor1502;
logic  invert0504;
logic  nor1503;
logic  invert0505;
logic  nor1504;
logic  invert0506;
logic  nor1505;
logic  invert0507;
logic  nor1506;
logic  invert0508;
logic  nor1507;
logic  invert0509;
logic  nor1508;
logic  invert0510;
logic  nor1509;
logic  invert0511;
logic  nor1510;
logic  invert0512;
logic  nor1511;
logic  invert0513;
logic  nor1512;
logic  invert0514;
logic  nor1513;
logic  invert0515;
logic  nor1514;
logic  invert0516;
logic  nor1515;
logic  invert0517;
logic  nor1516;
logic  invert0518;
logic  nor1517;
logic  invert0519;
logic  nor1518;
logic  invert0520;
logic  nor1519;
logic  invert0521;
logic  nor1520;
logic  invert0522;
logic  nor1521;
logic  invert0523;
logic  nor1522;
logic  invert0524;
logic  nor1523;
logic  invert0525;
logic  nor1524;
logic  invert0526;
logic  nor1525;
logic  invert0527;
logic  nor1526;
logic  invert0528;
logic  nor1527;
logic  invert0529;
logic  nor1528;
logic  invert0530;
logic  nor1529;
logic  invert0531;
logic  nor1530;
logic  invert0532;
logic  nor1531;
logic  invert0533;
logic  nor1532;
logic  invert0534;
logic  nor1533;
logic  invert0535;
logic  nor1534;
logic  invert0536;
logic  nor1535;
logic  invert0537;
logic  nor1536;
logic  invert0538;
logic  nor1537;
logic  invert0539;
logic  nor1538;
logic  invert0540;
logic  nor1539;
logic  invert0541;
logic  nor1540;
logic  invert0542;
logic  nor1541;
logic  invert0543;
logic  nor1542;
logic  invert0544;
logic  nor1543;
logic  invert0545;
logic  nor1544;
logic  invert0546;
logic  nor1545;
logic  invert0547;
logic  nor1546;
logic  invert0548;
logic  nor1547;
logic  invert0549;
logic  nor1548;
logic  invert0550;
logic  nor1549;
logic  invert0551;
logic  nor1550;
logic  invert0552;
logic  nor1551;
logic  invert0553;
logic  nor1552;
logic  invert0554;
logic  nor1553;
logic  invert0555;
logic  nor1554;
logic  invert0556;
logic  nor1555;
logic  invert0557;
logic  nor1556;
logic  invert0558;
logic  nor1557;
logic  invert0559;
logic  nor1558;
logic  invert0560;
logic  nor1559;
logic  invert0561;
logic  nor1560;
logic  invert0562;
logic  nor1561;
logic  invert0563;
logic  nor1562;
logic  invert0564;
logic  nor1563;
logic  invert0565;
logic  nor1564;
logic  invert0566;
logic  nor1565;
logic  invert0567;
logic  nor1566;
logic  invert0568;
logic  nor1567;
logic  invert0569;
logic  nor1568;
logic  invert0570;
logic  nor1569;
logic  invert0571;
logic  nor1570;
logic  invert0572;
logic  nor1571;
logic  invert0573;
logic  nor1572;
logic  invert0574;
logic  nor1573;
logic  invert0575;
logic  nor1574;
logic  invert0576;
logic  nor1575;
logic  invert0577;
logic  nor1576;
logic  invert0578;
logic  nor1577;
logic  invert0579;
logic  nor1578;
logic  invert0580;
logic  nor1579;
logic  invert0581;
logic  nor1580;
logic  invert0582;
logic  nor1581;
logic  invert0583;
logic  nor1582;
logic  invert0584;
logic  nor1583;
logic  invert0585;
logic  nor1584;
logic  invert0586;
logic  nor1585;
logic  invert0587;
logic  nor1586;
logic  invert0588;
logic  nor1587;
logic  invert0589;
logic  nor1588;
logic  invert0590;
logic  nor1589;
logic  invert0591;
logic  nor1590;
logic  invert0592;
logic  nor1591;
logic  invert0593;
logic  nor1592;
logic  invert0594;
logic  nor1593;
logic  invert0595;
logic  nor1594;
logic  invert0596;
logic  nor1595;
logic  invert0597;
logic  nor1596;
logic  invert0598;
logic  nor1597;
logic  invert0599;
logic  nor1598;
logic  invert0600;
logic  nor1599;
logic  invert0601;
logic  nor1600;
logic  invert0602;
logic  nor1601;
logic  invert0603;
logic  nor1602;
logic  invert0604;
logic  nor1603;
logic  invert0605;
logic  nor1604;
logic  invert0606;
logic  nor1605;
logic  invert0607;
logic  nor1606;
logic  invert0608;
logic  nor1607;
logic  invert0609;
logic  nor1608;
logic  invert0610;
logic  nor1609;
logic  invert0611;
logic  nor1610;
logic  invert0612;
logic  nor1611;
logic  invert0613;
logic  nor1612;
logic  invert0614;
logic  nor1613;
logic  invert0615;
logic  nor1614;
logic  invert0616;
logic  nor1615;
logic  invert0617;
logic  nor1616;
logic  invert0618;
logic  nor1617;
logic  invert0619;
logic  nor1618;
logic  invert0620;
logic  nor1619;
logic  invert0621;
logic  nor1620;
logic  invert0622;
logic  nor1621;
logic  invert0623;
logic  nor1622;
logic  invert0624;
logic  nor1623;
logic  invert0625;
logic  nor1624;
logic  invert0626;
logic  nor1625;
logic  invert0627;
logic  nor1626;
logic  invert0628;
logic  nor1627;
logic  invert0629;
logic  nor1628;
logic  invert0630;
logic  nor1629;
logic  invert0631;
logic  nor1630;
logic  invert0632;
logic  nor1631;
logic  invert0633;
logic  nor1632;
logic  invert0634;
logic  nor1633;
logic  invert0635;
logic  nor1634;
logic  invert0636;
logic  nor1635;
logic  invert0637;
logic  nor1636;
logic  invert0638;
logic  nor1637;
logic  invert0639;
logic  nor1638;
logic  invert0640;
logic  nor1639;
logic  invert0641;
logic  nor1640;
logic  invert0642;
logic  nor1641;
logic  invert0643;
logic  nor1642;
logic  invert0644;
logic  nor1643;
logic  invert0645;
logic  nor1644;
logic  invert0646;
logic  nor1645;
logic  invert0647;
logic  nor1646;
logic  invert0648;
logic  nor1647;
logic  invert0649;
logic  nor1648;
logic  invert0650;
logic  nor1649;
logic  invert0651;
logic  nor1650;
logic  invert0652;
logic  nor1651;
logic  invert0653;
logic  nor1652;
logic  invert0654;
logic  nor1653;
logic  invert0655;
logic  nor1654;
logic  invert0656;
logic  nor1655;
logic  invert0657;
logic  nor1656;
logic  invert0658;
logic  nor1657;
logic  invert0659;
logic  nor1658;
logic  invert0660;
logic  nor1659;
logic  invert0661;
logic  nor1660;
logic  invert0662;
logic  nor1661;
logic  invert0663;
logic  nor1662;
logic  invert0664;
logic  nor1663;
logic  invert0665;
logic  nor1664;
logic  invert0666;
logic  nor1665;
logic  invert0667;
logic  nor1666;
logic  invert0668;
logic  nor1667;
logic  invert0669;
logic  nor1668;
logic  invert0670;
logic  nor1669;
logic  invert0671;
logic  nor1670;
logic  invert0672;
logic  nor1671;
logic  invert0673;
logic  nor1672;
logic  invert0674;
logic  nor1673;
logic  invert0675;
logic  nor1674;
logic  invert0676;
logic  nor1675;
logic  invert0677;
logic  nor1676;
logic  invert0678;
logic  nor1677;
logic  invert0679;
logic  nor1678;
logic  invert0680;
logic  nor1679;
logic  invert0681;
logic  nor1680;
logic  invert0682;
logic  nor1681;
logic  invert0683;
logic  nor1682;
logic  invert0684;
logic  nor1683;
logic  invert0685;
logic  nor1684;
logic  invert0686;
logic  nor1685;
logic  invert0687;
logic  nor1686;
logic  invert0688;
logic  nor1687;
logic  invert0689;
logic  nor1688;
logic  invert0690;
logic  nor1689;
logic  invert0691;
logic  nor1690;
logic  invert0692;
logic  nor1691;
logic  invert0693;
logic  nor1692;
logic  invert0694;
logic  nor1693;
logic  invert0695;
logic  nor1694;
logic  invert0696;
logic  nor1695;
logic  invert0697;
logic  nor1696;
logic  invert0698;
logic  nor1697;
logic  invert0699;
logic  nor1698;
logic  invert0700;
logic  nor1699;
logic  invert0701;
logic  nor1700;
logic  invert0702;
logic  nor1701;
logic  invert0703;
logic  nor1702;
logic  invert0704;
logic  nor1703;
logic  invert0705;
logic  nor1704;
logic  invert0706;
logic  nor1705;
logic  invert0707;
logic  nor1706;
logic  invert0708;
logic  nor1707;
logic  invert0709;
logic  nor1708;
logic  invert0710;
logic  nor1709;
logic  invert0711;
logic  nor1710;
logic  invert0712;
logic  nor1711;
logic  invert0713;
logic  nor1712;
logic  invert0714;
logic  nor1713;
logic  invert0715;
logic  nor1714;
logic  invert0716;
logic  nor1715;
logic  invert0717;
logic  nor1716;
logic  invert0718;
logic  nor1717;
logic  invert0719;
logic  nor1718;
logic  invert0720;
logic  nor1719;
logic  invert0721;
logic  nor1720;
logic  invert0722;
logic  nor1721;
logic  invert0723;
logic  nor1722;
logic  invert0724;
logic  nor1723;
logic  invert0725;
logic  nor1724;
logic  invert0726;
logic  nor1725;
logic  invert0727;
logic  nor1726;
logic  invert0728;
logic  nor1727;
logic  invert0729;
logic  nor1728;
logic  invert0730;
logic  nor1729;
logic  invert0731;
logic  nor1730;
logic  invert0732;
logic  nor1731;
logic  invert0733;
logic  nor1732;
logic  invert0734;
logic  nor1733;
logic  invert0735;
logic  nor1734;
logic  invert0736;
logic  nor1735;
logic  invert0737;
logic  nor1736;
logic  invert0738;
logic  nor1737;
logic  invert0739;
logic  nor1738;
logic  invert0740;
logic  nor1739;
logic  invert0741;
logic  nor1740;
logic  invert0742;
logic  nor1741;
logic  invert0743;
logic  nor1742;
logic  invert0744;
logic  nor1743;
logic  invert0745;
logic  nor1744;
logic  invert0746;
logic  nor1745;
logic  invert0747;
logic  nor1746;
logic  invert0748;
logic  nor1747;
logic  invert0749;
logic  nor1748;
logic  invert0750;
logic  nor1749;
logic  invert0751;
logic  nor1750;
logic  invert0752;
logic  nor1751;
logic  invert0753;
logic  nor1752;
logic  invert0754;
logic  nor1753;
logic  invert0755;
logic  nor1754;
logic  invert0756;
logic  nor1755;
logic  invert0757;
logic  nor1756;
logic  invert0758;
logic  nor1757;
logic  invert0759;
logic  nor1758;
logic  invert0760;
logic  nor1759;
logic  invert0761;
logic  nor1760;
logic  invert0762;
logic  nor1761;
logic  invert0763;
logic  nor1762;
logic  invert0764;
logic  nor1763;
logic  invert0765;
logic  nor1764;
logic  invert0766;
logic  nor1765;
logic  invert0767;
logic  nor1766;
logic  invert0768;
logic  nor1767;
logic  invert0769;
logic  nor1768;
logic  invert0770;
logic  nor1769;
logic  invert0771;
logic  nor1770;
logic  invert0772;
logic  nor1771;
logic  invert0773;
logic  nor1772;
logic  invert0774;
logic  nor1773;
logic  invert0775;
logic  nor1774;
logic  invert0776;
logic  nor1775;
logic  invert0777;
logic  nor1776;
logic  invert0778;
logic  nor1777;
logic  invert0779;
logic  nor1778;
logic  invert0780;
logic  nor1779;
logic  invert0781;
logic  nor1780;
logic  invert0782;
logic  nor1781;
logic  invert0783;
logic  nor1782;
logic  invert0784;
logic  nor1783;
logic  invert0785;
logic  nor1784;
logic  invert0786;
logic  nor1785;
logic  invert0787;
logic  nor1786;
logic  invert0788;
logic  nor1787;
logic  invert0789;
logic  nor1788;
logic  invert0790;
logic  nor1789;
logic  invert0791;
logic  nor1790;
logic  invert0792;
logic  nor1791;
logic  invert0793;
logic  nor1792;
logic  invert0794;
logic  nor1793;
logic  invert0795;
logic  nor1794;
logic  invert0796;
logic  nor1795;
logic  invert0797;
logic  nor1796;
logic  invert0798;
logic  nor1797;
logic  invert0799;
logic  nor1798;
logic  invert0800;
logic  nor1799;
logic  invert0801;
logic  nor1800;
logic  invert0802;
logic  nor1801;
logic  invert0803;
logic  nor1802;
logic  invert0804;
logic  nor1803;
logic  invert0805;
logic  nor1804;
logic  invert0806;
logic  nor1805;
logic  invert0807;
logic  nor1806;
logic  invert0808;
logic  nor1807;
logic  invert0809;
logic  nor1808;
logic  invert0810;
logic  nor1809;
logic  invert0811;
logic  nor1810;
logic  invert0812;
logic  nor1811;
logic  invert0813;
logic  nor1812;
logic  invert0814;
logic  nor1813;
logic  invert0815;
logic  nor1814;
logic  invert0816;
logic  nor1815;
logic  invert0817;
logic  nor1816;
logic  invert0818;
logic  nor1817;
logic  invert0819;
logic  nor1818;
logic  invert0820;
logic  nor1819;
logic  invert0821;
logic  nor1820;
logic  invert0822;
logic  nor1821;
logic  invert0823;
logic  nor1822;
logic  invert0824;
logic  nor1823;
logic  invert0825;
logic  nor1824;
logic  invert0826;
logic  nor1825;
logic  invert0827;
logic  nor1826;
logic  invert0828;
logic  nor1827;
logic  invert0829;
logic  nor1828;
logic  invert0830;
logic  nor1829;
logic  invert0831;
logic  nor1830;
logic  invert0832;
logic  nor1831;
logic  invert0833;
logic  nor1832;
logic  invert0834;
logic  nor1833;
logic  invert0835;
logic  nor1834;
logic  invert0836;
logic  nor1835;
logic  invert0837;
logic  nor1836;
logic  invert0838;
logic  nor1837;
logic  invert0839;
logic  nor1838;
logic  invert0840;
logic  nor1839;
logic  invert0841;
logic  nor1840;
logic  invert0842;
logic  nor1841;
logic  invert0843;
logic  nor1842;
logic  invert0844;
logic  nor1843;
logic  invert0845;
logic  nor1844;
logic  invert0846;
logic  nor1845;
logic  invert0847;
logic  nor1846;
logic  invert0848;
logic  nor1847;
logic  invert0849;
logic  nor1848;
logic  invert0850;
logic  nor1849;
logic  invert0851;
logic  nor1850;
logic  invert0852;
logic  nor1851;
logic  invert0853;
logic  nor1852;
logic  invert0854;
logic  nor1853;
logic  invert0855;
logic  nor1854;
logic  invert0856;
logic  nor1855;
logic  invert0857;
logic  nor1856;
logic  invert0858;
logic  nor1857;
logic  invert0859;
logic  nor1858;
logic  invert0860;
logic  nor1859;
logic  invert0861;
logic  nor1860;
logic  invert0862;
logic  nor1861;
logic  invert0863;
logic  nor1862;
logic  invert0864;
logic  nor1863;
logic  invert0865;
logic  nor1864;
logic  invert0866;
logic  nor1865;
logic  invert0867;
logic  nor1866;
logic  invert0868;
logic  nor1867;
logic  invert0869;
logic  nor1868;
logic  invert0870;
logic  nor1869;
logic  invert0871;
logic  nor1870;
logic  invert0872;
logic  nor1871;
logic  invert0873;
logic  nor1872;
logic  invert0874;
logic  nor1873;
logic  invert0875;
logic  nor1874;
logic  invert0876;
logic  nor1875;
logic  invert0877;
logic  nor1876;
logic  invert0878;
logic  nor1877;
logic  invert0879;
logic  nor1878;
logic  invert0880;
logic  nor1879;
logic  invert0881;
logic  nor1880;
logic  invert0882;
logic  nor1881;
logic  invert0883;
logic  nor1882;
logic  invert0884;
logic  nor1883;
logic  invert0885;
logic  nor1884;
logic  invert0886;
logic  nor1885;
logic  invert0887;
logic  nor1886;
logic  invert0888;
logic  nor1887;
logic  invert0889;
logic  nor1888;
logic  invert0890;
logic  nor1889;
logic  invert0891;
logic  nor1890;
logic  invert0892;
logic  nor1891;
logic  invert0893;
logic  nor1892;
logic  invert0894;
logic  nor1893;
logic  invert0895;
logic  nor1894;
logic  invert0896;
logic  nor1895;
logic  invert0897;
logic  nor1896;
logic  invert0898;
logic  nor1897;
logic  invert0899;
logic  nor1898;
logic  invert0900;
logic  nor1899;
logic  invert0901;
logic  nor1900;
logic  invert0902;
logic  nor1901;
logic  invert0903;
logic  nor1902;
logic  invert0904;
logic  nor1903;
logic  invert0905;
logic  nor1904;
logic  invert0906;
logic  nor1905;
logic  invert0907;
logic  nor1906;
logic  invert0908;
logic  nor1907;
logic  invert0909;
logic  nor1908;
logic  invert0910;
logic  nor1909;
logic  invert0911;
logic  nor1910;
logic  invert0912;
logic  nor1911;
logic  invert0913;
logic  nor1912;
logic  invert0914;
logic  nor1913;
logic  invert0915;
logic  nor1914;
logic  invert0916;
logic  nor1915;
logic  invert0917;
logic  nor1916;
logic  invert0918;
logic  nor1917;
logic  invert0919;
logic  nor1918;
logic  invert0920;
logic  nor1919;
logic  invert0921;
logic  nor1920;
logic  invert0922;
logic  nor1921;
logic  invert0923;
logic  nor1922;
logic  invert0924;
logic  nor1923;
logic  invert0925;
logic  nor1924;
logic  invert0926;
logic  nor1925;
logic  invert0927;
logic  nor1926;
logic  invert0928;
logic  nor1927;
logic  invert0929;
logic  nor1928;
logic  invert0930;
logic  nor1929;
logic  invert0931;
logic  nor1930;
logic  invert0932;
logic  nor1931;
logic  invert0933;
logic  nor1932;
logic  invert0934;
logic  nor1933;
logic  invert0935;
logic  nor1934;
logic  invert0936;
logic  nor1935;
logic  invert0937;
logic  nor1936;
logic  invert0938;
logic  nor1937;
logic  invert0939;
logic  nor1938;
logic  invert0940;
logic  nor1939;
logic  invert0941;
logic  nor1940;
logic  invert0942;
logic  nor1941;
logic  invert0943;
logic  nor1942;
logic  invert0944;
logic  nor1943;
logic  invert0945;
logic  nor1944;
logic  invert0946;
logic  nor1945;
logic  invert0947;
logic  nor1946;
logic  invert0948;
logic  nor1947;
logic  invert0949;
logic  nor1948;
logic  invert0950;
logic  nor1949;
logic  invert0951;
logic  nor1950;
logic  invert0952;
logic  nor1951;
logic  invert0953;
logic  nor1952;
logic  invert0954;
logic  nor1953;
logic  invert0955;
logic  nor1954;
logic  invert0956;
logic  nor1955;
logic  invert0957;
logic  nor1956;
logic  invert0958;
logic  nor1957;
logic  invert0959;
logic  nor1958;
logic  invert0960;
logic  nor1959;
logic  invert0961;
logic  nor1960;
logic  invert0962;
logic  nor1961;
logic  invert0963;
logic  nor1962;
logic  invert0964;
logic  nor1963;
logic  invert0965;
logic  nor1964;
logic  invert0966;
logic  nor1965;
logic  invert0967;
logic  nor1966;
logic  invert0968;
logic  nor1967;
logic  invert0969;
logic  nor1968;
logic  invert0970;
logic  nor1969;
logic  invert0971;
logic  nor1970;
logic  invert0972;
logic  nor1971;
logic  invert0973;
logic  nor1972;
logic  invert0974;
logic  nor1973;
logic  invert0975;
logic  nor1974;
logic  invert0976;
logic  nor1975;
logic  invert0977;
logic  nor1976;
logic  invert0978;
logic  nor1977;
logic  invert0979;
logic  nor1978;
logic  invert0980;
logic  nor1979;
logic  invert0981;
logic  nor1980;
logic  invert0982;
logic  nor1981;
logic  invert0983;
logic  nor1982;
logic  invert0984;
logic  nor1983;
logic  invert0985;
logic  nor1984;
logic  invert0986;
logic  nor1985;
logic  invert0987;
logic  nor1986;
logic  invert0988;
logic  nor1987;
logic  invert0989;
logic  nor1988;
logic  invert0990;
logic  nor1989;
logic  invert0991;
logic  nor1990;
logic  invert0992;
logic  nor1991;
logic  invert0993;
logic  nor1992;
logic  invert0994;
logic  nor1993;
logic  invert0995;
logic  nor1994;
logic  invert0996;
logic  nor1995;
logic  invert0997;
logic  nor1996;
logic  invert0998;
logic  nor1997;
logic  invert0999;
logic  nor1998;
logic  invert1000;
logic  nor1999;
logic  invert1001;
logic  nor2000;
logic  invert1002;
logic  nor2001;
logic  invert1003;
logic  nor2002;
logic  invert1004;
logic  nor2003;
logic  invert1005;
logic  nor2004;
logic  invert1006;
logic  nor2005;
logic  invert1007;
logic  nor2006;
logic  invert1008;
logic  nor2007;
logic  invert1009;
logic  nor2008;
logic  invert1010;
logic  nor2009;
logic  invert1011;
logic  nor2010;
logic  invert1012;
logic  nor2011;
logic  invert1013;
logic  nor2012;
logic  invert1014;
logic  nor2013;
logic  invert1015;
logic  nor2014;
logic  invert1016;
logic  nor2015;
logic  invert1017;
logic  nor2016;
logic  invert1018;
logic  nor2017;
logic  invert1019;
logic  nor2018;
logic  invert1020;
logic  nor2019;
logic  invert1021;
logic  nor2020;
logic  invert1022;
logic  nor2021;
logic  invert1023;
// BuildXorTrees
// BuildXorTrees, FirstLevel, f = -1
assign xor0000 = (input_data[0001]^input_data[0000]^input_data[0003]^input_data[0002]); // EmitInputXorGate
assign xor0001 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); // EmitInputXorGate
assign xor0002 = (input_data[0009]^input_data[0008]^input_data[0011]^input_data[0010]); // EmitInputXorGate
assign xor0003 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); // EmitInputXorGate
assign xor0004 = (input_data[0019]^input_data[0018]^input_data[0017]^input_data[0016]); // EmitInputXorGate
assign xor0005 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); // EmitInputXorGate
assign xor0006 = (input_data[0025]^input_data[0024]^input_data[0027]^input_data[0026]); // EmitInputXorGate
assign xor0007 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); // EmitInputXorGate
assign xor0008 = (input_data[0035]^input_data[0034]^input_data[0033]^input_data[0032]); // EmitInputXorGate
assign xor0009 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); // EmitInputXorGate
assign xor0010 = (input_data[0041]^input_data[0040]^input_data[0043]^input_data[0042]); // EmitInputXorGate
assign xor0011 = (input_data[0046]^input_data[0045]^input_data[0044]^input_data[0047]); // EmitInputXorGate
assign xor0012 = (input_data[0051]^input_data[0050]^input_data[0049]^input_data[0048]); // EmitInputXorGate
assign xor0013 = (input_data[0053]^input_data[0052]^input_data[0055]^input_data[0054]); // EmitInputXorGate
assign xor0014 = (input_data[0059]^input_data[0058]^input_data[0057]^input_data[0056]); // EmitInputXorGate
assign xor0015 = (input_data[0063]^input_data[0062]^input_data[0061]^input_data[0060]); // EmitInputXorGate
assign xor0016 = (input_data[0065]^input_data[0064]^input_data[0067]^input_data[0066]); // EmitInputXorGate
assign xor0017 = (input_data[0069]^input_data[0068]^input_data[0071]^input_data[0070]); // EmitInputXorGate
assign xor0018 = (input_data[0072]^input_data[0075]^input_data[0074]^input_data[0073]); // EmitInputXorGate
assign xor0019 = (input_data[0079]^input_data[0078]^input_data[0077]^input_data[0076]); // EmitInputXorGate
assign xor0020 = (input_data[0081]^input_data[0080]^input_data[0083]^input_data[0082]); // EmitInputXorGate
assign xor0021 = (input_data[0085]^input_data[0084]^input_data[0087]^input_data[0086]); // EmitInputXorGate
assign xor0022 = (input_data[0088]^input_data[0091]^input_data[0090]^input_data[0089]); // EmitInputXorGate
assign xor0023 = (input_data[0095]^input_data[0094]^input_data[0093]^input_data[0092]); // EmitInputXorGate
assign xor0024 = (input_data[0097]^input_data[0096]^input_data[0099]^input_data[0098]); // EmitInputXorGate
assign xor0025 = (input_data[0101]^input_data[0100]^input_data[0103]^input_data[0102]); // EmitInputXorGate
assign xor0026 = (input_data[0105]^input_data[0104]^input_data[0107]^input_data[0106]); // EmitInputXorGate
assign xor0027 = (input_data[0111]^input_data[0110]^input_data[0109]^input_data[0108]); // EmitInputXorGate
assign xor0028 = (input_data[0114]^input_data[0113]^input_data[0112]^input_data[0115]); // EmitInputXorGate
assign xor0029 = (input_data[0117]^input_data[0116]^input_data[0119]^input_data[0118]); // EmitInputXorGate
assign xor0030 = (input_data[0121]^input_data[0120]^input_data[0123]^input_data[0122]); // EmitInputXorGate
assign xor0031 = (input_data[0127]^input_data[0126]^input_data[0125]^input_data[0124]); // EmitInputXorGate
assign xor0032 = (input_data[0131]^input_data[0130]^input_data[0129]^input_data[0128]); // EmitInputXorGate
assign xor0033 = (input_data[0133]^input_data[0132]^input_data[0135]^input_data[0134]); // EmitInputXorGate
assign xor0034 = (input_data[0139]^input_data[0138]^input_data[0137]^input_data[0136]); // EmitInputXorGate
assign xor0035 = (input_data[0141]^input_data[0140]^input_data[0143]^input_data[0142]); // EmitInputXorGate
assign xor0036 = (input_data[0145]^input_data[0144]^input_data[0147]^input_data[0146]); // EmitInputXorGate
assign xor0037 = (input_data[0149]^input_data[0148]^input_data[0151]^input_data[0150]); // EmitInputXorGate
assign xor0038 = (input_data[0155]^input_data[0154]^input_data[0153]^input_data[0152]); // EmitInputXorGate
assign xor0039 = (input_data[0159]^input_data[0158]^input_data[0157]^input_data[0156]); // EmitInputXorGate
assign xor0040 = (input_data[0161]^input_data[0160]^input_data[0163]^input_data[0162]); // EmitInputXorGate
assign xor0041 = (input_data[0165]^input_data[0164]^input_data[0167]^input_data[0166]); // EmitInputXorGate
assign xor0042 = (input_data[0169]^input_data[0168]^input_data[0171]^input_data[0170]); // EmitInputXorGate
assign xor0043 = (input_data[0175]^input_data[0174]^input_data[0173]^input_data[0172]); // EmitInputXorGate
assign xor0044 = (input_data[0177]^input_data[0176]^input_data[0179]^input_data[0178]); // EmitInputXorGate
assign xor0045 = (input_data[0181]^input_data[0180]^input_data[0183]^input_data[0182]); // EmitInputXorGate
assign xor0046 = (input_data[0187]^input_data[0186]^input_data[0185]^input_data[0184]); // EmitInputXorGate
assign xor0047 = (input_data[0191]^input_data[0190]^input_data[0189]^input_data[0188]); // EmitInputXorGate
assign xor0048 = (input_data[0193]^input_data[0192]^input_data[0195]^input_data[0194]); // EmitInputXorGate
assign xor0049 = (input_data[0196]^input_data[0199]^input_data[0198]^input_data[0197]); // EmitInputXorGate
assign xor0050 = (input_data[0201]^input_data[0200]^input_data[0203]^input_data[0202]); // EmitInputXorGate
assign xor0051 = (input_data[0205]^input_data[0204]^input_data[0207]^input_data[0206]); // EmitInputXorGate
assign xor0052 = (input_data[0211]^input_data[0210]^input_data[0209]^input_data[0208]); // EmitInputXorGate
assign xor0053 = (input_data[0215]^input_data[0214]^input_data[0213]^input_data[0212]); // EmitInputXorGate
assign xor0054 = (input_data[0217]^input_data[0216]^input_data[0219]^input_data[0218]); // EmitInputXorGate
assign xor0055 = (input_data[0221]^input_data[0220]^input_data[0223]^input_data[0222]); // EmitInputXorGate
assign xor0056 = (input_data[0224]^input_data[0227]^input_data[0226]^input_data[0225]); // EmitInputXorGate
assign xor0057 = (input_data[0231]^input_data[0230]^input_data[0229]^input_data[0228]); // EmitInputXorGate
assign xor0058 = (input_data[0233]^input_data[0232]^input_data[0235]^input_data[0234]); // EmitInputXorGate
assign xor0059 = (input_data[0236]^input_data[0239]^input_data[0238]^input_data[0237]); // EmitInputXorGate
assign xor0060 = (input_data[0242]^input_data[0241]^input_data[0240]^input_data[0243]); // EmitInputXorGate
assign xor0061 = (input_data[0245]^input_data[0244]^input_data[0247]^input_data[0246]); // EmitInputXorGate
assign xor0062 = (input_data[0249]^input_data[0248]^input_data[0251]^input_data[0250]); // EmitInputXorGate
assign xor0063 = (input_data[0255]^input_data[0254]^input_data[0253]^input_data[0252]); // EmitInputXorGate
assign xor0064 = (input_data[0259]^input_data[0258]^input_data[0257]^input_data[0256]); // EmitInputXorGate
assign xor0065 = (input_data[0261]^input_data[0260]^input_data[0263]^input_data[0262]); // EmitInputXorGate
assign xor0066 = (input_data[0265]^input_data[0264]^input_data[0267]^input_data[0266]); // EmitInputXorGate
assign xor0067 = (input_data[0269]^input_data[0268]^input_data[0271]^input_data[0270]); // EmitInputXorGate
assign xor0068 = (input_data[0275]^input_data[0274]^input_data[0273]^input_data[0272]); // EmitInputXorGate
assign xor0069 = (input_data[0278]^input_data[0277]^input_data[0276]^input_data[0279]); // EmitInputXorGate
assign xor0070 = (input_data[0281]^input_data[0280]^input_data[0283]^input_data[0282]); // EmitInputXorGate
assign xor0071 = (input_data[0284]^input_data[0287]^input_data[0286]^input_data[0285]); // EmitInputXorGate
assign xor0072 = (input_data[0291]^input_data[0290]^input_data[0289]^input_data[0288]); // EmitInputXorGate
assign xor0073 = (input_data[0293]^input_data[0292]^input_data[0295]^input_data[0294]); // EmitInputXorGate
assign xor0074 = (input_data[0296]^input_data[0299]^input_data[0298]^input_data[0297]); // EmitInputXorGate
assign xor0075 = (input_data[0301]^input_data[0300]^input_data[0303]^input_data[0302]); // EmitInputXorGate
assign xor0076 = (input_data[0305]^input_data[0304]^input_data[0307]^input_data[0306]); // EmitInputXorGate
assign xor0077 = (input_data[0310]^input_data[0309]^input_data[0308]^input_data[0311]); // EmitInputXorGate
assign xor0078 = (input_data[0313]^input_data[0312]^input_data[0315]^input_data[0314]); // EmitInputXorGate
assign xor0079 = (input_data[0319]^input_data[0318]^input_data[0317]^input_data[0316]); // EmitInputXorGate
assign xor0080 = (input_data[0322]^input_data[0321]^input_data[0320]^input_data[0323]); // EmitInputXorGate
assign xor0081 = (input_data[0325]^input_data[0324]^input_data[0327]^input_data[0326]); // EmitInputXorGate
assign xor0082 = (input_data[0329]^input_data[0328]^input_data[0331]^input_data[0330]); // EmitInputXorGate
assign xor0083 = (input_data[0335]^input_data[0334]^input_data[0333]^input_data[0332]); // EmitInputXorGate
assign xor0084 = (input_data[0339]^input_data[0338]^input_data[0337]^input_data[0336]); // EmitInputXorGate
assign xor0085 = (input_data[0341]^input_data[0340]^input_data[0343]^input_data[0342]); // EmitInputXorGate
assign xor0086 = (input_data[0345]^input_data[0344]^input_data[0347]^input_data[0346]); // EmitInputXorGate
assign xor0087 = (input_data[0348]^input_data[0351]^input_data[0350]^input_data[0349]); // EmitInputXorGate
assign xor0088 = (input_data[0355]^input_data[0354]^input_data[0353]^input_data[0352]); // EmitInputXorGate
assign xor0089 = (input_data[0357]^input_data[0356]^input_data[0359]^input_data[0358]); // EmitInputXorGate
assign xor0090 = (input_data[0361]^input_data[0360]^input_data[0363]^input_data[0362]); // EmitInputXorGate
assign xor0091 = (input_data[0365]^input_data[0364]^input_data[0367]^input_data[0366]); // EmitInputXorGate
assign xor0092 = (input_data[0371]^input_data[0370]^input_data[0369]^input_data[0368]); // EmitInputXorGate
assign xor0093 = (input_data[0373]^input_data[0372]^input_data[0375]^input_data[0374]); // EmitInputXorGate
assign xor0094 = (input_data[0377]^input_data[0376]^input_data[0379]^input_data[0378]); // EmitInputXorGate
assign xor0095 = (input_data[0383]^input_data[0382]^input_data[0381]^input_data[0380]); // EmitInputXorGate
assign xor0096 = (input_data[0385]^input_data[0384]^input_data[0387]^input_data[0386]); // EmitInputXorGate
assign xor0097 = (input_data[0389]^input_data[0388]^input_data[0391]^input_data[0390]); // EmitInputXorGate
assign xor0098 = (input_data[0395]^input_data[0394]^input_data[0393]^input_data[0392]); // EmitInputXorGate
assign xor0099 = (input_data[0399]^input_data[0398]^input_data[0397]^input_data[0396]); // EmitInputXorGate
assign xor0100 = (input_data[0401]^input_data[0400]^input_data[0403]^input_data[0402]); // EmitInputXorGate
assign xor0101 = (input_data[0405]^input_data[0404]^input_data[0407]^input_data[0406]); // EmitInputXorGate
assign xor0102 = (input_data[0411]^input_data[0410]^input_data[0409]^input_data[0408]); // EmitInputXorGate
assign xor0103 = (input_data[0413]^input_data[0412]^input_data[0415]^input_data[0414]); // EmitInputXorGate
assign xor0104 = (input_data[0417]^input_data[0416]^input_data[0419]^input_data[0418]); // EmitInputXorGate
assign xor0105 = (input_data[0421]^input_data[0420]^input_data[0423]^input_data[0422]); // EmitInputXorGate
assign xor0106 = (input_data[0426]^input_data[0425]^input_data[0424]^input_data[0427]); // EmitInputXorGate
assign xor0107 = (input_data[0430]^input_data[0429]^input_data[0428]^input_data[0431]); // EmitInputXorGate
assign xor0108 = (input_data[0433]^input_data[0432]^input_data[0435]^input_data[0434]); // EmitInputXorGate
assign xor0109 = (input_data[0439]^input_data[0438]^input_data[0437]^input_data[0436]); // EmitInputXorGate
assign xor0110 = (input_data[0441]^input_data[0440]^input_data[0443]^input_data[0442]); // EmitInputXorGate
assign xor0111 = (input_data[0445]^input_data[0444]^input_data[0447]^input_data[0446]); // EmitInputXorGate
assign xor0112 = (input_data[0449]^input_data[0448]^input_data[0451]^input_data[0450]); // EmitInputXorGate
assign xor0113 = (input_data[0455]^input_data[0454]^input_data[0453]^input_data[0452]); // EmitInputXorGate
assign xor0114 = (input_data[0459]^input_data[0458]^input_data[0457]^input_data[0456]); // EmitInputXorGate
assign xor0115 = (input_data[0461]^input_data[0460]^input_data[0463]^input_data[0462]); // EmitInputXorGate
assign xor0116 = (input_data[0465]^input_data[0464]^input_data[0467]^input_data[0466]); // EmitInputXorGate
assign xor0117 = (input_data[0468]^input_data[0471]^input_data[0470]^input_data[0469]); // EmitInputXorGate
assign xor0118 = (input_data[0475]^input_data[0474]^input_data[0473]^input_data[0472]); // EmitInputXorGate
assign xor0119 = (input_data[0477]^input_data[0476]^input_data[0479]^input_data[0478]); // EmitInputXorGate
assign xor0120 = (input_data[0481]^input_data[0480]^input_data[0483]^input_data[0482]); // EmitInputXorGate
assign xor0121 = (input_data[0486]^input_data[0485]^input_data[0484]^input_data[0487]); // EmitInputXorGate
assign xor0122 = (input_data[0491]^input_data[0490]^input_data[0489]^input_data[0488]); // EmitInputXorGate
assign xor0123 = (input_data[0493]^input_data[0492]^input_data[0495]^input_data[0494]); // EmitInputXorGate
assign xor0124 = (input_data[0499]^input_data[0498]^input_data[0497]^input_data[0496]); // EmitInputXorGate
assign xor0125 = (input_data[0500]^input_data[0503]^input_data[0502]^input_data[0501]); // EmitInputXorGate
assign xor0126 = (input_data[0505]^input_data[0504]^input_data[0507]^input_data[0506]); // EmitInputXorGate
assign xor0127 = (input_data[0509]^input_data[0508]^input_data[0511]^input_data[0510]); // EmitInputXorGate
assign xor0128 = (input_data[0512]^input_data[0515]^input_data[0514]^input_data[0513]); // EmitInputXorGate
assign xor0129 = (input_data[0519]^input_data[0518]^input_data[0517]^input_data[0516]); // EmitInputXorGate
assign xor0130 = (input_data[0521]^input_data[0520]^input_data[0523]^input_data[0522]); // EmitInputXorGate
assign xor0131 = (input_data[0525]^input_data[0524]^input_data[0527]^input_data[0526]); // EmitInputXorGate
assign xor0132 = (input_data[0529]^input_data[0528]^input_data[0531]^input_data[0530]); // EmitInputXorGate
assign xor0133 = (input_data[0535]^input_data[0534]^input_data[0533]^input_data[0532]); // EmitInputXorGate
assign xor0134 = (input_data[0539]^input_data[0538]^input_data[0537]^input_data[0536]); // EmitInputXorGate
assign xor0135 = (input_data[0541]^input_data[0540]^input_data[0543]^input_data[0542]); // EmitInputXorGate
assign xor0136 = (input_data[0545]^input_data[0544]^input_data[0547]^input_data[0546]); // EmitInputXorGate
assign xor0137 = (input_data[0551]^input_data[0550]^input_data[0549]^input_data[0548]); // EmitInputXorGate
assign xor0138 = (input_data[0554]^input_data[0553]^input_data[0552]^input_data[0555]); // EmitInputXorGate
assign xor0139 = (input_data[0557]^input_data[0556]^input_data[0559]^input_data[0558]); // EmitInputXorGate
assign xor0140 = (input_data[0561]^input_data[0560]^input_data[0563]^input_data[0562]); // EmitInputXorGate
assign xor0141 = (input_data[0567]^input_data[0566]^input_data[0565]^input_data[0564]); // EmitInputXorGate
assign xor0142 = (input_data[0571]^input_data[0570]^input_data[0569]^input_data[0568]); // EmitInputXorGate
assign xor0143 = (input_data[0573]^input_data[0572]^input_data[0575]^input_data[0574]); // EmitInputXorGate
assign xor0144 = (input_data[0579]^input_data[0578]^input_data[0577]^input_data[0576]); // EmitInputXorGate
assign xor0145 = (input_data[0581]^input_data[0580]^input_data[0583]^input_data[0582]); // EmitInputXorGate
assign xor0146 = (input_data[0585]^input_data[0584]^input_data[0587]^input_data[0586]); // EmitInputXorGate
assign xor0147 = (input_data[0589]^input_data[0588]^input_data[0591]^input_data[0590]); // EmitInputXorGate
assign xor0148 = (input_data[0595]^input_data[0594]^input_data[0593]^input_data[0592]); // EmitInputXorGate
assign xor0149 = (input_data[0599]^input_data[0598]^input_data[0597]^input_data[0596]); // EmitInputXorGate
assign xor0150 = (input_data[0601]^input_data[0600]^input_data[0603]^input_data[0602]); // EmitInputXorGate
assign xor0151 = (input_data[0605]^input_data[0604]^input_data[0607]^input_data[0606]); // EmitInputXorGate
assign xor0152 = (input_data[0609]^input_data[0608]^input_data[0611]^input_data[0610]); // EmitInputXorGate
assign xor0153 = (input_data[0613]^input_data[0612]^input_data[0615]^input_data[0614]); // EmitInputXorGate
assign xor0154 = (input_data[0619]^input_data[0618]^input_data[0617]^input_data[0616]); // EmitInputXorGate
assign xor0155 = (input_data[0621]^input_data[0620]^input_data[0623]^input_data[0622]); // EmitInputXorGate
assign xor0156 = (input_data[0625]^input_data[0624]^input_data[0627]^input_data[0626]); // EmitInputXorGate
assign xor0157 = (input_data[0629]^input_data[0628]^input_data[0631]^input_data[0630]); // EmitInputXorGate
assign xor0158 = (input_data[0635]^input_data[0634]^input_data[0633]^input_data[0632]); // EmitInputXorGate
assign xor0159 = (input_data[0639]^input_data[0638]^input_data[0637]^input_data[0636]); // EmitInputXorGate
assign xor0160 = (input_data[0641]^input_data[0640]^input_data[0643]^input_data[0642]); // EmitInputXorGate
assign xor0161 = (input_data[0645]^input_data[0644]^input_data[0647]^input_data[0646]); // EmitInputXorGate
assign xor0162 = (input_data[0651]^input_data[0650]^input_data[0649]^input_data[0648]); // EmitInputXorGate
assign xor0163 = (input_data[0655]^input_data[0654]^input_data[0653]^input_data[0652]); // EmitInputXorGate
assign xor0164 = (input_data[0657]^input_data[0656]^input_data[0659]^input_data[0658]); // EmitInputXorGate
assign xor0165 = (input_data[0661]^input_data[0660]^input_data[0663]^input_data[0662]); // EmitInputXorGate
assign xor0166 = (input_data[0664]^input_data[0667]^input_data[0666]^input_data[0665]); // EmitInputXorGate
assign xor0167 = (input_data[0671]^input_data[0670]^input_data[0669]^input_data[0668]); // EmitInputXorGate
assign xor0168 = (input_data[0673]^input_data[0672]^input_data[0675]^input_data[0674]); // EmitInputXorGate
assign xor0169 = (input_data[0676]^input_data[0679]^input_data[0678]^input_data[0677]); // EmitInputXorGate
assign xor0170 = (input_data[0682]^input_data[0681]^input_data[0680]^input_data[0683]); // EmitInputXorGate
assign xor0171 = (input_data[0685]^input_data[0684]^input_data[0687]^input_data[0686]); // EmitInputXorGate
assign xor0172 = (input_data[0689]^input_data[0688]^input_data[0691]^input_data[0690]); // EmitInputXorGate
assign xor0173 = (input_data[0695]^input_data[0694]^input_data[0693]^input_data[0692]); // EmitInputXorGate
assign xor0174 = (input_data[0699]^input_data[0698]^input_data[0697]^input_data[0696]); // EmitInputXorGate
assign xor0175 = (input_data[0701]^input_data[0700]^input_data[0703]^input_data[0702]); // EmitInputXorGate
assign xor0176 = (input_data[0705]^input_data[0704]^input_data[0707]^input_data[0706]); // EmitInputXorGate
assign xor0177 = (input_data[0709]^input_data[0708]^input_data[0711]^input_data[0710]); // EmitInputXorGate
assign xor0178 = (input_data[0715]^input_data[0714]^input_data[0713]^input_data[0712]); // EmitInputXorGate
assign xor0179 = (input_data[0719]^input_data[0718]^input_data[0717]^input_data[0716]); // EmitInputXorGate
assign xor0180 = (input_data[0721]^input_data[0720]^input_data[0723]^input_data[0722]); // EmitInputXorGate
assign xor0181 = (input_data[0725]^input_data[0724]^input_data[0727]^input_data[0726]); // EmitInputXorGate
assign xor0182 = (input_data[0731]^input_data[0730]^input_data[0729]^input_data[0728]); // EmitInputXorGate
assign xor0183 = (input_data[0735]^input_data[0734]^input_data[0733]^input_data[0732]); // EmitInputXorGate
assign xor0184 = (input_data[0737]^input_data[0736]^input_data[0739]^input_data[0738]); // EmitInputXorGate
assign xor0185 = (input_data[0741]^input_data[0740]^input_data[0743]^input_data[0742]); // EmitInputXorGate
assign xor0186 = (input_data[0745]^input_data[0744]^input_data[0747]^input_data[0746]); // EmitInputXorGate
assign xor0187 = (input_data[0750]^input_data[0749]^input_data[0748]^input_data[0751]); // EmitInputXorGate
assign xor0188 = (input_data[0753]^input_data[0752]^input_data[0755]^input_data[0754]); // EmitInputXorGate
assign xor0189 = (input_data[0759]^input_data[0758]^input_data[0757]^input_data[0756]); // EmitInputXorGate
assign xor0190 = (input_data[0762]^input_data[0761]^input_data[0760]^input_data[0763]); // EmitInputXorGate
assign xor0191 = (input_data[0765]^input_data[0764]^input_data[0767]^input_data[0766]); // EmitInputXorGate
assign xor0192 = (input_data[0769]^input_data[0768]^input_data[0771]^input_data[0770]); // EmitInputXorGate
assign xor0193 = (input_data[0775]^input_data[0774]^input_data[0773]^input_data[0772]); // EmitInputXorGate
assign xor0194 = (input_data[0779]^input_data[0778]^input_data[0777]^input_data[0776]); // EmitInputXorGate
assign xor0195 = (input_data[0781]^input_data[0780]^input_data[0783]^input_data[0782]); // EmitInputXorGate
assign xor0196 = (input_data[0785]^input_data[0784]^input_data[0787]^input_data[0786]); // EmitInputXorGate
assign xor0197 = (input_data[0788]^input_data[0791]^input_data[0790]^input_data[0789]); // EmitInputXorGate
assign xor0198 = (input_data[0795]^input_data[0794]^input_data[0793]^input_data[0792]); // EmitInputXorGate
assign xor0199 = (input_data[0797]^input_data[0796]^input_data[0799]^input_data[0798]); // EmitInputXorGate
assign xor0200 = (input_data[0803]^input_data[0802]^input_data[0801]^input_data[0800]); // EmitInputXorGate
assign xor0201 = (input_data[0805]^input_data[0804]^input_data[0807]^input_data[0806]); // EmitInputXorGate
assign xor0202 = (input_data[0809]^input_data[0808]^input_data[0811]^input_data[0810]); // EmitInputXorGate
assign xor0203 = (input_data[0815]^input_data[0814]^input_data[0813]^input_data[0812]); // EmitInputXorGate
assign xor0204 = (input_data[0819]^input_data[0818]^input_data[0817]^input_data[0816]); // EmitInputXorGate
assign xor0205 = (input_data[0821]^input_data[0820]^input_data[0823]^input_data[0822]); // EmitInputXorGate
assign xor0206 = (input_data[0825]^input_data[0824]^input_data[0827]^input_data[0826]); // EmitInputXorGate
assign xor0207 = (input_data[0829]^input_data[0828]^input_data[0831]^input_data[0830]); // EmitInputXorGate
assign xor0208 = (input_data[0835]^input_data[0834]^input_data[0833]^input_data[0832]); // EmitInputXorGate
assign xor0209 = (input_data[0839]^input_data[0838]^input_data[0837]^input_data[0836]); // EmitInputXorGate
assign xor0210 = (input_data[0841]^input_data[0840]^input_data[0843]^input_data[0842]); // EmitInputXorGate
assign xor0211 = (input_data[0845]^input_data[0844]^input_data[0847]^input_data[0846]); // EmitInputXorGate
assign xor0212 = (input_data[0851]^input_data[0850]^input_data[0849]^input_data[0848]); // EmitInputXorGate
assign xor0213 = (input_data[0853]^input_data[0852]^input_data[0855]^input_data[0854]); // EmitInputXorGate
assign xor0214 = (input_data[0857]^input_data[0856]^input_data[0859]^input_data[0858]); // EmitInputXorGate
assign xor0215 = (input_data[0861]^input_data[0860]^input_data[0863]^input_data[0862]); // EmitInputXorGate
assign xor0216 = (input_data[0866]^input_data[0865]^input_data[0864]^input_data[0867]); // EmitInputXorGate
assign xor0217 = (input_data[0870]^input_data[0869]^input_data[0868]^input_data[0871]); // EmitInputXorGate
assign xor0218 = (input_data[0873]^input_data[0872]^input_data[0875]^input_data[0874]); // EmitInputXorGate
assign xor0219 = (input_data[0879]^input_data[0878]^input_data[0877]^input_data[0876]); // EmitInputXorGate
assign xor0220 = (input_data[0881]^input_data[0880]^input_data[0883]^input_data[0882]); // EmitInputXorGate
assign xor0221 = (input_data[0885]^input_data[0884]^input_data[0887]^input_data[0886]); // EmitInputXorGate
assign xor0222 = (input_data[0889]^input_data[0888]^input_data[0891]^input_data[0890]); // EmitInputXorGate
assign xor0223 = (input_data[0895]^input_data[0894]^input_data[0893]^input_data[0892]); // EmitInputXorGate
assign xor0224 = (input_data[0899]^input_data[0898]^input_data[0897]^input_data[0896]); // EmitInputXorGate
assign xor0225 = (input_data[0901]^input_data[0900]^input_data[0903]^input_data[0902]); // EmitInputXorGate
assign xor0226 = (input_data[0905]^input_data[0904]^input_data[0907]^input_data[0906]); // EmitInputXorGate
assign xor0227 = (input_data[0908]^input_data[0911]^input_data[0910]^input_data[0909]); // EmitInputXorGate
assign xor0228 = (input_data[0915]^input_data[0914]^input_data[0913]^input_data[0912]); // EmitInputXorGate
assign xor0229 = (input_data[0917]^input_data[0916]^input_data[0919]^input_data[0918]); // EmitInputXorGate
assign xor0230 = (input_data[0921]^input_data[0920]^input_data[0923]^input_data[0922]); // EmitInputXorGate
assign xor0231 = (input_data[0925]^input_data[0924]^input_data[0927]^input_data[0926]); // EmitInputXorGate
assign xor0232 = (input_data[0931]^input_data[0930]^input_data[0929]^input_data[0928]); // EmitInputXorGate
assign xor0233 = (input_data[0934]^input_data[0933]^input_data[0932]^input_data[0935]); // EmitInputXorGate
assign xor0234 = (input_data[0937]^input_data[0936]^input_data[0939]^input_data[0938]); // EmitInputXorGate
assign xor0235 = (input_data[0943]^input_data[0942]^input_data[0941]^input_data[0940]); // EmitInputXorGate
assign xor0236 = (input_data[0945]^input_data[0944]^input_data[0947]^input_data[0946]); // EmitInputXorGate
assign xor0237 = (input_data[0949]^input_data[0948]^input_data[0951]^input_data[0950]); // EmitInputXorGate
assign xor0238 = (input_data[0952]^input_data[0955]^input_data[0954]^input_data[0953]); // EmitInputXorGate
assign xor0239 = (input_data[0959]^input_data[0958]^input_data[0957]^input_data[0956]); // EmitInputXorGate
assign xor0240 = (input_data[0961]^input_data[0960]^input_data[0963]^input_data[0962]); // EmitInputXorGate
assign xor0241 = (input_data[0965]^input_data[0964]^input_data[0967]^input_data[0966]); // EmitInputXorGate
assign xor0242 = (input_data[0969]^input_data[0968]^input_data[0971]^input_data[0970]); // EmitInputXorGate
assign xor0243 = (input_data[0975]^input_data[0974]^input_data[0973]^input_data[0972]); // EmitInputXorGate
assign xor0244 = (input_data[0979]^input_data[0978]^input_data[0977]^input_data[0976]); // EmitInputXorGate
assign xor0245 = (input_data[0981]^input_data[0980]^input_data[0983]^input_data[0982]); // EmitInputXorGate
assign xor0246 = (input_data[0985]^input_data[0984]^input_data[0987]^input_data[0986]); // EmitInputXorGate
assign xor0247 = (input_data[0991]^input_data[0990]^input_data[0989]^input_data[0988]); // EmitInputXorGate
assign xor0248 = (input_data[0994]^input_data[0993]^input_data[0992]^input_data[0995]); // EmitInputXorGate
assign xor0249 = (input_data[0997]^input_data[0996]^input_data[0999]^input_data[0998]); // EmitInputXorGate
assign xor0250 = (input_data[1001]^input_data[1000]^input_data[1003]^input_data[1002]); // EmitInputXorGate
assign xor0251 = (input_data[1005]^input_data[1004]^input_data[1007]^input_data[1006]); // EmitInputXorGate
assign xor0252 = (input_data[1008]^input_data[1011]^input_data[1010]^input_data[1009]); // EmitInputXorGate
assign xor0253 = (input_data[1015]^input_data[1014]^input_data[1013]^input_data[1012]); // EmitInputXorGate
assign xor0254 = (input_data[1017]^input_data[1016]^input_data[1019]^input_data[1018]); // EmitInputXorGate
assign xor0255 = (input_data[1021]^input_data[1020]^input_data[1023]^input_data[1022]); // EmitInputXorGate
// BuildXorTrees, FirstLevel, f = 0
assign xor0256 = (input_data[0005]^input_data[0007]^input_data[0001]^input_data[0003]); // EmitInputXorGate
assign xor0257 = (input_data[0009]^input_data[0015]^input_data[0011]^input_data[0013]); // EmitInputXorGate
assign xor0258 = (input_data[0019]^input_data[0017]^input_data[0021]^input_data[0023]); // EmitInputXorGate
assign xor0259 = (input_data[0025]^input_data[0027]^input_data[0031]^input_data[0029]); // EmitInputXorGate
assign xor0260 = (input_data[0035]^input_data[0037]^input_data[0033]^input_data[0039]); // EmitInputXorGate
assign xor0261 = (input_data[0041]^input_data[0043]^input_data[0045]^input_data[0047]); // EmitInputXorGate
assign xor0262 = (input_data[0051]^input_data[0053]^input_data[0049]^input_data[0055]); // EmitInputXorGate
assign xor0263 = (input_data[0063]^input_data[0059]^input_data[0061]^input_data[0057]); // EmitInputXorGate
assign xor0264 = (input_data[0069]^input_data[0065]^input_data[0071]^input_data[0067]); // EmitInputXorGate
assign xor0265 = (input_data[0079]^input_data[0075]^input_data[0077]^input_data[0073]); // EmitInputXorGate
assign xor0266 = (input_data[0085]^input_data[0087]^input_data[0081]^input_data[0083]); // EmitInputXorGate
assign xor0267 = (input_data[0095]^input_data[0091]^input_data[0093]^input_data[0089]); // EmitInputXorGate
assign xor0268 = (input_data[0097]^input_data[0101]^input_data[0103]^input_data[0099]); // EmitInputXorGate
assign xor0269 = (input_data[0105]^input_data[0107]^input_data[0111]^input_data[0109]); // EmitInputXorGate
assign xor0270 = (input_data[0117]^input_data[0113]^input_data[0119]^input_data[0115]); // EmitInputXorGate
assign xor0271 = (input_data[0127]^input_data[0121]^input_data[0123]^input_data[0125]); // EmitInputXorGate
assign xor0272 = (input_data[0131]^input_data[0133]^input_data[0129]^input_data[0135]); // EmitInputXorGate
assign xor0273 = (input_data[0139]^input_data[0141]^input_data[0137]^input_data[0143]); // EmitInputXorGate
assign xor0274 = (input_data[0149]^input_data[0145]^input_data[0147]^input_data[0151]); // EmitInputXorGate
assign xor0275 = (input_data[0159]^input_data[0155]^input_data[0157]^input_data[0153]); // EmitInputXorGate
assign xor0276 = (input_data[0165]^input_data[0167]^input_data[0161]^input_data[0163]); // EmitInputXorGate
assign xor0277 = (input_data[0169]^input_data[0175]^input_data[0171]^input_data[0173]); // EmitInputXorGate
assign xor0278 = (input_data[0181]^input_data[0183]^input_data[0177]^input_data[0179]); // EmitInputXorGate
assign xor0279 = (input_data[0187]^input_data[0191]^input_data[0189]^input_data[0185]); // EmitInputXorGate
assign xor0280 = (input_data[0193]^input_data[0199]^input_data[0195]^input_data[0197]); // EmitInputXorGate
assign xor0281 = (input_data[0205]^input_data[0207]^input_data[0201]^input_data[0203]); // EmitInputXorGate
assign xor0282 = (input_data[0215]^input_data[0211]^input_data[0213]^input_data[0209]); // EmitInputXorGate
assign xor0283 = (input_data[0217]^input_data[0221]^input_data[0223]^input_data[0219]); // EmitInputXorGate
assign xor0284 = (input_data[0231]^input_data[0227]^input_data[0229]^input_data[0225]); // EmitInputXorGate
assign xor0285 = (input_data[0233]^input_data[0239]^input_data[0235]^input_data[0237]); // EmitInputXorGate
assign xor0286 = (input_data[0245]^input_data[0247]^input_data[0241]^input_data[0243]); // EmitInputXorGate
assign xor0287 = (input_data[0249]^input_data[0255]^input_data[0251]^input_data[0253]); // EmitInputXorGate
assign xor0288 = (input_data[0259]^input_data[0257]^input_data[0261]^input_data[0263]); // EmitInputXorGate
assign xor0289 = (input_data[0269]^input_data[0265]^input_data[0267]^input_data[0271]); // EmitInputXorGate
assign xor0290 = (input_data[0275]^input_data[0277]^input_data[0273]^input_data[0279]); // EmitInputXorGate
assign xor0291 = (input_data[0287]^input_data[0281]^input_data[0283]^input_data[0285]); // EmitInputXorGate
assign xor0292 = (input_data[0291]^input_data[0293]^input_data[0289]^input_data[0295]); // EmitInputXorGate
assign xor0293 = (input_data[0301]^input_data[0303]^input_data[0299]^input_data[0297]); // EmitInputXorGate
assign xor0294 = (input_data[0309]^input_data[0305]^input_data[0307]^input_data[0311]); // EmitInputXorGate
assign xor0295 = (input_data[0313]^input_data[0319]^input_data[0315]^input_data[0317]); // EmitInputXorGate
assign xor0296 = (input_data[0325]^input_data[0327]^input_data[0321]^input_data[0323]); // EmitInputXorGate
assign xor0297 = (input_data[0329]^input_data[0335]^input_data[0331]^input_data[0333]); // EmitInputXorGate
assign xor0298 = (input_data[0339]^input_data[0341]^input_data[0343]^input_data[0337]); // EmitInputXorGate
assign xor0299 = (input_data[0345]^input_data[0351]^input_data[0347]^input_data[0349]); // EmitInputXorGate
assign xor0300 = (input_data[0355]^input_data[0357]^input_data[0353]^input_data[0359]); // EmitInputXorGate
assign xor0301 = (input_data[0365]^input_data[0367]^input_data[0361]^input_data[0363]); // EmitInputXorGate
assign xor0302 = (input_data[0371]^input_data[0373]^input_data[0369]^input_data[0375]); // EmitInputXorGate
assign xor0303 = (input_data[0377]^input_data[0383]^input_data[0379]^input_data[0381]); // EmitInputXorGate
assign xor0304 = (input_data[0389]^input_data[0385]^input_data[0387]^input_data[0391]); // EmitInputXorGate
assign xor0305 = (input_data[0399]^input_data[0395]^input_data[0397]^input_data[0393]); // EmitInputXorGate
assign xor0306 = (input_data[0405]^input_data[0407]^input_data[0401]^input_data[0403]); // EmitInputXorGate
assign xor0307 = (input_data[0411]^input_data[0413]^input_data[0409]^input_data[0415]); // EmitInputXorGate
assign xor0308 = (input_data[0417]^input_data[0421]^input_data[0423]^input_data[0419]); // EmitInputXorGate
assign xor0309 = (input_data[0429]^input_data[0425]^input_data[0427]^input_data[0431]); // EmitInputXorGate
assign xor0310 = (input_data[0433]^input_data[0439]^input_data[0435]^input_data[0437]); // EmitInputXorGate
assign xor0311 = (input_data[0445]^input_data[0447]^input_data[0441]^input_data[0443]); // EmitInputXorGate
assign xor0312 = (input_data[0449]^input_data[0455]^input_data[0451]^input_data[0453]); // EmitInputXorGate
assign xor0313 = (input_data[0459]^input_data[0461]^input_data[0457]^input_data[0463]); // EmitInputXorGate
assign xor0314 = (input_data[0465]^input_data[0467]^input_data[0471]^input_data[0469]); // EmitInputXorGate
assign xor0315 = (input_data[0475]^input_data[0477]^input_data[0473]^input_data[0479]); // EmitInputXorGate
assign xor0316 = (input_data[0481]^input_data[0483]^input_data[0485]^input_data[0487]); // EmitInputXorGate
assign xor0317 = (input_data[0491]^input_data[0493]^input_data[0489]^input_data[0495]); // EmitInputXorGate
assign xor0318 = (input_data[0503]^input_data[0499]^input_data[0497]^input_data[0501]); // EmitInputXorGate
assign xor0319 = (input_data[0509]^input_data[0505]^input_data[0507]^input_data[0511]); // EmitInputXorGate
assign xor0320 = (input_data[0519]^input_data[0515]^input_data[0517]^input_data[0513]); // EmitInputXorGate
assign xor0321 = (input_data[0525]^input_data[0527]^input_data[0521]^input_data[0523]); // EmitInputXorGate
assign xor0322 = (input_data[0529]^input_data[0535]^input_data[0531]^input_data[0533]); // EmitInputXorGate
assign xor0323 = (input_data[0539]^input_data[0541]^input_data[0543]^input_data[0537]); // EmitInputXorGate
assign xor0324 = (input_data[0545]^input_data[0551]^input_data[0547]^input_data[0549]); // EmitInputXorGate
assign xor0325 = (input_data[0557]^input_data[0553]^input_data[0559]^input_data[0555]); // EmitInputXorGate
assign xor0326 = (input_data[0567]^input_data[0561]^input_data[0563]^input_data[0565]); // EmitInputXorGate
assign xor0327 = (input_data[0571]^input_data[0573]^input_data[0569]^input_data[0575]); // EmitInputXorGate
assign xor0328 = (input_data[0579]^input_data[0581]^input_data[0577]^input_data[0583]); // EmitInputXorGate
assign xor0329 = (input_data[0589]^input_data[0585]^input_data[0587]^input_data[0591]); // EmitInputXorGate
assign xor0330 = (input_data[0599]^input_data[0595]^input_data[0597]^input_data[0593]); // EmitInputXorGate
assign xor0331 = (input_data[0601]^input_data[0603]^input_data[0605]^input_data[0607]); // EmitInputXorGate
assign xor0332 = (input_data[0613]^input_data[0609]^input_data[0615]^input_data[0611]); // EmitInputXorGate
assign xor0333 = (input_data[0619]^input_data[0621]^input_data[0617]^input_data[0623]); // EmitInputXorGate
assign xor0334 = (input_data[0629]^input_data[0625]^input_data[0627]^input_data[0631]); // EmitInputXorGate
assign xor0335 = (input_data[0639]^input_data[0635]^input_data[0637]^input_data[0633]); // EmitInputXorGate
assign xor0336 = (input_data[0645]^input_data[0647]^input_data[0641]^input_data[0643]); // EmitInputXorGate
assign xor0337 = (input_data[0655]^input_data[0651]^input_data[0653]^input_data[0649]); // EmitInputXorGate
assign xor0338 = (input_data[0657]^input_data[0661]^input_data[0663]^input_data[0659]); // EmitInputXorGate
assign xor0339 = (input_data[0671]^input_data[0667]^input_data[0669]^input_data[0665]); // EmitInputXorGate
assign xor0340 = (input_data[0673]^input_data[0679]^input_data[0675]^input_data[0677]); // EmitInputXorGate
assign xor0341 = (input_data[0685]^input_data[0687]^input_data[0681]^input_data[0683]); // EmitInputXorGate
assign xor0342 = (input_data[0689]^input_data[0695]^input_data[0691]^input_data[0693]); // EmitInputXorGate
assign xor0343 = (input_data[0699]^input_data[0697]^input_data[0701]^input_data[0703]); // EmitInputXorGate
assign xor0344 = (input_data[0709]^input_data[0705]^input_data[0707]^input_data[0711]); // EmitInputXorGate
assign xor0345 = (input_data[0719]^input_data[0715]^input_data[0717]^input_data[0713]); // EmitInputXorGate
assign xor0346 = (input_data[0725]^input_data[0727]^input_data[0721]^input_data[0723]); // EmitInputXorGate
assign xor0347 = (input_data[0735]^input_data[0731]^input_data[0733]^input_data[0729]); // EmitInputXorGate
assign xor0348 = (input_data[0741]^input_data[0743]^input_data[0737]^input_data[0739]); // EmitInputXorGate
assign xor0349 = (input_data[0749]^input_data[0745]^input_data[0747]^input_data[0751]); // EmitInputXorGate
assign xor0350 = (input_data[0753]^input_data[0759]^input_data[0755]^input_data[0757]); // EmitInputXorGate
assign xor0351 = (input_data[0765]^input_data[0767]^input_data[0761]^input_data[0763]); // EmitInputXorGate
assign xor0352 = (input_data[0769]^input_data[0775]^input_data[0771]^input_data[0773]); // EmitInputXorGate
assign xor0353 = (input_data[0779]^input_data[0781]^input_data[0783]^input_data[0777]); // EmitInputXorGate
assign xor0354 = (input_data[0785]^input_data[0791]^input_data[0787]^input_data[0789]); // EmitInputXorGate
assign xor0355 = (input_data[0795]^input_data[0797]^input_data[0793]^input_data[0799]); // EmitInputXorGate
assign xor0356 = (input_data[0803]^input_data[0805]^input_data[0807]^input_data[0801]); // EmitInputXorGate
assign xor0357 = (input_data[0809]^input_data[0815]^input_data[0811]^input_data[0813]); // EmitInputXorGate
assign xor0358 = (input_data[0819]^input_data[0817]^input_data[0821]^input_data[0823]); // EmitInputXorGate
assign xor0359 = (input_data[0829]^input_data[0825]^input_data[0827]^input_data[0831]); // EmitInputXorGate
assign xor0360 = (input_data[0839]^input_data[0835]^input_data[0837]^input_data[0833]); // EmitInputXorGate
assign xor0361 = (input_data[0845]^input_data[0847]^input_data[0841]^input_data[0843]); // EmitInputXorGate
assign xor0362 = (input_data[0851]^input_data[0853]^input_data[0849]^input_data[0855]); // EmitInputXorGate
assign xor0363 = (input_data[0857]^input_data[0861]^input_data[0863]^input_data[0859]); // EmitInputXorGate
assign xor0364 = (input_data[0869]^input_data[0865]^input_data[0867]^input_data[0871]); // EmitInputXorGate
assign xor0365 = (input_data[0873]^input_data[0879]^input_data[0875]^input_data[0877]); // EmitInputXorGate
assign xor0366 = (input_data[0885]^input_data[0887]^input_data[0881]^input_data[0883]); // EmitInputXorGate
assign xor0367 = (input_data[0889]^input_data[0895]^input_data[0891]^input_data[0893]); // EmitInputXorGate
assign xor0368 = (input_data[0899]^input_data[0897]^input_data[0901]^input_data[0903]); // EmitInputXorGate
assign xor0369 = (input_data[0905]^input_data[0907]^input_data[0911]^input_data[0909]); // EmitInputXorGate
assign xor0370 = (input_data[0915]^input_data[0917]^input_data[0913]^input_data[0919]); // EmitInputXorGate
assign xor0371 = (input_data[0925]^input_data[0927]^input_data[0921]^input_data[0923]); // EmitInputXorGate
assign xor0372 = (input_data[0931]^input_data[0933]^input_data[0929]^input_data[0935]); // EmitInputXorGate
assign xor0373 = (input_data[0943]^input_data[0937]^input_data[0939]^input_data[0941]); // EmitInputXorGate
assign xor0374 = (input_data[0949]^input_data[0945]^input_data[0947]^input_data[0951]); // EmitInputXorGate
assign xor0375 = (input_data[0959]^input_data[0955]^input_data[0957]^input_data[0953]); // EmitInputXorGate
assign xor0376 = (input_data[0965]^input_data[0967]^input_data[0961]^input_data[0963]); // EmitInputXorGate
assign xor0377 = (input_data[0969]^input_data[0975]^input_data[0971]^input_data[0973]); // EmitInputXorGate
assign xor0378 = (input_data[0979]^input_data[0981]^input_data[0977]^input_data[0983]); // EmitInputXorGate
assign xor0379 = (input_data[0985]^input_data[0987]^input_data[0991]^input_data[0989]); // EmitInputXorGate
assign xor0380 = (input_data[0997]^input_data[0993]^input_data[0999]^input_data[0995]); // EmitInputXorGate
assign xor0381 = (input_data[1005]^input_data[1007]^input_data[1001]^input_data[1003]); // EmitInputXorGate
assign xor0382 = (input_data[1015]^input_data[1011]^input_data[1013]^input_data[1009]); // EmitInputXorGate
assign xor0383 = (input_data[1017]^input_data[1021]^input_data[1023]^input_data[1019]); // EmitInputXorGate
// BuildXorTrees, FirstLevel, f = 1
assign xor0384 = (input_data[0007]^input_data[0006]^input_data[0003]^input_data[0002]); // EmitInputXorGate
assign xor0385 = (input_data[0015]^input_data[0014]^input_data[0011]^input_data[0010]); // EmitInputXorGate
assign xor0386 = (input_data[0019]^input_data[0018]^input_data[0023]^input_data[0022]); // EmitInputXorGate
assign xor0387 = (input_data[0027]^input_data[0031]^input_data[0030]^input_data[0026]); // EmitInputXorGate
assign xor0388 = (input_data[0035]^input_data[0034]^input_data[0039]^input_data[0038]); // EmitInputXorGate
assign xor0389 = (input_data[0046]^input_data[0043]^input_data[0042]^input_data[0047]); // EmitInputXorGate
assign xor0390 = (input_data[0051]^input_data[0050]^input_data[0055]^input_data[0054]); // EmitInputXorGate
assign xor0391 = (input_data[0063]^input_data[0062]^input_data[0059]^input_data[0058]); // EmitInputXorGate
assign xor0392 = (input_data[0071]^input_data[0067]^input_data[0066]^input_data[0070]); // EmitInputXorGate
assign xor0393 = (input_data[0079]^input_data[0078]^input_data[0075]^input_data[0074]); // EmitInputXorGate
assign xor0394 = (input_data[0087]^input_data[0086]^input_data[0083]^input_data[0082]); // EmitInputXorGate
assign xor0395 = (input_data[0095]^input_data[0094]^input_data[0091]^input_data[0090]); // EmitInputXorGate
assign xor0396 = (input_data[0103]^input_data[0102]^input_data[0099]^input_data[0098]); // EmitInputXorGate
assign xor0397 = (input_data[0107]^input_data[0111]^input_data[0106]^input_data[0110]); // EmitInputXorGate
assign xor0398 = (input_data[0114]^input_data[0119]^input_data[0118]^input_data[0115]); // EmitInputXorGate
assign xor0399 = (input_data[0127]^input_data[0126]^input_data[0123]^input_data[0122]); // EmitInputXorGate
assign xor0400 = (input_data[0131]^input_data[0130]^input_data[0135]^input_data[0134]); // EmitInputXorGate
assign xor0401 = (input_data[0139]^input_data[0138]^input_data[0143]^input_data[0142]); // EmitInputXorGate
assign xor0402 = (input_data[0147]^input_data[0151]^input_data[0150]^input_data[0146]); // EmitInputXorGate
assign xor0403 = (input_data[0159]^input_data[0158]^input_data[0155]^input_data[0154]); // EmitInputXorGate
assign xor0404 = (input_data[0167]^input_data[0166]^input_data[0163]^input_data[0162]); // EmitInputXorGate
assign xor0405 = (input_data[0175]^input_data[0174]^input_data[0171]^input_data[0170]); // EmitInputXorGate
assign xor0406 = (input_data[0183]^input_data[0182]^input_data[0179]^input_data[0178]); // EmitInputXorGate
assign xor0407 = (input_data[0187]^input_data[0186]^input_data[0191]^input_data[0190]); // EmitInputXorGate
assign xor0408 = (input_data[0199]^input_data[0198]^input_data[0195]^input_data[0194]); // EmitInputXorGate
assign xor0409 = (input_data[0207]^input_data[0206]^input_data[0203]^input_data[0202]); // EmitInputXorGate
assign xor0410 = (input_data[0215]^input_data[0214]^input_data[0211]^input_data[0210]); // EmitInputXorGate
assign xor0411 = (input_data[0223]^input_data[0222]^input_data[0219]^input_data[0218]); // EmitInputXorGate
assign xor0412 = (input_data[0231]^input_data[0227]^input_data[0226]^input_data[0230]); // EmitInputXorGate
assign xor0413 = (input_data[0239]^input_data[0238]^input_data[0235]^input_data[0234]); // EmitInputXorGate
assign xor0414 = (input_data[0242]^input_data[0247]^input_data[0246]^input_data[0243]); // EmitInputXorGate
assign xor0415 = (input_data[0255]^input_data[0254]^input_data[0251]^input_data[0250]); // EmitInputXorGate
assign xor0416 = (input_data[0259]^input_data[0258]^input_data[0263]^input_data[0262]); // EmitInputXorGate
assign xor0417 = (input_data[0267]^input_data[0271]^input_data[0266]^input_data[0270]); // EmitInputXorGate
assign xor0418 = (input_data[0278]^input_data[0275]^input_data[0274]^input_data[0279]); // EmitInputXorGate
assign xor0419 = (input_data[0287]^input_data[0286]^input_data[0283]^input_data[0282]); // EmitInputXorGate
assign xor0420 = (input_data[0291]^input_data[0290]^input_data[0295]^input_data[0294]); // EmitInputXorGate
assign xor0421 = (input_data[0303]^input_data[0302]^input_data[0299]^input_data[0298]); // EmitInputXorGate
assign xor0422 = (input_data[0310]^input_data[0307]^input_data[0311]^input_data[0306]); // EmitInputXorGate
assign xor0423 = (input_data[0319]^input_data[0318]^input_data[0315]^input_data[0314]); // EmitInputXorGate
assign xor0424 = (input_data[0322]^input_data[0327]^input_data[0326]^input_data[0323]); // EmitInputXorGate
assign xor0425 = (input_data[0335]^input_data[0334]^input_data[0331]^input_data[0330]); // EmitInputXorGate
assign xor0426 = (input_data[0339]^input_data[0338]^input_data[0343]^input_data[0342]); // EmitInputXorGate
assign xor0427 = (input_data[0351]^input_data[0347]^input_data[0346]^input_data[0350]); // EmitInputXorGate
assign xor0428 = (input_data[0355]^input_data[0354]^input_data[0359]^input_data[0358]); // EmitInputXorGate
assign xor0429 = (input_data[0367]^input_data[0366]^input_data[0363]^input_data[0362]); // EmitInputXorGate
assign xor0430 = (input_data[0371]^input_data[0370]^input_data[0375]^input_data[0374]); // EmitInputXorGate
assign xor0431 = (input_data[0383]^input_data[0382]^input_data[0379]^input_data[0378]); // EmitInputXorGate
assign xor0432 = (input_data[0387]^input_data[0391]^input_data[0386]^input_data[0390]); // EmitInputXorGate
assign xor0433 = (input_data[0399]^input_data[0398]^input_data[0395]^input_data[0394]); // EmitInputXorGate
assign xor0434 = (input_data[0407]^input_data[0406]^input_data[0403]^input_data[0402]); // EmitInputXorGate
assign xor0435 = (input_data[0411]^input_data[0410]^input_data[0415]^input_data[0414]); // EmitInputXorGate
assign xor0436 = (input_data[0423]^input_data[0422]^input_data[0419]^input_data[0418]); // EmitInputXorGate
assign xor0437 = (input_data[0430]^input_data[0426]^input_data[0427]^input_data[0431]); // EmitInputXorGate
assign xor0438 = (input_data[0439]^input_data[0438]^input_data[0435]^input_data[0434]); // EmitInputXorGate
assign xor0439 = (input_data[0447]^input_data[0446]^input_data[0443]^input_data[0442]); // EmitInputXorGate
assign xor0440 = (input_data[0455]^input_data[0454]^input_data[0451]^input_data[0450]); // EmitInputXorGate
assign xor0441 = (input_data[0459]^input_data[0458]^input_data[0463]^input_data[0462]); // EmitInputXorGate
assign xor0442 = (input_data[0467]^input_data[0471]^input_data[0466]^input_data[0470]); // EmitInputXorGate
assign xor0443 = (input_data[0475]^input_data[0474]^input_data[0479]^input_data[0478]); // EmitInputXorGate
assign xor0444 = (input_data[0486]^input_data[0483]^input_data[0482]^input_data[0487]); // EmitInputXorGate
assign xor0445 = (input_data[0491]^input_data[0490]^input_data[0495]^input_data[0494]); // EmitInputXorGate
assign xor0446 = (input_data[0503]^input_data[0502]^input_data[0499]^input_data[0498]); // EmitInputXorGate
assign xor0447 = (input_data[0507]^input_data[0511]^input_data[0506]^input_data[0510]); // EmitInputXorGate
assign xor0448 = (input_data[0519]^input_data[0518]^input_data[0515]^input_data[0514]); // EmitInputXorGate
assign xor0449 = (input_data[0527]^input_data[0526]^input_data[0523]^input_data[0522]); // EmitInputXorGate
assign xor0450 = (input_data[0535]^input_data[0534]^input_data[0531]^input_data[0530]); // EmitInputXorGate
assign xor0451 = (input_data[0539]^input_data[0538]^input_data[0543]^input_data[0542]); // EmitInputXorGate
assign xor0452 = (input_data[0551]^input_data[0547]^input_data[0550]^input_data[0546]); // EmitInputXorGate
assign xor0453 = (input_data[0554]^input_data[0559]^input_data[0558]^input_data[0555]); // EmitInputXorGate
assign xor0454 = (input_data[0567]^input_data[0566]^input_data[0563]^input_data[0562]); // EmitInputXorGate
assign xor0455 = (input_data[0571]^input_data[0570]^input_data[0575]^input_data[0574]); // EmitInputXorGate
assign xor0456 = (input_data[0579]^input_data[0578]^input_data[0583]^input_data[0582]); // EmitInputXorGate
assign xor0457 = (input_data[0587]^input_data[0591]^input_data[0586]^input_data[0590]); // EmitInputXorGate
assign xor0458 = (input_data[0599]^input_data[0598]^input_data[0595]^input_data[0594]); // EmitInputXorGate
assign xor0459 = (input_data[0603]^input_data[0602]^input_data[0607]^input_data[0606]); // EmitInputXorGate
assign xor0460 = (input_data[0615]^input_data[0614]^input_data[0611]^input_data[0610]); // EmitInputXorGate
assign xor0461 = (input_data[0619]^input_data[0618]^input_data[0623]^input_data[0622]); // EmitInputXorGate
assign xor0462 = (input_data[0627]^input_data[0631]^input_data[0626]^input_data[0630]); // EmitInputXorGate
assign xor0463 = (input_data[0639]^input_data[0638]^input_data[0635]^input_data[0634]); // EmitInputXorGate
assign xor0464 = (input_data[0647]^input_data[0646]^input_data[0643]^input_data[0642]); // EmitInputXorGate
assign xor0465 = (input_data[0655]^input_data[0654]^input_data[0651]^input_data[0650]); // EmitInputXorGate
assign xor0466 = (input_data[0663]^input_data[0662]^input_data[0659]^input_data[0658]); // EmitInputXorGate
assign xor0467 = (input_data[0671]^input_data[0667]^input_data[0666]^input_data[0670]); // EmitInputXorGate
assign xor0468 = (input_data[0679]^input_data[0678]^input_data[0675]^input_data[0674]); // EmitInputXorGate
assign xor0469 = (input_data[0682]^input_data[0687]^input_data[0686]^input_data[0683]); // EmitInputXorGate
assign xor0470 = (input_data[0695]^input_data[0694]^input_data[0691]^input_data[0690]); // EmitInputXorGate
assign xor0471 = (input_data[0699]^input_data[0698]^input_data[0703]^input_data[0702]); // EmitInputXorGate
assign xor0472 = (input_data[0707]^input_data[0711]^input_data[0710]^input_data[0706]); // EmitInputXorGate
assign xor0473 = (input_data[0719]^input_data[0718]^input_data[0715]^input_data[0714]); // EmitInputXorGate
assign xor0474 = (input_data[0727]^input_data[0726]^input_data[0723]^input_data[0722]); // EmitInputXorGate
assign xor0475 = (input_data[0735]^input_data[0734]^input_data[0731]^input_data[0730]); // EmitInputXorGate
assign xor0476 = (input_data[0743]^input_data[0742]^input_data[0739]^input_data[0738]); // EmitInputXorGate
assign xor0477 = (input_data[0750]^input_data[0747]^input_data[0751]^input_data[0746]); // EmitInputXorGate
assign xor0478 = (input_data[0759]^input_data[0758]^input_data[0755]^input_data[0754]); // EmitInputXorGate
assign xor0479 = (input_data[0762]^input_data[0767]^input_data[0766]^input_data[0763]); // EmitInputXorGate
assign xor0480 = (input_data[0775]^input_data[0774]^input_data[0771]^input_data[0770]); // EmitInputXorGate
assign xor0481 = (input_data[0779]^input_data[0778]^input_data[0783]^input_data[0782]); // EmitInputXorGate
assign xor0482 = (input_data[0791]^input_data[0787]^input_data[0786]^input_data[0790]); // EmitInputXorGate
assign xor0483 = (input_data[0795]^input_data[0794]^input_data[0799]^input_data[0798]); // EmitInputXorGate
assign xor0484 = (input_data[0803]^input_data[0802]^input_data[0807]^input_data[0806]); // EmitInputXorGate
assign xor0485 = (input_data[0815]^input_data[0814]^input_data[0811]^input_data[0810]); // EmitInputXorGate
assign xor0486 = (input_data[0819]^input_data[0818]^input_data[0823]^input_data[0822]); // EmitInputXorGate
assign xor0487 = (input_data[0827]^input_data[0831]^input_data[0826]^input_data[0830]); // EmitInputXorGate
assign xor0488 = (input_data[0839]^input_data[0838]^input_data[0835]^input_data[0834]); // EmitInputXorGate
assign xor0489 = (input_data[0847]^input_data[0846]^input_data[0843]^input_data[0842]); // EmitInputXorGate
assign xor0490 = (input_data[0851]^input_data[0850]^input_data[0855]^input_data[0854]); // EmitInputXorGate
assign xor0491 = (input_data[0863]^input_data[0862]^input_data[0859]^input_data[0858]); // EmitInputXorGate
assign xor0492 = (input_data[0870]^input_data[0866]^input_data[0867]^input_data[0871]); // EmitInputXorGate
assign xor0493 = (input_data[0879]^input_data[0878]^input_data[0875]^input_data[0874]); // EmitInputXorGate
assign xor0494 = (input_data[0887]^input_data[0886]^input_data[0883]^input_data[0882]); // EmitInputXorGate
assign xor0495 = (input_data[0895]^input_data[0894]^input_data[0891]^input_data[0890]); // EmitInputXorGate
assign xor0496 = (input_data[0899]^input_data[0898]^input_data[0903]^input_data[0902]); // EmitInputXorGate
assign xor0497 = (input_data[0907]^input_data[0911]^input_data[0906]^input_data[0910]); // EmitInputXorGate
assign xor0498 = (input_data[0915]^input_data[0914]^input_data[0919]^input_data[0918]); // EmitInputXorGate
assign xor0499 = (input_data[0927]^input_data[0926]^input_data[0923]^input_data[0922]); // EmitInputXorGate
assign xor0500 = (input_data[0934]^input_data[0931]^input_data[0930]^input_data[0935]); // EmitInputXorGate
assign xor0501 = (input_data[0943]^input_data[0942]^input_data[0939]^input_data[0938]); // EmitInputXorGate
assign xor0502 = (input_data[0947]^input_data[0951]^input_data[0946]^input_data[0950]); // EmitInputXorGate
assign xor0503 = (input_data[0959]^input_data[0958]^input_data[0955]^input_data[0954]); // EmitInputXorGate
assign xor0504 = (input_data[0967]^input_data[0966]^input_data[0963]^input_data[0962]); // EmitInputXorGate
assign xor0505 = (input_data[0975]^input_data[0974]^input_data[0971]^input_data[0970]); // EmitInputXorGate
assign xor0506 = (input_data[0979]^input_data[0978]^input_data[0983]^input_data[0982]); // EmitInputXorGate
assign xor0507 = (input_data[0987]^input_data[0991]^input_data[0990]^input_data[0986]); // EmitInputXorGate
assign xor0508 = (input_data[0994]^input_data[0999]^input_data[0998]^input_data[0995]); // EmitInputXorGate
assign xor0509 = (input_data[1007]^input_data[1006]^input_data[1003]^input_data[1002]); // EmitInputXorGate
assign xor0510 = (input_data[1015]^input_data[1014]^input_data[1011]^input_data[1010]); // EmitInputXorGate
assign xor0511 = (input_data[1023]^input_data[1022]^input_data[1019]^input_data[1018]); // EmitInputXorGate
// BuildXorTrees, FirstLevel, f = 2
assign xor0512 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); // EmitInputXorGate
assign xor0513 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); // EmitInputXorGate
assign xor0514 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); // EmitInputXorGate
assign xor0515 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); // EmitInputXorGate
assign xor0516 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); // EmitInputXorGate
assign xor0517 = (input_data[0046]^input_data[0045]^input_data[0044]^input_data[0047]); // EmitInputXorGate
assign xor0518 = (input_data[0053]^input_data[0052]^input_data[0055]^input_data[0054]); // EmitInputXorGate
assign xor0519 = (input_data[0063]^input_data[0062]^input_data[0061]^input_data[0060]); // EmitInputXorGate
assign xor0520 = (input_data[0069]^input_data[0068]^input_data[0071]^input_data[0070]); // EmitInputXorGate
assign xor0521 = (input_data[0079]^input_data[0078]^input_data[0077]^input_data[0076]); // EmitInputXorGate
assign xor0522 = (input_data[0085]^input_data[0084]^input_data[0087]^input_data[0086]); // EmitInputXorGate
assign xor0523 = (input_data[0095]^input_data[0094]^input_data[0093]^input_data[0092]); // EmitInputXorGate
assign xor0524 = (input_data[0101]^input_data[0100]^input_data[0103]^input_data[0102]); // EmitInputXorGate
assign xor0525 = (input_data[0111]^input_data[0110]^input_data[0109]^input_data[0108]); // EmitInputXorGate
assign xor0526 = (input_data[0117]^input_data[0116]^input_data[0119]^input_data[0118]); // EmitInputXorGate
assign xor0527 = (input_data[0127]^input_data[0126]^input_data[0125]^input_data[0124]); // EmitInputXorGate
assign xor0528 = (input_data[0133]^input_data[0132]^input_data[0135]^input_data[0134]); // EmitInputXorGate
assign xor0529 = (input_data[0141]^input_data[0140]^input_data[0143]^input_data[0142]); // EmitInputXorGate
assign xor0530 = (input_data[0149]^input_data[0148]^input_data[0151]^input_data[0150]); // EmitInputXorGate
assign xor0531 = (input_data[0159]^input_data[0158]^input_data[0157]^input_data[0156]); // EmitInputXorGate
assign xor0532 = (input_data[0165]^input_data[0164]^input_data[0167]^input_data[0166]); // EmitInputXorGate
assign xor0533 = (input_data[0175]^input_data[0174]^input_data[0173]^input_data[0172]); // EmitInputXorGate
assign xor0534 = (input_data[0181]^input_data[0180]^input_data[0183]^input_data[0182]); // EmitInputXorGate
assign xor0535 = (input_data[0191]^input_data[0190]^input_data[0189]^input_data[0188]); // EmitInputXorGate
assign xor0536 = (input_data[0196]^input_data[0199]^input_data[0198]^input_data[0197]); // EmitInputXorGate
assign xor0537 = (input_data[0205]^input_data[0204]^input_data[0207]^input_data[0206]); // EmitInputXorGate
assign xor0538 = (input_data[0215]^input_data[0214]^input_data[0213]^input_data[0212]); // EmitInputXorGate
assign xor0539 = (input_data[0221]^input_data[0220]^input_data[0223]^input_data[0222]); // EmitInputXorGate
assign xor0540 = (input_data[0231]^input_data[0230]^input_data[0229]^input_data[0228]); // EmitInputXorGate
assign xor0541 = (input_data[0236]^input_data[0239]^input_data[0238]^input_data[0237]); // EmitInputXorGate
assign xor0542 = (input_data[0245]^input_data[0244]^input_data[0247]^input_data[0246]); // EmitInputXorGate
assign xor0543 = (input_data[0255]^input_data[0254]^input_data[0253]^input_data[0252]); // EmitInputXorGate
assign xor0544 = (input_data[0261]^input_data[0260]^input_data[0263]^input_data[0262]); // EmitInputXorGate
assign xor0545 = (input_data[0269]^input_data[0268]^input_data[0271]^input_data[0270]); // EmitInputXorGate
assign xor0546 = (input_data[0278]^input_data[0277]^input_data[0276]^input_data[0279]); // EmitInputXorGate
assign xor0547 = (input_data[0284]^input_data[0287]^input_data[0286]^input_data[0285]); // EmitInputXorGate
assign xor0548 = (input_data[0293]^input_data[0292]^input_data[0295]^input_data[0294]); // EmitInputXorGate
assign xor0549 = (input_data[0301]^input_data[0300]^input_data[0303]^input_data[0302]); // EmitInputXorGate
assign xor0550 = (input_data[0310]^input_data[0309]^input_data[0308]^input_data[0311]); // EmitInputXorGate
assign xor0551 = (input_data[0319]^input_data[0318]^input_data[0317]^input_data[0316]); // EmitInputXorGate
assign xor0552 = (input_data[0325]^input_data[0324]^input_data[0327]^input_data[0326]); // EmitInputXorGate
assign xor0553 = (input_data[0335]^input_data[0334]^input_data[0333]^input_data[0332]); // EmitInputXorGate
assign xor0554 = (input_data[0341]^input_data[0340]^input_data[0343]^input_data[0342]); // EmitInputXorGate
assign xor0555 = (input_data[0348]^input_data[0351]^input_data[0350]^input_data[0349]); // EmitInputXorGate
assign xor0556 = (input_data[0357]^input_data[0356]^input_data[0359]^input_data[0358]); // EmitInputXorGate
assign xor0557 = (input_data[0365]^input_data[0364]^input_data[0367]^input_data[0366]); // EmitInputXorGate
assign xor0558 = (input_data[0373]^input_data[0372]^input_data[0375]^input_data[0374]); // EmitInputXorGate
assign xor0559 = (input_data[0383]^input_data[0382]^input_data[0381]^input_data[0380]); // EmitInputXorGate
assign xor0560 = (input_data[0389]^input_data[0388]^input_data[0391]^input_data[0390]); // EmitInputXorGate
assign xor0561 = (input_data[0399]^input_data[0398]^input_data[0397]^input_data[0396]); // EmitInputXorGate
assign xor0562 = (input_data[0405]^input_data[0404]^input_data[0407]^input_data[0406]); // EmitInputXorGate
assign xor0563 = (input_data[0413]^input_data[0412]^input_data[0415]^input_data[0414]); // EmitInputXorGate
assign xor0564 = (input_data[0421]^input_data[0420]^input_data[0423]^input_data[0422]); // EmitInputXorGate
assign xor0565 = (input_data[0430]^input_data[0429]^input_data[0428]^input_data[0431]); // EmitInputXorGate
assign xor0566 = (input_data[0439]^input_data[0438]^input_data[0437]^input_data[0436]); // EmitInputXorGate
assign xor0567 = (input_data[0445]^input_data[0444]^input_data[0447]^input_data[0446]); // EmitInputXorGate
assign xor0568 = (input_data[0455]^input_data[0454]^input_data[0453]^input_data[0452]); // EmitInputXorGate
assign xor0569 = (input_data[0461]^input_data[0460]^input_data[0463]^input_data[0462]); // EmitInputXorGate
assign xor0570 = (input_data[0468]^input_data[0471]^input_data[0470]^input_data[0469]); // EmitInputXorGate
assign xor0571 = (input_data[0477]^input_data[0476]^input_data[0479]^input_data[0478]); // EmitInputXorGate
assign xor0572 = (input_data[0486]^input_data[0485]^input_data[0484]^input_data[0487]); // EmitInputXorGate
assign xor0573 = (input_data[0493]^input_data[0492]^input_data[0495]^input_data[0494]); // EmitInputXorGate
assign xor0574 = (input_data[0500]^input_data[0503]^input_data[0502]^input_data[0501]); // EmitInputXorGate
assign xor0575 = (input_data[0509]^input_data[0508]^input_data[0511]^input_data[0510]); // EmitInputXorGate
assign xor0576 = (input_data[0519]^input_data[0518]^input_data[0517]^input_data[0516]); // EmitInputXorGate
assign xor0577 = (input_data[0525]^input_data[0524]^input_data[0527]^input_data[0526]); // EmitInputXorGate
assign xor0578 = (input_data[0535]^input_data[0534]^input_data[0533]^input_data[0532]); // EmitInputXorGate
assign xor0579 = (input_data[0541]^input_data[0540]^input_data[0543]^input_data[0542]); // EmitInputXorGate
assign xor0580 = (input_data[0551]^input_data[0550]^input_data[0549]^input_data[0548]); // EmitInputXorGate
assign xor0581 = (input_data[0557]^input_data[0556]^input_data[0559]^input_data[0558]); // EmitInputXorGate
assign xor0582 = (input_data[0567]^input_data[0566]^input_data[0565]^input_data[0564]); // EmitInputXorGate
assign xor0583 = (input_data[0573]^input_data[0572]^input_data[0575]^input_data[0574]); // EmitInputXorGate
assign xor0584 = (input_data[0581]^input_data[0580]^input_data[0583]^input_data[0582]); // EmitInputXorGate
assign xor0585 = (input_data[0589]^input_data[0588]^input_data[0591]^input_data[0590]); // EmitInputXorGate
assign xor0586 = (input_data[0599]^input_data[0598]^input_data[0597]^input_data[0596]); // EmitInputXorGate
assign xor0587 = (input_data[0605]^input_data[0604]^input_data[0607]^input_data[0606]); // EmitInputXorGate
assign xor0588 = (input_data[0613]^input_data[0612]^input_data[0615]^input_data[0614]); // EmitInputXorGate
assign xor0589 = (input_data[0621]^input_data[0620]^input_data[0623]^input_data[0622]); // EmitInputXorGate
assign xor0590 = (input_data[0629]^input_data[0628]^input_data[0631]^input_data[0630]); // EmitInputXorGate
assign xor0591 = (input_data[0639]^input_data[0638]^input_data[0637]^input_data[0636]); // EmitInputXorGate
assign xor0592 = (input_data[0645]^input_data[0644]^input_data[0647]^input_data[0646]); // EmitInputXorGate
assign xor0593 = (input_data[0655]^input_data[0654]^input_data[0653]^input_data[0652]); // EmitInputXorGate
assign xor0594 = (input_data[0661]^input_data[0660]^input_data[0663]^input_data[0662]); // EmitInputXorGate
assign xor0595 = (input_data[0671]^input_data[0670]^input_data[0669]^input_data[0668]); // EmitInputXorGate
assign xor0596 = (input_data[0676]^input_data[0679]^input_data[0678]^input_data[0677]); // EmitInputXorGate
assign xor0597 = (input_data[0685]^input_data[0684]^input_data[0687]^input_data[0686]); // EmitInputXorGate
assign xor0598 = (input_data[0695]^input_data[0694]^input_data[0693]^input_data[0692]); // EmitInputXorGate
assign xor0599 = (input_data[0701]^input_data[0700]^input_data[0703]^input_data[0702]); // EmitInputXorGate
assign xor0600 = (input_data[0709]^input_data[0708]^input_data[0711]^input_data[0710]); // EmitInputXorGate
assign xor0601 = (input_data[0719]^input_data[0718]^input_data[0717]^input_data[0716]); // EmitInputXorGate
assign xor0602 = (input_data[0725]^input_data[0724]^input_data[0727]^input_data[0726]); // EmitInputXorGate
assign xor0603 = (input_data[0735]^input_data[0734]^input_data[0733]^input_data[0732]); // EmitInputXorGate
assign xor0604 = (input_data[0741]^input_data[0740]^input_data[0743]^input_data[0742]); // EmitInputXorGate
assign xor0605 = (input_data[0750]^input_data[0749]^input_data[0748]^input_data[0751]); // EmitInputXorGate
assign xor0606 = (input_data[0759]^input_data[0758]^input_data[0757]^input_data[0756]); // EmitInputXorGate
assign xor0607 = (input_data[0765]^input_data[0764]^input_data[0767]^input_data[0766]); // EmitInputXorGate
assign xor0608 = (input_data[0775]^input_data[0774]^input_data[0773]^input_data[0772]); // EmitInputXorGate
assign xor0609 = (input_data[0781]^input_data[0780]^input_data[0783]^input_data[0782]); // EmitInputXorGate
assign xor0610 = (input_data[0788]^input_data[0791]^input_data[0790]^input_data[0789]); // EmitInputXorGate
assign xor0611 = (input_data[0797]^input_data[0796]^input_data[0799]^input_data[0798]); // EmitInputXorGate
assign xor0612 = (input_data[0805]^input_data[0804]^input_data[0807]^input_data[0806]); // EmitInputXorGate
assign xor0613 = (input_data[0815]^input_data[0814]^input_data[0813]^input_data[0812]); // EmitInputXorGate
assign xor0614 = (input_data[0821]^input_data[0820]^input_data[0823]^input_data[0822]); // EmitInputXorGate
assign xor0615 = (input_data[0829]^input_data[0828]^input_data[0831]^input_data[0830]); // EmitInputXorGate
assign xor0616 = (input_data[0839]^input_data[0838]^input_data[0837]^input_data[0836]); // EmitInputXorGate
assign xor0617 = (input_data[0845]^input_data[0844]^input_data[0847]^input_data[0846]); // EmitInputXorGate
assign xor0618 = (input_data[0853]^input_data[0852]^input_data[0855]^input_data[0854]); // EmitInputXorGate
assign xor0619 = (input_data[0861]^input_data[0860]^input_data[0863]^input_data[0862]); // EmitInputXorGate
assign xor0620 = (input_data[0870]^input_data[0869]^input_data[0868]^input_data[0871]); // EmitInputXorGate
assign xor0621 = (input_data[0879]^input_data[0878]^input_data[0877]^input_data[0876]); // EmitInputXorGate
assign xor0622 = (input_data[0885]^input_data[0884]^input_data[0887]^input_data[0886]); // EmitInputXorGate
assign xor0623 = (input_data[0895]^input_data[0894]^input_data[0893]^input_data[0892]); // EmitInputXorGate
assign xor0624 = (input_data[0901]^input_data[0900]^input_data[0903]^input_data[0902]); // EmitInputXorGate
assign xor0625 = (input_data[0908]^input_data[0911]^input_data[0910]^input_data[0909]); // EmitInputXorGate
assign xor0626 = (input_data[0917]^input_data[0916]^input_data[0919]^input_data[0918]); // EmitInputXorGate
assign xor0627 = (input_data[0925]^input_data[0924]^input_data[0927]^input_data[0926]); // EmitInputXorGate
assign xor0628 = (input_data[0934]^input_data[0933]^input_data[0932]^input_data[0935]); // EmitInputXorGate
assign xor0629 = (input_data[0943]^input_data[0942]^input_data[0941]^input_data[0940]); // EmitInputXorGate
assign xor0630 = (input_data[0949]^input_data[0948]^input_data[0951]^input_data[0950]); // EmitInputXorGate
assign xor0631 = (input_data[0959]^input_data[0958]^input_data[0957]^input_data[0956]); // EmitInputXorGate
assign xor0632 = (input_data[0965]^input_data[0964]^input_data[0967]^input_data[0966]); // EmitInputXorGate
assign xor0633 = (input_data[0975]^input_data[0974]^input_data[0973]^input_data[0972]); // EmitInputXorGate
assign xor0634 = (input_data[0981]^input_data[0980]^input_data[0983]^input_data[0982]); // EmitInputXorGate
assign xor0635 = (input_data[0991]^input_data[0990]^input_data[0989]^input_data[0988]); // EmitInputXorGate
assign xor0636 = (input_data[0997]^input_data[0996]^input_data[0999]^input_data[0998]); // EmitInputXorGate
assign xor0637 = (input_data[1005]^input_data[1004]^input_data[1007]^input_data[1006]); // EmitInputXorGate
assign xor0638 = (input_data[1015]^input_data[1014]^input_data[1013]^input_data[1012]); // EmitInputXorGate
assign xor0639 = (input_data[1021]^input_data[1020]^input_data[1023]^input_data[1022]); // EmitInputXorGate
// BuildXorTrees, ParityBits, i = 0
assign xor0640 = (xor0257^xor0258^xor0256^xor0259); // MakeXorFrom
assign xor0641 = (xor0260^xor0263^xor0261^xor0262); // MakeXorFrom
assign xor0642 = (xor0265^xor0266^xor0264^xor0267); // MakeXorFrom
assign xor0643 = (xor0270^xor0268^xor0271^xor0269); // MakeXorFrom
assign xor0644 = (xor0275^xor0273^xor0274^xor0272); // MakeXorFrom
assign xor0645 = (xor0278^xor0276^xor0279^xor0277); // MakeXorFrom
assign xor0646 = (xor0283^xor0281^xor0282^xor0280); // MakeXorFrom
assign xor0647 = (xor0285^xor0286^xor0284^xor0287); // MakeXorFrom
assign xor0648 = (xor0288^xor0291^xor0289^xor0290); // MakeXorFrom
assign xor0649 = (xor0295^xor0293^xor0294^xor0292); // MakeXorFrom
assign xor0650 = (xor0296^xor0299^xor0297^xor0298); // MakeXorFrom
assign xor0651 = (xor0302^xor0300^xor0303^xor0301); // MakeXorFrom
assign xor0652 = (xor0307^xor0305^xor0306^xor0304); // MakeXorFrom
assign xor0653 = (xor0309^xor0310^xor0308^xor0311); // MakeXorFrom
assign xor0654 = (xor0312^xor0315^xor0313^xor0314); // MakeXorFrom
assign xor0655 = (xor0317^xor0318^xor0316^xor0319); // MakeXorFrom
assign xor0656 = (xor0322^xor0320^xor0323^xor0321); // MakeXorFrom
assign xor0657 = (xor0327^xor0325^xor0326^xor0324); // MakeXorFrom
assign xor0658 = (xor0330^xor0328^xor0331^xor0329); // MakeXorFrom
assign xor0659 = (xor0335^xor0333^xor0334^xor0332); // MakeXorFrom
assign xor0660 = (xor0337^xor0338^xor0336^xor0339); // MakeXorFrom
assign xor0661 = (xor0340^xor0343^xor0341^xor0342); // MakeXorFrom
assign xor0662 = (xor0347^xor0345^xor0346^xor0344); // MakeXorFrom
assign xor0663 = (xor0350^xor0348^xor0351^xor0349); // MakeXorFrom
assign xor0664 = (xor0355^xor0353^xor0354^xor0352); // MakeXorFrom
assign xor0665 = (xor0358^xor0356^xor0359^xor0357); // MakeXorFrom
assign xor0666 = (xor0363^xor0361^xor0362^xor0360); // MakeXorFrom
assign xor0667 = (xor0365^xor0366^xor0364^xor0367); // MakeXorFrom
assign xor0668 = (xor0368^xor0371^xor0369^xor0370); // MakeXorFrom
assign xor0669 = (xor0375^xor0373^xor0374^xor0372); // MakeXorFrom
assign xor0670 = (xor0376^xor0379^xor0377^xor0378); // MakeXorFrom
assign xor0671 = (xor0383^xor0381^xor0382^xor0380); // MakeXorFrom
assign xor0672 = (xor0643^xor0641^xor0642^xor0640); // MakeXorFrom
assign xor0673 = (xor0644^xor0647^xor0645^xor0646); // MakeXorFrom
assign xor0674 = (xor0651^xor0649^xor0650^xor0648); // MakeXorFrom
assign xor0675 = (xor0654^xor0652^xor0655^xor0653); // MakeXorFrom
assign xor0676 = (xor0659^xor0657^xor0658^xor0656); // MakeXorFrom
assign xor0677 = (xor0661^xor0662^xor0660^xor0663); // MakeXorFrom
assign xor0678 = (xor0664^xor0667^xor0665^xor0666); // MakeXorFrom
assign xor0679 = (xor0671^xor0669^xor0670^xor0668); // MakeXorFrom
assign xor0680 = (xor0672^xor0675^xor0673^xor0674); // MakeXorFrom
assign xor0681 = (xor0679^xor0677^xor0678^xor0676); // MakeXorFrom
assign xor0682 = (xor0680^xor0681); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 1
assign xor0683 = (xor0386^xor0384^xor0387^xor0385); // MakeXorFrom
assign xor0684 = (xor0391^xor0389^xor0390^xor0388); // MakeXorFrom
assign xor0685 = (xor0393^xor0394^xor0392^xor0395); // MakeXorFrom
assign xor0686 = (xor0396^xor0399^xor0397^xor0398); // MakeXorFrom
assign xor0687 = (xor0403^xor0401^xor0402^xor0400); // MakeXorFrom
assign xor0688 = (xor0404^xor0407^xor0405^xor0406); // MakeXorFrom
assign xor0689 = (xor0411^xor0409^xor0410^xor0408); // MakeXorFrom
assign xor0690 = (xor0414^xor0412^xor0415^xor0413); // MakeXorFrom
assign xor0691 = (xor0419^xor0417^xor0418^xor0416); // MakeXorFrom
assign xor0692 = (xor0421^xor0422^xor0420^xor0423); // MakeXorFrom
assign xor0693 = (xor0424^xor0427^xor0425^xor0426); // MakeXorFrom
assign xor0694 = (xor0431^xor0429^xor0430^xor0428); // MakeXorFrom
assign xor0695 = (xor0434^xor0432^xor0435^xor0433); // MakeXorFrom
assign xor0696 = (xor0439^xor0437^xor0438^xor0436); // MakeXorFrom
assign xor0697 = (xor0441^xor0442^xor0440^xor0443); // MakeXorFrom
assign xor0698 = (xor0447^xor0445^xor0446^xor0444); // MakeXorFrom
assign xor0699 = (xor0449^xor0450^xor0448^xor0451); // MakeXorFrom
assign xor0700 = (xor0452^xor0455^xor0453^xor0454); // MakeXorFrom
assign xor0701 = (xor0459^xor0457^xor0458^xor0456); // MakeXorFrom
assign xor0702 = (xor0462^xor0460^xor0463^xor0461); // MakeXorFrom
assign xor0703 = (xor0467^xor0465^xor0466^xor0464); // MakeXorFrom
assign xor0704 = (xor0470^xor0468^xor0471^xor0469); // MakeXorFrom
assign xor0705 = (xor0475^xor0473^xor0474^xor0472); // MakeXorFrom
assign xor0706 = (xor0477^xor0478^xor0476^xor0479); // MakeXorFrom
assign xor0707 = (xor0480^xor0483^xor0481^xor0482); // MakeXorFrom
assign xor0708 = (xor0487^xor0485^xor0486^xor0484); // MakeXorFrom
assign xor0709 = (xor0490^xor0488^xor0491^xor0489); // MakeXorFrom
assign xor0710 = (xor0495^xor0493^xor0494^xor0492); // MakeXorFrom
assign xor0711 = (xor0498^xor0496^xor0499^xor0497); // MakeXorFrom
assign xor0712 = (xor0501^xor0502^xor0500^xor0503); // MakeXorFrom
assign xor0713 = (xor0504^xor0507^xor0505^xor0506); // MakeXorFrom
assign xor0714 = (xor0511^xor0509^xor0510^xor0508); // MakeXorFrom
assign xor0715 = (xor0685^xor0686^xor0683^xor0684); // MakeXorFrom
assign xor0716 = (xor0689^xor0690^xor0687^xor0688); // MakeXorFrom
assign xor0717 = (xor0692^xor0693^xor0694^xor0691); // MakeXorFrom
assign xor0718 = (xor0697^xor0698^xor0695^xor0696); // MakeXorFrom
assign xor0719 = (xor0701^xor0702^xor0700^xor0699); // MakeXorFrom
assign xor0720 = (xor0706^xor0703^xor0704^xor0705); // MakeXorFrom
assign xor0721 = (xor0709^xor0710^xor0707^xor0708); // MakeXorFrom
assign xor0722 = (xor0713^xor0714^xor0711^xor0712); // MakeXorFrom
assign xor0723 = (xor0716^xor0717^xor0718^xor0715); // MakeXorFrom
assign xor0724 = (xor0721^xor0722^xor0719^xor0720); // MakeXorFrom
assign xor0725 = (xor0723^xor0724); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 2
assign xor0726 = (xor0514^xor0512^xor0515^xor0513); // MakeXorFrom
assign xor0727 = (xor0519^xor0517^xor0518^xor0516); // MakeXorFrom
assign xor0728 = (xor0521^xor0522^xor0520^xor0523); // MakeXorFrom
assign xor0729 = (xor0527^xor0525^xor0526^xor0524); // MakeXorFrom
assign xor0730 = (xor0529^xor0530^xor0528^xor0531); // MakeXorFrom
assign xor0731 = (xor0532^xor0535^xor0533^xor0534); // MakeXorFrom
assign xor0732 = (xor0539^xor0537^xor0538^xor0536); // MakeXorFrom
assign xor0733 = (xor0542^xor0540^xor0543^xor0541); // MakeXorFrom
assign xor0734 = (xor0547^xor0545^xor0546^xor0544); // MakeXorFrom
assign xor0735 = (xor0550^xor0548^xor0551^xor0549); // MakeXorFrom
assign xor0736 = (xor0552^xor0555^xor0553^xor0554); // MakeXorFrom
assign xor0737 = (xor0557^xor0558^xor0556^xor0559); // MakeXorFrom
assign xor0738 = (xor0560^xor0563^xor0561^xor0562); // MakeXorFrom
assign xor0739 = (xor0567^xor0565^xor0566^xor0564); // MakeXorFrom
assign xor0740 = (xor0570^xor0568^xor0571^xor0569); // MakeXorFrom
assign xor0741 = (xor0575^xor0573^xor0574^xor0572); // MakeXorFrom
assign xor0742 = (xor0577^xor0578^xor0576^xor0579); // MakeXorFrom
assign xor0743 = (xor0580^xor0583^xor0581^xor0582); // MakeXorFrom
assign xor0744 = (xor0585^xor0586^xor0584^xor0587); // MakeXorFrom
assign xor0745 = (xor0588^xor0591^xor0589^xor0590); // MakeXorFrom
assign xor0746 = (xor0595^xor0593^xor0594^xor0592); // MakeXorFrom
assign xor0747 = (xor0598^xor0596^xor0599^xor0597); // MakeXorFrom
assign xor0748 = (xor0603^xor0601^xor0602^xor0600); // MakeXorFrom
assign xor0749 = (xor0605^xor0606^xor0604^xor0607); // MakeXorFrom
assign xor0750 = (xor0611^xor0609^xor0610^xor0608); // MakeXorFrom
assign xor0751 = (xor0613^xor0614^xor0612^xor0615); // MakeXorFrom
assign xor0752 = (xor0616^xor0619^xor0617^xor0618); // MakeXorFrom
assign xor0753 = (xor0623^xor0621^xor0622^xor0620); // MakeXorFrom
assign xor0754 = (xor0626^xor0624^xor0627^xor0625); // MakeXorFrom
assign xor0755 = (xor0631^xor0629^xor0630^xor0628); // MakeXorFrom
assign xor0756 = (xor0633^xor0634^xor0632^xor0635); // MakeXorFrom
assign xor0757 = (xor0639^xor0637^xor0638^xor0636); // MakeXorFrom
assign xor0758 = (xor0729^xor0727^xor0728^xor0726); // MakeXorFrom
assign xor0759 = (xor0731^xor0732^xor0730^xor0733); // MakeXorFrom
assign xor0760 = (xor0734^xor0737^xor0735^xor0736); // MakeXorFrom
assign xor0761 = (xor0741^xor0739^xor0740^xor0738); // MakeXorFrom
assign xor0762 = (xor0744^xor0742^xor0745^xor0743); // MakeXorFrom
assign xor0763 = (xor0749^xor0747^xor0748^xor0746); // MakeXorFrom
assign xor0764 = (xor0751^xor0752^xor0750^xor0753); // MakeXorFrom
assign xor0765 = (xor0757^xor0755^xor0756^xor0754); // MakeXorFrom
assign xor0766 = (xor0761^xor0759^xor0760^xor0758); // MakeXorFrom
assign xor0767 = (xor0762^xor0765^xor0763^xor0764); // MakeXorFrom
assign xor0768 = (xor0767^xor0766); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 3
assign xor0769 = (xor0002^xor0010^xor0006^xor0014); // MakeXorFrom
assign xor0770 = (xor0030^xor0018^xor0026^xor0022); // MakeXorFrom
assign xor0771 = (xor0038^xor0046^xor0034^xor0042); // MakeXorFrom
assign xor0772 = (xor0054^xor0062^xor0058^xor0050); // MakeXorFrom
assign xor0773 = (xor0066^xor0074^xor0078^xor0070); // MakeXorFrom
assign xor0774 = (xor0086^xor0094^xor0082^xor0090); // MakeXorFrom
assign xor0775 = (xor0110^xor0106^xor0098^xor0102); // MakeXorFrom
assign xor0776 = (xor0118^xor0126^xor0114^xor0122); // MakeXorFrom
assign xor0777 = (xor0138^xor0134^xor0142^xor0130); // MakeXorFrom
assign xor0778 = (xor0146^xor0154^xor0150^xor0158); // MakeXorFrom
assign xor0779 = (xor0166^xor0174^xor0162^xor0170); // MakeXorFrom
assign xor0780 = (xor0182^xor0190^xor0178^xor0186); // MakeXorFrom
assign xor0781 = (xor0194^xor0202^xor0198^xor0206); // MakeXorFrom
assign xor0782 = (xor0222^xor0210^xor0218^xor0214); // MakeXorFrom
assign xor0783 = (xor0230^xor0238^xor0226^xor0234); // MakeXorFrom
assign xor0784 = (xor0250^xor0246^xor0254^xor0242); // MakeXorFrom
assign xor0785 = (xor0519^xor0517^xor0515^xor0513); // MakeXorFrom
assign xor0786 = (xor0521^xor0527^xor0525^xor0523); // MakeXorFrom
assign xor0787 = (xor0529^xor0535^xor0533^xor0531); // MakeXorFrom
assign xor0788 = (xor0539^xor0537^xor0543^xor0541); // MakeXorFrom
assign xor0789 = (xor0547^xor0545^xor0551^xor0549); // MakeXorFrom
assign xor0790 = (xor0557^xor0555^xor0553^xor0559); // MakeXorFrom
assign xor0791 = (xor0567^xor0565^xor0563^xor0561); // MakeXorFrom
assign xor0792 = (xor0575^xor0573^xor0571^xor0569); // MakeXorFrom
assign xor0793 = (xor0577^xor0583^xor0581^xor0579); // MakeXorFrom
assign xor0794 = (xor0585^xor0591^xor0589^xor0587); // MakeXorFrom
assign xor0795 = (xor0595^xor0593^xor0599^xor0597); // MakeXorFrom
assign xor0796 = (xor0605^xor0603^xor0601^xor0607); // MakeXorFrom
assign xor0797 = (xor0613^xor0611^xor0609^xor0615); // MakeXorFrom
assign xor0798 = (xor0623^xor0621^xor0619^xor0617); // MakeXorFrom
assign xor0799 = (xor0631^xor0629^xor0627^xor0625); // MakeXorFrom
assign xor0800 = (xor0633^xor0639^xor0637^xor0635); // MakeXorFrom
assign xor0801 = (xor0769^xor0772^xor0770^xor0771); // MakeXorFrom
assign xor0802 = (xor0775^xor0776^xor0773^xor0774); // MakeXorFrom
assign xor0803 = (xor0777^xor0780^xor0778^xor0779); // MakeXorFrom
assign xor0804 = (xor0782^xor0783^xor0784^xor0781); // MakeXorFrom
assign xor0805 = (xor0787^xor0788^xor0785^xor0786); // MakeXorFrom
assign xor0806 = (xor0790^xor0791^xor0789^xor0792); // MakeXorFrom
assign xor0807 = (xor0795^xor0796^xor0793^xor0794); // MakeXorFrom
assign xor0808 = (xor0800^xor0797^xor0798^xor0799); // MakeXorFrom
assign xor0809 = (xor0803^xor0804^xor0801^xor0802); // MakeXorFrom
assign xor0810 = (xor0808^xor0805^xor0806^xor0807); // MakeXorFrom
assign xor0811 = (xor0810^xor0809); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 4
assign xor0812 = (xor0006^xor0014^xor0004^xor0012); // MakeXorFrom
assign xor0813 = (xor0030^xor0020^xor0028^xor0022); // MakeXorFrom
assign xor0814 = (xor0038^xor0046^xor0036^xor0044); // MakeXorFrom
assign xor0815 = (xor0054^xor0062^xor0052^xor0060); // MakeXorFrom
assign xor0816 = (xor0076^xor0078^xor0070^xor0068); // MakeXorFrom
assign xor0817 = (xor0086^xor0094^xor0084^xor0092); // MakeXorFrom
assign xor0818 = (xor0110^xor0100^xor0108^xor0102); // MakeXorFrom
assign xor0819 = (xor0118^xor0126^xor0116^xor0124); // MakeXorFrom
assign xor0820 = (xor0134^xor0142^xor0132^xor0140); // MakeXorFrom
assign xor0821 = (xor0156^xor0150^xor0158^xor0148); // MakeXorFrom
assign xor0822 = (xor0166^xor0174^xor0164^xor0172); // MakeXorFrom
assign xor0823 = (xor0182^xor0190^xor0180^xor0188); // MakeXorFrom
assign xor0824 = (xor0204^xor0198^xor0206^xor0196); // MakeXorFrom
assign xor0825 = (xor0222^xor0212^xor0220^xor0214); // MakeXorFrom
assign xor0826 = (xor0230^xor0238^xor0228^xor0236); // MakeXorFrom
assign xor0827 = (xor0246^xor0254^xor0244^xor0252); // MakeXorFrom
assign xor0828 = (xor0514^xor0519^xor0518^xor0515); // MakeXorFrom
assign xor0829 = (xor0522^xor0527^xor0526^xor0523); // MakeXorFrom
assign xor0830 = (xor0530^xor0535^xor0534^xor0531); // MakeXorFrom
assign xor0831 = (xor0539^xor0542^xor0538^xor0543); // MakeXorFrom
assign xor0832 = (xor0550^xor0547^xor0546^xor0551); // MakeXorFrom
assign xor0833 = (xor0558^xor0555^xor0554^xor0559); // MakeXorFrom
assign xor0834 = (xor0567^xor0566^xor0563^xor0562); // MakeXorFrom
assign xor0835 = (xor0570^xor0575^xor0574^xor0571); // MakeXorFrom
assign xor0836 = (xor0578^xor0583^xor0579^xor0582); // MakeXorFrom
assign xor0837 = (xor0586^xor0591^xor0590^xor0587); // MakeXorFrom
assign xor0838 = (xor0598^xor0595^xor0594^xor0599); // MakeXorFrom
assign xor0839 = (xor0606^xor0603^xor0602^xor0607); // MakeXorFrom
assign xor0840 = (xor0614^xor0611^xor0610^xor0615); // MakeXorFrom
assign xor0841 = (xor0623^xor0619^xor0622^xor0618); // MakeXorFrom
assign xor0842 = (xor0626^xor0631^xor0630^xor0627); // MakeXorFrom
assign xor0843 = (xor0634^xor0639^xor0638^xor0635); // MakeXorFrom
assign xor0844 = (xor0815^xor0813^xor0814^xor0812); // MakeXorFrom
assign xor0845 = (xor0818^xor0816^xor0819^xor0817); // MakeXorFrom
assign xor0846 = (xor0823^xor0821^xor0822^xor0820); // MakeXorFrom
assign xor0847 = (xor0825^xor0826^xor0824^xor0827); // MakeXorFrom
assign xor0848 = (xor0828^xor0831^xor0829^xor0830); // MakeXorFrom
assign xor0849 = (xor0835^xor0833^xor0834^xor0832); // MakeXorFrom
assign xor0850 = (xor0836^xor0839^xor0837^xor0838); // MakeXorFrom
assign xor0851 = (xor0843^xor0841^xor0842^xor0840); // MakeXorFrom
assign xor0852 = (xor0846^xor0844^xor0847^xor0845); // MakeXorFrom
assign xor0853 = (xor0851^xor0849^xor0850^xor0848); // MakeXorFrom
assign xor0854 = (xor0853^xor0852); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 5
assign xor0855 = (xor0010^xor0008^xor0014^xor0012); // MakeXorFrom
assign xor0856 = (xor0030^xor0028^xor0026^xor0024); // MakeXorFrom
assign xor0857 = (xor0040^xor0046^xor0044^xor0042); // MakeXorFrom
assign xor0858 = (xor0056^xor0062^xor0060^xor0058); // MakeXorFrom
assign xor0859 = (xor0076^xor0074^xor0072^xor0078); // MakeXorFrom
assign xor0860 = (xor0094^xor0092^xor0090^xor0088); // MakeXorFrom
assign xor0861 = (xor0110^xor0108^xor0106^xor0104); // MakeXorFrom
assign xor0862 = (xor0120^xor0126^xor0124^xor0122); // MakeXorFrom
assign xor0863 = (xor0138^xor0136^xor0142^xor0140); // MakeXorFrom
assign xor0864 = (xor0156^xor0154^xor0152^xor0158); // MakeXorFrom
assign xor0865 = (xor0174^xor0172^xor0170^xor0168); // MakeXorFrom
assign xor0866 = (xor0184^xor0190^xor0188^xor0186); // MakeXorFrom
assign xor0867 = (xor0204^xor0202^xor0200^xor0206); // MakeXorFrom
assign xor0868 = (xor0222^xor0220^xor0218^xor0216); // MakeXorFrom
assign xor0869 = (xor0232^xor0238^xor0236^xor0234); // MakeXorFrom
assign xor0870 = (xor0250^xor0248^xor0254^xor0252); // MakeXorFrom
assign xor0871 = (xor0731^xor0729^xor0727^xor0733); // MakeXorFrom
assign xor0872 = (xor0741^xor0739^xor0737^xor0735); // MakeXorFrom
assign xor0873 = (xor0749^xor0747^xor0745^xor0743); // MakeXorFrom
assign xor0874 = (xor0751^xor0757^xor0755^xor0753); // MakeXorFrom
assign xor0875 = (xor0856^xor0857^xor0858^xor0855); // MakeXorFrom
assign xor0876 = (xor0861^xor0859^xor0862^xor0860); // MakeXorFrom
assign xor0877 = (xor0863^xor0864^xor0865^xor0866); // MakeXorFrom
assign xor0878 = (xor0869^xor0867^xor0870^xor0868); // MakeXorFrom
assign xor0879 = (xor0873^xor0874^xor0871^xor0872); // MakeXorFrom
assign xor0880 = (xor0877^xor0878^xor0875^xor0876); // MakeXorFrom
assign xor0881 = xor0879;
assign xor0882 = (xor0881^xor0880); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 6
assign xor0883 = (xor0020^xor0018^xor0016^xor0022); // MakeXorFrom
assign xor0884 = (xor0048^xor0054^xor0052^xor0050); // MakeXorFrom
assign xor0885 = (xor0086^xor0084^xor0082^xor0080); // MakeXorFrom
assign xor0886 = (xor0118^xor0116^xor0114^xor0112); // MakeXorFrom
assign xor0887 = (xor0146^xor0144^xor0150^xor0148); // MakeXorFrom
assign xor0888 = (xor0176^xor0182^xor0180^xor0178); // MakeXorFrom
assign xor0889 = (xor0212^xor0210^xor0208^xor0214); // MakeXorFrom
assign xor0890 = (xor0240^xor0246^xor0244^xor0242); // MakeXorFrom
assign xor0891 = (xor0521^xor0520^xor0525^xor0524); // MakeXorFrom
assign xor0892 = (xor0537^xor0540^xor0536^xor0541); // MakeXorFrom
assign xor0893 = (xor0552^xor0557^xor0556^xor0553); // MakeXorFrom
assign xor0894 = (xor0568^xor0573^xor0569^xor0572); // MakeXorFrom
assign xor0895 = (xor0588^xor0585^xor0584^xor0589); // MakeXorFrom
assign xor0896 = (xor0605^xor0604^xor0601^xor0600); // MakeXorFrom
assign xor0897 = (xor0616^xor0621^xor0617^xor0620); // MakeXorFrom
assign xor0898 = (xor0633^xor0632^xor0637^xor0636); // MakeXorFrom
assign xor0899 = (xor0835^xor0833^xor0831^xor0829); // MakeXorFrom
assign xor0900 = (xor0843^xor0841^xor0839^xor0837); // MakeXorFrom
assign xor0901 = (xor0856^xor0862^xor0860^xor0858); // MakeXorFrom
assign xor0902 = (xor0864^xor0870^xor0868^xor0866); // MakeXorFrom
assign xor0903 = (xor0884^xor0885^xor0886^xor0883); // MakeXorFrom
assign xor0904 = (xor0889^xor0890^xor0887^xor0888); // MakeXorFrom
assign xor0905 = (xor0894^xor0891^xor0892^xor0893); // MakeXorFrom
assign xor0906 = (xor0897^xor0898^xor0895^xor0896); // MakeXorFrom
assign xor0907 = (xor0899^xor0901^xor0902^xor0900); // MakeXorFrom
assign xor0908 = (xor0905^xor0906^xor0903^xor0904); // MakeXorFrom
assign xor0909 = xor0907;
assign xor0910 = (xor0908^xor0909); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 7
assign xor0911 = (xor0038^xor0036^xor0034^xor0032); // MakeXorFrom
assign xor0912 = (xor0100^xor0098^xor0102^xor0096); // MakeXorFrom
assign xor0913 = (xor0166^xor0164^xor0162^xor0160); // MakeXorFrom
assign xor0914 = (xor0230^xor0228^xor0226^xor0224); // MakeXorFrom
assign xor0915 = (xor0529^xor0532^xor0528^xor0533); // MakeXorFrom
assign xor0916 = (xor0560^xor0565^xor0564^xor0561); // MakeXorFrom
assign xor0917 = (xor0596^xor0593^xor0592^xor0597); // MakeXorFrom
assign xor0918 = (xor0624^xor0629^xor0628^xor0625); // MakeXorFrom
assign xor0919 = (xor0835^xor0834^xor0831^xor0830); // MakeXorFrom
assign xor0920 = (xor0843^xor0839^xor0842^xor0838); // MakeXorFrom
assign xor0921 = (xor0861^xor0862^xor0857^xor0858); // MakeXorFrom
assign xor0922 = (xor0869^xor0870^xor0865^xor0866); // MakeXorFrom
assign xor0923 = (xor0884^xor0890^xor0888^xor0886); // MakeXorFrom
assign xor0924 = (xor0894^xor0892^xor0898^xor0896); // MakeXorFrom
assign xor0925 = (xor0913^xor0914^xor0911^xor0912); // MakeXorFrom
assign xor0926 = (xor0915^xor0916^xor0917^xor0918); // MakeXorFrom
assign xor0927 = (xor0921^xor0922^xor0919^xor0920); // MakeXorFrom
assign xor0928 = (xor0923^xor0924); // MakeXorFrom
assign xor0929 = (xor0926^xor0927^xor0928^xor0925); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 8
assign xor0930 = (xor0066^xor0064^xor0070^xor0068); // MakeXorFrom
assign xor0931 = (xor0194^xor0192^xor0198^xor0196); // MakeXorFrom
assign xor0932 = (xor0548^xor0545^xor0544^xor0549); // MakeXorFrom
assign xor0933 = (xor0613^xor0609^xor0612^xor0608); // MakeXorFrom
assign xor0934 = (xor0851^xor0849^xor0878^xor0876); // MakeXorFrom
assign xor0935 = (xor0889^xor0890^xor0885^xor0886); // MakeXorFrom
assign xor0936 = (xor0894^xor0897^xor0898^xor0893); // MakeXorFrom
assign xor0937 = (xor0916^xor0914^xor0912^xor0918); // MakeXorFrom
assign xor0938 = (xor0933^xor0931^xor0932^xor0930); // MakeXorFrom
assign xor0939 = (xor0936^xor0934^xor0937^xor0935); // MakeXorFrom
assign xor0940 = (xor0939^xor0938); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 9
assign xor0941 = (xor0128^xor0134^xor0132^xor0130); // MakeXorFrom
assign xor0942 = (xor0580^xor0577^xor0576^xor0581); // MakeXorFrom
assign xor0943 = (xor0836^xor0841^xor0837^xor0840); // MakeXorFrom
assign xor0944 = (xor0863^xor0864^xor0867^xor0868); // MakeXorFrom
assign xor0945 = (xor0913^xor0906^xor0914^xor0904); // MakeXorFrom
assign xor0946 = (xor0922^xor0920^xor0917^xor0918); // MakeXorFrom
assign xor0947 = (xor0933^xor0931); // MakeXorFrom
assign xor0948 = (xor0943^xor0944^xor0941^xor0942); // MakeXorFrom
assign xor0949 = (xor0946^xor0947^xor0945); // MakeXorFrom
assign xor0950 = (xor0949^xor0948); // MakeXorFrom
// BuildXorTrees, BuildCheckBit
// BuildCheckBit: building inverse max-parity tree
assign xor0951 = (xor0002^xor0000^xor0006^xor0004); // MakeXorFrom
assign xor0952 = (xor0512^xor0517^xor0516^xor0513); // MakeXorFrom
assign xor0953 = (xor0828^xor0833^xor0832^xor0829); // MakeXorFrom
assign xor0954 = (xor0856^xor0859^xor0860^xor0855); // MakeXorFrom
assign xor0955 = (xor0905^xor0903^xor0911^xor0912); // MakeXorFrom
assign xor0956 = (xor0915^xor0916^xor0921^xor0919); // MakeXorFrom
assign xor0957 = (xor0932^xor0930); // MakeXorFrom
assign xor0958 = (xor0953^xor0954^xor0951^xor0952); // MakeXorFrom
assign xor0959 = (xor0957^xor0955^xor0956); // MakeXorFrom
assign xor0960 = (xor0959^xor0958); // MakeXorFrom
// BuildCheckBit: building check-bit tree
assign xor0961 = (xor0960^xor0950); // MakeXorFrom
assign ecc_parity[-1] = xor0961;
assign ecc_parity[0] = xor0682;
assign ecc_parity[1] = xor0725;
assign ecc_parity[2] = xor0768;
assign ecc_parity[3] = xor0811;
assign ecc_parity[4] = xor0854;
assign ecc_parity[5] = xor0882;
assign ecc_parity[6] = xor0910;
assign ecc_parity[7] = xor0929;
assign ecc_parity[8] = xor0940;
assign ecc_parity[9] = xor0950;
assign input_data[0] = i_chk    [0];
assign input_data[1] = i_chk    [1];
assign input_data[2] = i_chk    [2];
assign input_data[3] = i_data   [0];
assign o_data    [0] = corrected[3];
assign input_data[4] = i_chk    [3];
assign input_data[5] = i_data   [1];
assign o_data    [1] = corrected[5];
assign input_data[6] = i_data   [2];
assign o_data    [2] = corrected[6];
assign input_data[7] = i_data   [3];
assign o_data    [3] = corrected[7];
assign input_data[8] = i_chk    [4];
assign input_data[9] = i_data   [4];
assign o_data    [4] = corrected[9];
assign input_data[10] = i_data   [5];
assign o_data    [5] = corrected[10];
assign input_data[11] = i_data   [6];
assign o_data    [6] = corrected[11];
assign input_data[12] = i_data   [7];
assign o_data    [7] = corrected[12];
assign input_data[13] = i_data   [8];
assign o_data    [8] = corrected[13];
assign input_data[14] = i_data   [9];
assign o_data    [9] = corrected[14];
assign input_data[15] = i_data   [10];
assign o_data    [10] = corrected[15];
assign input_data[16] = i_chk    [5];
assign input_data[17] = i_data   [11];
assign o_data    [11] = corrected[17];
assign input_data[18] = i_data   [12];
assign o_data    [12] = corrected[18];
assign input_data[19] = i_data   [13];
assign o_data    [13] = corrected[19];
assign input_data[20] = i_data   [14];
assign o_data    [14] = corrected[20];
assign input_data[21] = i_data   [15];
assign o_data    [15] = corrected[21];
assign input_data[22] = i_data   [16];
assign o_data    [16] = corrected[22];
assign input_data[23] = i_data   [17];
assign o_data    [17] = corrected[23];
assign input_data[24] = i_data   [18];
assign o_data    [18] = corrected[24];
assign input_data[25] = i_data   [19];
assign o_data    [19] = corrected[25];
assign input_data[26] = i_data   [20];
assign o_data    [20] = corrected[26];
assign input_data[27] = i_data   [21];
assign o_data    [21] = corrected[27];
assign input_data[28] = i_data   [22];
assign o_data    [22] = corrected[28];
assign input_data[29] = i_data   [23];
assign o_data    [23] = corrected[29];
assign input_data[30] = i_data   [24];
assign o_data    [24] = corrected[30];
assign input_data[31] = i_data   [25];
assign o_data    [25] = corrected[31];
assign input_data[32] = i_chk    [6];
assign input_data[33] = i_data   [26];
assign o_data    [26] = corrected[33];
assign input_data[34] = i_data   [27];
assign o_data    [27] = corrected[34];
assign input_data[35] = i_data   [28];
assign o_data    [28] = corrected[35];
assign input_data[36] = i_data   [29];
assign o_data    [29] = corrected[36];
assign input_data[37] = i_data   [30];
assign o_data    [30] = corrected[37];
assign input_data[38] = i_data   [31];
assign o_data    [31] = corrected[38];
assign input_data[39] = i_data   [32];
assign o_data    [32] = corrected[39];
assign input_data[40] = i_data   [33];
assign o_data    [33] = corrected[40];
assign input_data[41] = i_data   [34];
assign o_data    [34] = corrected[41];
assign input_data[42] = i_data   [35];
assign o_data    [35] = corrected[42];
assign input_data[43] = i_data   [36];
assign o_data    [36] = corrected[43];
assign input_data[44] = i_data   [37];
assign o_data    [37] = corrected[44];
assign input_data[45] = i_data   [38];
assign o_data    [38] = corrected[45];
assign input_data[46] = i_data   [39];
assign o_data    [39] = corrected[46];
assign input_data[47] = i_data   [40];
assign o_data    [40] = corrected[47];
assign input_data[48] = i_data   [41];
assign o_data    [41] = corrected[48];
assign input_data[49] = i_data   [42];
assign o_data    [42] = corrected[49];
assign input_data[50] = i_data   [43];
assign o_data    [43] = corrected[50];
assign input_data[51] = i_data   [44];
assign o_data    [44] = corrected[51];
assign input_data[52] = i_data   [45];
assign o_data    [45] = corrected[52];
assign input_data[53] = i_data   [46];
assign o_data    [46] = corrected[53];
assign input_data[54] = i_data   [47];
assign o_data    [47] = corrected[54];
assign input_data[55] = i_data   [48];
assign o_data    [48] = corrected[55];
assign input_data[56] = i_data   [49];
assign o_data    [49] = corrected[56];
assign input_data[57] = i_data   [50];
assign o_data    [50] = corrected[57];
assign input_data[58] = i_data   [51];
assign o_data    [51] = corrected[58];
assign input_data[59] = i_data   [52];
assign o_data    [52] = corrected[59];
assign input_data[60] = i_data   [53];
assign o_data    [53] = corrected[60];
assign input_data[61] = i_data   [54];
assign o_data    [54] = corrected[61];
assign input_data[62] = i_data   [55];
assign o_data    [55] = corrected[62];
assign input_data[63] = i_data   [56];
assign o_data    [56] = corrected[63];
assign input_data[64] = i_chk    [7];
assign input_data[65] = i_data   [57];
assign o_data    [57] = corrected[65];
assign input_data[66] = i_data   [58];
assign o_data    [58] = corrected[66];
assign input_data[67] = i_data   [59];
assign o_data    [59] = corrected[67];
assign input_data[68] = i_data   [60];
assign o_data    [60] = corrected[68];
assign input_data[69] = i_data   [61];
assign o_data    [61] = corrected[69];
assign input_data[70] = i_data   [62];
assign o_data    [62] = corrected[70];
assign input_data[71] = i_data   [63];
assign o_data    [63] = corrected[71];
assign input_data[72] = i_data   [64];
assign o_data    [64] = corrected[72];
assign input_data[73] = i_data   [65];
assign o_data    [65] = corrected[73];
assign input_data[74] = i_data   [66];
assign o_data    [66] = corrected[74];
assign input_data[75] = i_data   [67];
assign o_data    [67] = corrected[75];
assign input_data[76] = i_data   [68];
assign o_data    [68] = corrected[76];
assign input_data[77] = i_data   [69];
assign o_data    [69] = corrected[77];
assign input_data[78] = i_data   [70];
assign o_data    [70] = corrected[78];
assign input_data[79] = i_data   [71];
assign o_data    [71] = corrected[79];
assign input_data[80] = i_data   [72];
assign o_data    [72] = corrected[80];
assign input_data[81] = i_data   [73];
assign o_data    [73] = corrected[81];
assign input_data[82] = i_data   [74];
assign o_data    [74] = corrected[82];
assign input_data[83] = i_data   [75];
assign o_data    [75] = corrected[83];
assign input_data[84] = i_data   [76];
assign o_data    [76] = corrected[84];
assign input_data[85] = i_data   [77];
assign o_data    [77] = corrected[85];
assign input_data[86] = i_data   [78];
assign o_data    [78] = corrected[86];
assign input_data[87] = i_data   [79];
assign o_data    [79] = corrected[87];
assign input_data[88] = i_data   [80];
assign o_data    [80] = corrected[88];
assign input_data[89] = i_data   [81];
assign o_data    [81] = corrected[89];
assign input_data[90] = i_data   [82];
assign o_data    [82] = corrected[90];
assign input_data[91] = i_data   [83];
assign o_data    [83] = corrected[91];
assign input_data[92] = i_data   [84];
assign o_data    [84] = corrected[92];
assign input_data[93] = i_data   [85];
assign o_data    [85] = corrected[93];
assign input_data[94] = i_data   [86];
assign o_data    [86] = corrected[94];
assign input_data[95] = i_data   [87];
assign o_data    [87] = corrected[95];
assign input_data[96] = i_data   [88];
assign o_data    [88] = corrected[96];
assign input_data[97] = i_data   [89];
assign o_data    [89] = corrected[97];
assign input_data[98] = i_data   [90];
assign o_data    [90] = corrected[98];
assign input_data[99] = i_data   [91];
assign o_data    [91] = corrected[99];
assign input_data[100] = i_data   [92];
assign o_data    [92] = corrected[100];
assign input_data[101] = i_data   [93];
assign o_data    [93] = corrected[101];
assign input_data[102] = i_data   [94];
assign o_data    [94] = corrected[102];
assign input_data[103] = i_data   [95];
assign o_data    [95] = corrected[103];
assign input_data[104] = i_data   [96];
assign o_data    [96] = corrected[104];
assign input_data[105] = i_data   [97];
assign o_data    [97] = corrected[105];
assign input_data[106] = i_data   [98];
assign o_data    [98] = corrected[106];
assign input_data[107] = i_data   [99];
assign o_data    [99] = corrected[107];
assign input_data[108] = i_data   [100];
assign o_data    [100] = corrected[108];
assign input_data[109] = i_data   [101];
assign o_data    [101] = corrected[109];
assign input_data[110] = i_data   [102];
assign o_data    [102] = corrected[110];
assign input_data[111] = i_data   [103];
assign o_data    [103] = corrected[111];
assign input_data[112] = i_data   [104];
assign o_data    [104] = corrected[112];
assign input_data[113] = i_data   [105];
assign o_data    [105] = corrected[113];
assign input_data[114] = i_data   [106];
assign o_data    [106] = corrected[114];
assign input_data[115] = i_data   [107];
assign o_data    [107] = corrected[115];
assign input_data[116] = i_data   [108];
assign o_data    [108] = corrected[116];
assign input_data[117] = i_data   [109];
assign o_data    [109] = corrected[117];
assign input_data[118] = i_data   [110];
assign o_data    [110] = corrected[118];
assign input_data[119] = i_data   [111];
assign o_data    [111] = corrected[119];
assign input_data[120] = i_data   [112];
assign o_data    [112] = corrected[120];
assign input_data[121] = i_data   [113];
assign o_data    [113] = corrected[121];
assign input_data[122] = i_data   [114];
assign o_data    [114] = corrected[122];
assign input_data[123] = i_data   [115];
assign o_data    [115] = corrected[123];
assign input_data[124] = i_data   [116];
assign o_data    [116] = corrected[124];
assign input_data[125] = i_data   [117];
assign o_data    [117] = corrected[125];
assign input_data[126] = i_data   [118];
assign o_data    [118] = corrected[126];
assign input_data[127] = i_data   [119];
assign o_data    [119] = corrected[127];
assign input_data[128] = i_chk    [8];
assign input_data[129] = i_data   [120];
assign o_data    [120] = corrected[129];
assign input_data[130] = i_data   [121];
assign o_data    [121] = corrected[130];
assign input_data[131] = i_data   [122];
assign o_data    [122] = corrected[131];
assign input_data[132] = i_data   [123];
assign o_data    [123] = corrected[132];
assign input_data[133] = i_data   [124];
assign o_data    [124] = corrected[133];
assign input_data[134] = i_data   [125];
assign o_data    [125] = corrected[134];
assign input_data[135] = i_data   [126];
assign o_data    [126] = corrected[135];
assign input_data[136] = i_data   [127];
assign o_data    [127] = corrected[136];
assign input_data[137] = i_data   [128];
assign o_data    [128] = corrected[137];
assign input_data[138] = i_data   [129];
assign o_data    [129] = corrected[138];
assign input_data[139] = i_data   [130];
assign o_data    [130] = corrected[139];
assign input_data[140] = i_data   [131];
assign o_data    [131] = corrected[140];
assign input_data[141] = i_data   [132];
assign o_data    [132] = corrected[141];
assign input_data[142] = i_data   [133];
assign o_data    [133] = corrected[142];
assign input_data[143] = i_data   [134];
assign o_data    [134] = corrected[143];
assign input_data[144] = i_data   [135];
assign o_data    [135] = corrected[144];
assign input_data[145] = i_data   [136];
assign o_data    [136] = corrected[145];
assign input_data[146] = i_data   [137];
assign o_data    [137] = corrected[146];
assign input_data[147] = i_data   [138];
assign o_data    [138] = corrected[147];
assign input_data[148] = i_data   [139];
assign o_data    [139] = corrected[148];
assign input_data[149] = i_data   [140];
assign o_data    [140] = corrected[149];
assign input_data[150] = i_data   [141];
assign o_data    [141] = corrected[150];
assign input_data[151] = i_data   [142];
assign o_data    [142] = corrected[151];
assign input_data[152] = i_data   [143];
assign o_data    [143] = corrected[152];
assign input_data[153] = i_data   [144];
assign o_data    [144] = corrected[153];
assign input_data[154] = i_data   [145];
assign o_data    [145] = corrected[154];
assign input_data[155] = i_data   [146];
assign o_data    [146] = corrected[155];
assign input_data[156] = i_data   [147];
assign o_data    [147] = corrected[156];
assign input_data[157] = i_data   [148];
assign o_data    [148] = corrected[157];
assign input_data[158] = i_data   [149];
assign o_data    [149] = corrected[158];
assign input_data[159] = i_data   [150];
assign o_data    [150] = corrected[159];
assign input_data[160] = i_data   [151];
assign o_data    [151] = corrected[160];
assign input_data[161] = i_data   [152];
assign o_data    [152] = corrected[161];
assign input_data[162] = i_data   [153];
assign o_data    [153] = corrected[162];
assign input_data[163] = i_data   [154];
assign o_data    [154] = corrected[163];
assign input_data[164] = i_data   [155];
assign o_data    [155] = corrected[164];
assign input_data[165] = i_data   [156];
assign o_data    [156] = corrected[165];
assign input_data[166] = i_data   [157];
assign o_data    [157] = corrected[166];
assign input_data[167] = i_data   [158];
assign o_data    [158] = corrected[167];
assign input_data[168] = i_data   [159];
assign o_data    [159] = corrected[168];
assign input_data[169] = i_data   [160];
assign o_data    [160] = corrected[169];
assign input_data[170] = i_data   [161];
assign o_data    [161] = corrected[170];
assign input_data[171] = i_data   [162];
assign o_data    [162] = corrected[171];
assign input_data[172] = i_data   [163];
assign o_data    [163] = corrected[172];
assign input_data[173] = i_data   [164];
assign o_data    [164] = corrected[173];
assign input_data[174] = i_data   [165];
assign o_data    [165] = corrected[174];
assign input_data[175] = i_data   [166];
assign o_data    [166] = corrected[175];
assign input_data[176] = i_data   [167];
assign o_data    [167] = corrected[176];
assign input_data[177] = i_data   [168];
assign o_data    [168] = corrected[177];
assign input_data[178] = i_data   [169];
assign o_data    [169] = corrected[178];
assign input_data[179] = i_data   [170];
assign o_data    [170] = corrected[179];
assign input_data[180] = i_data   [171];
assign o_data    [171] = corrected[180];
assign input_data[181] = i_data   [172];
assign o_data    [172] = corrected[181];
assign input_data[182] = i_data   [173];
assign o_data    [173] = corrected[182];
assign input_data[183] = i_data   [174];
assign o_data    [174] = corrected[183];
assign input_data[184] = i_data   [175];
assign o_data    [175] = corrected[184];
assign input_data[185] = i_data   [176];
assign o_data    [176] = corrected[185];
assign input_data[186] = i_data   [177];
assign o_data    [177] = corrected[186];
assign input_data[187] = i_data   [178];
assign o_data    [178] = corrected[187];
assign input_data[188] = i_data   [179];
assign o_data    [179] = corrected[188];
assign input_data[189] = i_data   [180];
assign o_data    [180] = corrected[189];
assign input_data[190] = i_data   [181];
assign o_data    [181] = corrected[190];
assign input_data[191] = i_data   [182];
assign o_data    [182] = corrected[191];
assign input_data[192] = i_data   [183];
assign o_data    [183] = corrected[192];
assign input_data[193] = i_data   [184];
assign o_data    [184] = corrected[193];
assign input_data[194] = i_data   [185];
assign o_data    [185] = corrected[194];
assign input_data[195] = i_data   [186];
assign o_data    [186] = corrected[195];
assign input_data[196] = i_data   [187];
assign o_data    [187] = corrected[196];
assign input_data[197] = i_data   [188];
assign o_data    [188] = corrected[197];
assign input_data[198] = i_data   [189];
assign o_data    [189] = corrected[198];
assign input_data[199] = i_data   [190];
assign o_data    [190] = corrected[199];
assign input_data[200] = i_data   [191];
assign o_data    [191] = corrected[200];
assign input_data[201] = i_data   [192];
assign o_data    [192] = corrected[201];
assign input_data[202] = i_data   [193];
assign o_data    [193] = corrected[202];
assign input_data[203] = i_data   [194];
assign o_data    [194] = corrected[203];
assign input_data[204] = i_data   [195];
assign o_data    [195] = corrected[204];
assign input_data[205] = i_data   [196];
assign o_data    [196] = corrected[205];
assign input_data[206] = i_data   [197];
assign o_data    [197] = corrected[206];
assign input_data[207] = i_data   [198];
assign o_data    [198] = corrected[207];
assign input_data[208] = i_data   [199];
assign o_data    [199] = corrected[208];
assign input_data[209] = i_data   [200];
assign o_data    [200] = corrected[209];
assign input_data[210] = i_data   [201];
assign o_data    [201] = corrected[210];
assign input_data[211] = i_data   [202];
assign o_data    [202] = corrected[211];
assign input_data[212] = i_data   [203];
assign o_data    [203] = corrected[212];
assign input_data[213] = i_data   [204];
assign o_data    [204] = corrected[213];
assign input_data[214] = i_data   [205];
assign o_data    [205] = corrected[214];
assign input_data[215] = i_data   [206];
assign o_data    [206] = corrected[215];
assign input_data[216] = i_data   [207];
assign o_data    [207] = corrected[216];
assign input_data[217] = i_data   [208];
assign o_data    [208] = corrected[217];
assign input_data[218] = i_data   [209];
assign o_data    [209] = corrected[218];
assign input_data[219] = i_data   [210];
assign o_data    [210] = corrected[219];
assign input_data[220] = i_data   [211];
assign o_data    [211] = corrected[220];
assign input_data[221] = i_data   [212];
assign o_data    [212] = corrected[221];
assign input_data[222] = i_data   [213];
assign o_data    [213] = corrected[222];
assign input_data[223] = i_data   [214];
assign o_data    [214] = corrected[223];
assign input_data[224] = i_data   [215];
assign o_data    [215] = corrected[224];
assign input_data[225] = i_data   [216];
assign o_data    [216] = corrected[225];
assign input_data[226] = i_data   [217];
assign o_data    [217] = corrected[226];
assign input_data[227] = i_data   [218];
assign o_data    [218] = corrected[227];
assign input_data[228] = i_data   [219];
assign o_data    [219] = corrected[228];
assign input_data[229] = i_data   [220];
assign o_data    [220] = corrected[229];
assign input_data[230] = i_data   [221];
assign o_data    [221] = corrected[230];
assign input_data[231] = i_data   [222];
assign o_data    [222] = corrected[231];
assign input_data[232] = i_data   [223];
assign o_data    [223] = corrected[232];
assign input_data[233] = i_data   [224];
assign o_data    [224] = corrected[233];
assign input_data[234] = i_data   [225];
assign o_data    [225] = corrected[234];
assign input_data[235] = i_data   [226];
assign o_data    [226] = corrected[235];
assign input_data[236] = i_data   [227];
assign o_data    [227] = corrected[236];
assign input_data[237] = i_data   [228];
assign o_data    [228] = corrected[237];
assign input_data[238] = i_data   [229];
assign o_data    [229] = corrected[238];
assign input_data[239] = i_data   [230];
assign o_data    [230] = corrected[239];
assign input_data[240] = i_data   [231];
assign o_data    [231] = corrected[240];
assign input_data[241] = i_data   [232];
assign o_data    [232] = corrected[241];
assign input_data[242] = i_data   [233];
assign o_data    [233] = corrected[242];
assign input_data[243] = i_data   [234];
assign o_data    [234] = corrected[243];
assign input_data[244] = i_data   [235];
assign o_data    [235] = corrected[244];
assign input_data[245] = i_data   [236];
assign o_data    [236] = corrected[245];
assign input_data[246] = i_data   [237];
assign o_data    [237] = corrected[246];
assign input_data[247] = i_data   [238];
assign o_data    [238] = corrected[247];
assign input_data[248] = i_data   [239];
assign o_data    [239] = corrected[248];
assign input_data[249] = i_data   [240];
assign o_data    [240] = corrected[249];
assign input_data[250] = i_data   [241];
assign o_data    [241] = corrected[250];
assign input_data[251] = i_data   [242];
assign o_data    [242] = corrected[251];
assign input_data[252] = i_data   [243];
assign o_data    [243] = corrected[252];
assign input_data[253] = i_data   [244];
assign o_data    [244] = corrected[253];
assign input_data[254] = i_data   [245];
assign o_data    [245] = corrected[254];
assign input_data[255] = i_data   [246];
assign o_data    [246] = corrected[255];
assign input_data[256] = i_chk    [9];
assign input_data[257] = i_data   [247];
assign o_data    [247] = corrected[257];
assign input_data[258] = i_data   [248];
assign o_data    [248] = corrected[258];
assign input_data[259] = i_data   [249];
assign o_data    [249] = corrected[259];
assign input_data[260] = i_data   [250];
assign o_data    [250] = corrected[260];
assign input_data[261] = i_data   [251];
assign o_data    [251] = corrected[261];
assign input_data[262] = i_data   [252];
assign o_data    [252] = corrected[262];
assign input_data[263] = i_data   [253];
assign o_data    [253] = corrected[263];
assign input_data[264] = i_data   [254];
assign o_data    [254] = corrected[264];
assign input_data[265] = i_data   [255];
assign o_data    [255] = corrected[265];
assign input_data[266] = i_data   [256];
assign o_data    [256] = corrected[266];
assign input_data[267] = i_data   [257];
assign o_data    [257] = corrected[267];
assign input_data[268] = i_data   [258];
assign o_data    [258] = corrected[268];
assign input_data[269] = i_data   [259];
assign o_data    [259] = corrected[269];
assign input_data[270] = i_data   [260];
assign o_data    [260] = corrected[270];
assign input_data[271] = i_data   [261];
assign o_data    [261] = corrected[271];
assign input_data[272] = i_data   [262];
assign o_data    [262] = corrected[272];
assign input_data[273] = i_data   [263];
assign o_data    [263] = corrected[273];
assign input_data[274] = i_data   [264];
assign o_data    [264] = corrected[274];
assign input_data[275] = i_data   [265];
assign o_data    [265] = corrected[275];
assign input_data[276] = i_data   [266];
assign o_data    [266] = corrected[276];
assign input_data[277] = i_data   [267];
assign o_data    [267] = corrected[277];
assign input_data[278] = i_data   [268];
assign o_data    [268] = corrected[278];
assign input_data[279] = i_data   [269];
assign o_data    [269] = corrected[279];
assign input_data[280] = i_data   [270];
assign o_data    [270] = corrected[280];
assign input_data[281] = i_data   [271];
assign o_data    [271] = corrected[281];
assign input_data[282] = i_data   [272];
assign o_data    [272] = corrected[282];
assign input_data[283] = i_data   [273];
assign o_data    [273] = corrected[283];
assign input_data[284] = i_data   [274];
assign o_data    [274] = corrected[284];
assign input_data[285] = i_data   [275];
assign o_data    [275] = corrected[285];
assign input_data[286] = i_data   [276];
assign o_data    [276] = corrected[286];
assign input_data[287] = i_data   [277];
assign o_data    [277] = corrected[287];
assign input_data[288] = i_data   [278];
assign o_data    [278] = corrected[288];
assign input_data[289] = i_data   [279];
assign o_data    [279] = corrected[289];
assign input_data[290] = i_data   [280];
assign o_data    [280] = corrected[290];
assign input_data[291] = i_data   [281];
assign o_data    [281] = corrected[291];
assign input_data[292] = i_data   [282];
assign o_data    [282] = corrected[292];
assign input_data[293] = i_data   [283];
assign o_data    [283] = corrected[293];
assign input_data[294] = i_data   [284];
assign o_data    [284] = corrected[294];
assign input_data[295] = i_data   [285];
assign o_data    [285] = corrected[295];
assign input_data[296] = i_data   [286];
assign o_data    [286] = corrected[296];
assign input_data[297] = i_data   [287];
assign o_data    [287] = corrected[297];
assign input_data[298] = i_data   [288];
assign o_data    [288] = corrected[298];
assign input_data[299] = i_data   [289];
assign o_data    [289] = corrected[299];
assign input_data[300] = i_data   [290];
assign o_data    [290] = corrected[300];
assign input_data[301] = i_data   [291];
assign o_data    [291] = corrected[301];
assign input_data[302] = i_data   [292];
assign o_data    [292] = corrected[302];
assign input_data[303] = i_data   [293];
assign o_data    [293] = corrected[303];
assign input_data[304] = i_data   [294];
assign o_data    [294] = corrected[304];
assign input_data[305] = i_data   [295];
assign o_data    [295] = corrected[305];
assign input_data[306] = i_data   [296];
assign o_data    [296] = corrected[306];
assign input_data[307] = i_data   [297];
assign o_data    [297] = corrected[307];
assign input_data[308] = i_data   [298];
assign o_data    [298] = corrected[308];
assign input_data[309] = i_data   [299];
assign o_data    [299] = corrected[309];
assign input_data[310] = i_data   [300];
assign o_data    [300] = corrected[310];
assign input_data[311] = i_data   [301];
assign o_data    [301] = corrected[311];
assign input_data[312] = i_data   [302];
assign o_data    [302] = corrected[312];
assign input_data[313] = i_data   [303];
assign o_data    [303] = corrected[313];
assign input_data[314] = i_data   [304];
assign o_data    [304] = corrected[314];
assign input_data[315] = i_data   [305];
assign o_data    [305] = corrected[315];
assign input_data[316] = i_data   [306];
assign o_data    [306] = corrected[316];
assign input_data[317] = i_data   [307];
assign o_data    [307] = corrected[317];
assign input_data[318] = i_data   [308];
assign o_data    [308] = corrected[318];
assign input_data[319] = i_data   [309];
assign o_data    [309] = corrected[319];
assign input_data[320] = i_data   [310];
assign o_data    [310] = corrected[320];
assign input_data[321] = i_data   [311];
assign o_data    [311] = corrected[321];
assign input_data[322] = i_data   [312];
assign o_data    [312] = corrected[322];
assign input_data[323] = i_data   [313];
assign o_data    [313] = corrected[323];
assign input_data[324] = i_data   [314];
assign o_data    [314] = corrected[324];
assign input_data[325] = i_data   [315];
assign o_data    [315] = corrected[325];
assign input_data[326] = i_data   [316];
assign o_data    [316] = corrected[326];
assign input_data[327] = i_data   [317];
assign o_data    [317] = corrected[327];
assign input_data[328] = i_data   [318];
assign o_data    [318] = corrected[328];
assign input_data[329] = i_data   [319];
assign o_data    [319] = corrected[329];
assign input_data[330] = i_data   [320];
assign o_data    [320] = corrected[330];
assign input_data[331] = i_data   [321];
assign o_data    [321] = corrected[331];
assign input_data[332] = i_data   [322];
assign o_data    [322] = corrected[332];
assign input_data[333] = i_data   [323];
assign o_data    [323] = corrected[333];
assign input_data[334] = i_data   [324];
assign o_data    [324] = corrected[334];
assign input_data[335] = i_data   [325];
assign o_data    [325] = corrected[335];
assign input_data[336] = i_data   [326];
assign o_data    [326] = corrected[336];
assign input_data[337] = i_data   [327];
assign o_data    [327] = corrected[337];
assign input_data[338] = i_data   [328];
assign o_data    [328] = corrected[338];
assign input_data[339] = i_data   [329];
assign o_data    [329] = corrected[339];
assign input_data[340] = i_data   [330];
assign o_data    [330] = corrected[340];
assign input_data[341] = i_data   [331];
assign o_data    [331] = corrected[341];
assign input_data[342] = i_data   [332];
assign o_data    [332] = corrected[342];
assign input_data[343] = i_data   [333];
assign o_data    [333] = corrected[343];
assign input_data[344] = i_data   [334];
assign o_data    [334] = corrected[344];
assign input_data[345] = i_data   [335];
assign o_data    [335] = corrected[345];
assign input_data[346] = i_data   [336];
assign o_data    [336] = corrected[346];
assign input_data[347] = i_data   [337];
assign o_data    [337] = corrected[347];
assign input_data[348] = i_data   [338];
assign o_data    [338] = corrected[348];
assign input_data[349] = i_data   [339];
assign o_data    [339] = corrected[349];
assign input_data[350] = i_data   [340];
assign o_data    [340] = corrected[350];
assign input_data[351] = i_data   [341];
assign o_data    [341] = corrected[351];
assign input_data[352] = i_data   [342];
assign o_data    [342] = corrected[352];
assign input_data[353] = i_data   [343];
assign o_data    [343] = corrected[353];
assign input_data[354] = i_data   [344];
assign o_data    [344] = corrected[354];
assign input_data[355] = i_data   [345];
assign o_data    [345] = corrected[355];
assign input_data[356] = i_data   [346];
assign o_data    [346] = corrected[356];
assign input_data[357] = i_data   [347];
assign o_data    [347] = corrected[357];
assign input_data[358] = i_data   [348];
assign o_data    [348] = corrected[358];
assign input_data[359] = i_data   [349];
assign o_data    [349] = corrected[359];
assign input_data[360] = i_data   [350];
assign o_data    [350] = corrected[360];
assign input_data[361] = i_data   [351];
assign o_data    [351] = corrected[361];
assign input_data[362] = i_data   [352];
assign o_data    [352] = corrected[362];
assign input_data[363] = i_data   [353];
assign o_data    [353] = corrected[363];
assign input_data[364] = i_data   [354];
assign o_data    [354] = corrected[364];
assign input_data[365] = i_data   [355];
assign o_data    [355] = corrected[365];
assign input_data[366] = i_data   [356];
assign o_data    [356] = corrected[366];
assign input_data[367] = i_data   [357];
assign o_data    [357] = corrected[367];
assign input_data[368] = i_data   [358];
assign o_data    [358] = corrected[368];
assign input_data[369] = i_data   [359];
assign o_data    [359] = corrected[369];
assign input_data[370] = i_data   [360];
assign o_data    [360] = corrected[370];
assign input_data[371] = i_data   [361];
assign o_data    [361] = corrected[371];
assign input_data[372] = i_data   [362];
assign o_data    [362] = corrected[372];
assign input_data[373] = i_data   [363];
assign o_data    [363] = corrected[373];
assign input_data[374] = i_data   [364];
assign o_data    [364] = corrected[374];
assign input_data[375] = i_data   [365];
assign o_data    [365] = corrected[375];
assign input_data[376] = i_data   [366];
assign o_data    [366] = corrected[376];
assign input_data[377] = i_data   [367];
assign o_data    [367] = corrected[377];
assign input_data[378] = i_data   [368];
assign o_data    [368] = corrected[378];
assign input_data[379] = i_data   [369];
assign o_data    [369] = corrected[379];
assign input_data[380] = i_data   [370];
assign o_data    [370] = corrected[380];
assign input_data[381] = i_data   [371];
assign o_data    [371] = corrected[381];
assign input_data[382] = i_data   [372];
assign o_data    [372] = corrected[382];
assign input_data[383] = i_data   [373];
assign o_data    [373] = corrected[383];
assign input_data[384] = i_data   [374];
assign o_data    [374] = corrected[384];
assign input_data[385] = i_data   [375];
assign o_data    [375] = corrected[385];
assign input_data[386] = i_data   [376];
assign o_data    [376] = corrected[386];
assign input_data[387] = i_data   [377];
assign o_data    [377] = corrected[387];
assign input_data[388] = i_data   [378];
assign o_data    [378] = corrected[388];
assign input_data[389] = i_data   [379];
assign o_data    [379] = corrected[389];
assign input_data[390] = i_data   [380];
assign o_data    [380] = corrected[390];
assign input_data[391] = i_data   [381];
assign o_data    [381] = corrected[391];
assign input_data[392] = i_data   [382];
assign o_data    [382] = corrected[392];
assign input_data[393] = i_data   [383];
assign o_data    [383] = corrected[393];
assign input_data[394] = i_data   [384];
assign o_data    [384] = corrected[394];
assign input_data[395] = i_data   [385];
assign o_data    [385] = corrected[395];
assign input_data[396] = i_data   [386];
assign o_data    [386] = corrected[396];
assign input_data[397] = i_data   [387];
assign o_data    [387] = corrected[397];
assign input_data[398] = i_data   [388];
assign o_data    [388] = corrected[398];
assign input_data[399] = i_data   [389];
assign o_data    [389] = corrected[399];
assign input_data[400] = i_data   [390];
assign o_data    [390] = corrected[400];
assign input_data[401] = i_data   [391];
assign o_data    [391] = corrected[401];
assign input_data[402] = i_data   [392];
assign o_data    [392] = corrected[402];
assign input_data[403] = i_data   [393];
assign o_data    [393] = corrected[403];
assign input_data[404] = i_data   [394];
assign o_data    [394] = corrected[404];
assign input_data[405] = i_data   [395];
assign o_data    [395] = corrected[405];
assign input_data[406] = i_data   [396];
assign o_data    [396] = corrected[406];
assign input_data[407] = i_data   [397];
assign o_data    [397] = corrected[407];
assign input_data[408] = i_data   [398];
assign o_data    [398] = corrected[408];
assign input_data[409] = i_data   [399];
assign o_data    [399] = corrected[409];
assign input_data[410] = i_data   [400];
assign o_data    [400] = corrected[410];
assign input_data[411] = i_data   [401];
assign o_data    [401] = corrected[411];
assign input_data[412] = i_data   [402];
assign o_data    [402] = corrected[412];
assign input_data[413] = i_data   [403];
assign o_data    [403] = corrected[413];
assign input_data[414] = i_data   [404];
assign o_data    [404] = corrected[414];
assign input_data[415] = i_data   [405];
assign o_data    [405] = corrected[415];
assign input_data[416] = i_data   [406];
assign o_data    [406] = corrected[416];
assign input_data[417] = i_data   [407];
assign o_data    [407] = corrected[417];
assign input_data[418] = i_data   [408];
assign o_data    [408] = corrected[418];
assign input_data[419] = i_data   [409];
assign o_data    [409] = corrected[419];
assign input_data[420] = i_data   [410];
assign o_data    [410] = corrected[420];
assign input_data[421] = i_data   [411];
assign o_data    [411] = corrected[421];
assign input_data[422] = i_data   [412];
assign o_data    [412] = corrected[422];
assign input_data[423] = i_data   [413];
assign o_data    [413] = corrected[423];
assign input_data[424] = i_data   [414];
assign o_data    [414] = corrected[424];
assign input_data[425] = i_data   [415];
assign o_data    [415] = corrected[425];
assign input_data[426] = i_data   [416];
assign o_data    [416] = corrected[426];
assign input_data[427] = i_data   [417];
assign o_data    [417] = corrected[427];
assign input_data[428] = i_data   [418];
assign o_data    [418] = corrected[428];
assign input_data[429] = i_data   [419];
assign o_data    [419] = corrected[429];
assign input_data[430] = i_data   [420];
assign o_data    [420] = corrected[430];
assign input_data[431] = i_data   [421];
assign o_data    [421] = corrected[431];
assign input_data[432] = i_data   [422];
assign o_data    [422] = corrected[432];
assign input_data[433] = i_data   [423];
assign o_data    [423] = corrected[433];
assign input_data[434] = i_data   [424];
assign o_data    [424] = corrected[434];
assign input_data[435] = i_data   [425];
assign o_data    [425] = corrected[435];
assign input_data[436] = i_data   [426];
assign o_data    [426] = corrected[436];
assign input_data[437] = i_data   [427];
assign o_data    [427] = corrected[437];
assign input_data[438] = i_data   [428];
assign o_data    [428] = corrected[438];
assign input_data[439] = i_data   [429];
assign o_data    [429] = corrected[439];
assign input_data[440] = i_data   [430];
assign o_data    [430] = corrected[440];
assign input_data[441] = i_data   [431];
assign o_data    [431] = corrected[441];
assign input_data[442] = i_data   [432];
assign o_data    [432] = corrected[442];
assign input_data[443] = i_data   [433];
assign o_data    [433] = corrected[443];
assign input_data[444] = i_data   [434];
assign o_data    [434] = corrected[444];
assign input_data[445] = i_data   [435];
assign o_data    [435] = corrected[445];
assign input_data[446] = i_data   [436];
assign o_data    [436] = corrected[446];
assign input_data[447] = i_data   [437];
assign o_data    [437] = corrected[447];
assign input_data[448] = i_data   [438];
assign o_data    [438] = corrected[448];
assign input_data[449] = i_data   [439];
assign o_data    [439] = corrected[449];
assign input_data[450] = i_data   [440];
assign o_data    [440] = corrected[450];
assign input_data[451] = i_data   [441];
assign o_data    [441] = corrected[451];
assign input_data[452] = i_data   [442];
assign o_data    [442] = corrected[452];
assign input_data[453] = i_data   [443];
assign o_data    [443] = corrected[453];
assign input_data[454] = i_data   [444];
assign o_data    [444] = corrected[454];
assign input_data[455] = i_data   [445];
assign o_data    [445] = corrected[455];
assign input_data[456] = i_data   [446];
assign o_data    [446] = corrected[456];
assign input_data[457] = i_data   [447];
assign o_data    [447] = corrected[457];
assign input_data[458] = i_data   [448];
assign o_data    [448] = corrected[458];
assign input_data[459] = i_data   [449];
assign o_data    [449] = corrected[459];
assign input_data[460] = i_data   [450];
assign o_data    [450] = corrected[460];
assign input_data[461] = i_data   [451];
assign o_data    [451] = corrected[461];
assign input_data[462] = i_data   [452];
assign o_data    [452] = corrected[462];
assign input_data[463] = i_data   [453];
assign o_data    [453] = corrected[463];
assign input_data[464] = i_data   [454];
assign o_data    [454] = corrected[464];
assign input_data[465] = i_data   [455];
assign o_data    [455] = corrected[465];
assign input_data[466] = i_data   [456];
assign o_data    [456] = corrected[466];
assign input_data[467] = i_data   [457];
assign o_data    [457] = corrected[467];
assign input_data[468] = i_data   [458];
assign o_data    [458] = corrected[468];
assign input_data[469] = i_data   [459];
assign o_data    [459] = corrected[469];
assign input_data[470] = i_data   [460];
assign o_data    [460] = corrected[470];
assign input_data[471] = i_data   [461];
assign o_data    [461] = corrected[471];
assign input_data[472] = i_data   [462];
assign o_data    [462] = corrected[472];
assign input_data[473] = i_data   [463];
assign o_data    [463] = corrected[473];
assign input_data[474] = i_data   [464];
assign o_data    [464] = corrected[474];
assign input_data[475] = i_data   [465];
assign o_data    [465] = corrected[475];
assign input_data[476] = i_data   [466];
assign o_data    [466] = corrected[476];
assign input_data[477] = i_data   [467];
assign o_data    [467] = corrected[477];
assign input_data[478] = i_data   [468];
assign o_data    [468] = corrected[478];
assign input_data[479] = i_data   [469];
assign o_data    [469] = corrected[479];
assign input_data[480] = i_data   [470];
assign o_data    [470] = corrected[480];
assign input_data[481] = i_data   [471];
assign o_data    [471] = corrected[481];
assign input_data[482] = i_data   [472];
assign o_data    [472] = corrected[482];
assign input_data[483] = i_data   [473];
assign o_data    [473] = corrected[483];
assign input_data[484] = i_data   [474];
assign o_data    [474] = corrected[484];
assign input_data[485] = i_data   [475];
assign o_data    [475] = corrected[485];
assign input_data[486] = i_data   [476];
assign o_data    [476] = corrected[486];
assign input_data[487] = i_data   [477];
assign o_data    [477] = corrected[487];
assign input_data[488] = i_data   [478];
assign o_data    [478] = corrected[488];
assign input_data[489] = i_data   [479];
assign o_data    [479] = corrected[489];
assign input_data[490] = i_data   [480];
assign o_data    [480] = corrected[490];
assign input_data[491] = i_data   [481];
assign o_data    [481] = corrected[491];
assign input_data[492] = i_data   [482];
assign o_data    [482] = corrected[492];
assign input_data[493] = i_data   [483];
assign o_data    [483] = corrected[493];
assign input_data[494] = i_data   [484];
assign o_data    [484] = corrected[494];
assign input_data[495] = i_data   [485];
assign o_data    [485] = corrected[495];
assign input_data[496] = i_data   [486];
assign o_data    [486] = corrected[496];
assign input_data[497] = i_data   [487];
assign o_data    [487] = corrected[497];
assign input_data[498] = i_data   [488];
assign o_data    [488] = corrected[498];
assign input_data[499] = i_data   [489];
assign o_data    [489] = corrected[499];
assign input_data[500] = i_data   [490];
assign o_data    [490] = corrected[500];
assign input_data[501] = i_data   [491];
assign o_data    [491] = corrected[501];
assign input_data[502] = i_data   [492];
assign o_data    [492] = corrected[502];
assign input_data[503] = i_data   [493];
assign o_data    [493] = corrected[503];
assign input_data[504] = i_data   [494];
assign o_data    [494] = corrected[504];
assign input_data[505] = i_data   [495];
assign o_data    [495] = corrected[505];
assign input_data[506] = i_data   [496];
assign o_data    [496] = corrected[506];
assign input_data[507] = i_data   [497];
assign o_data    [497] = corrected[507];
assign input_data[508] = i_data   [498];
assign o_data    [498] = corrected[508];
assign input_data[509] = i_data   [499];
assign o_data    [499] = corrected[509];
assign input_data[510] = i_data   [500];
assign o_data    [500] = corrected[510];
assign input_data[511] = i_data   [501];
assign o_data    [501] = corrected[511];
assign input_data[512] = i_chk    [10];
assign input_data[513] = i_data   [502];
assign o_data    [502] = corrected[513];
assign input_data[514] = i_data   [503];
assign o_data    [503] = corrected[514];
assign input_data[515] = i_data   [504];
assign o_data    [504] = corrected[515];
assign input_data[516] = i_data   [505];
assign o_data    [505] = corrected[516];
assign input_data[517] = i_data   [506];
assign o_data    [506] = corrected[517];
assign input_data[518] = i_data   [507];
assign o_data    [507] = corrected[518];
assign input_data[519] = i_data   [508];
assign o_data    [508] = corrected[519];
assign input_data[520] = i_data   [509];
assign o_data    [509] = corrected[520];
assign input_data[521] = i_data   [510];
assign o_data    [510] = corrected[521];
assign input_data[522] = i_data   [511];
assign o_data    [511] = corrected[522];
assign input_data[523] = i_data   [512];
assign o_data    [512] = corrected[523];
assign input_data[524] = i_data   [513];
assign o_data    [513] = corrected[524];
assign input_data[525] = i_data   [514];
assign o_data    [514] = corrected[525];
assign input_data[526] = i_data   [515];
assign o_data    [515] = corrected[526];
assign input_data[527] = i_data   [516];
assign o_data    [516] = corrected[527];
assign input_data[528] = i_data   [517];
assign o_data    [517] = corrected[528];
assign input_data[529] = i_data   [518];
assign o_data    [518] = corrected[529];
assign input_data[530] = i_data   [519];
assign o_data    [519] = corrected[530];
assign input_data[531] = i_data   [520];
assign o_data    [520] = corrected[531];
assign input_data[532] = i_data   [521];
assign o_data    [521] = corrected[532];
assign input_data[533] = i_data   [522];
assign o_data    [522] = corrected[533];
assign input_data[534] = i_data   [523];
assign o_data    [523] = corrected[534];
assign input_data[535] = i_data   [524];
assign o_data    [524] = corrected[535];
assign input_data[536] = i_data   [525];
assign o_data    [525] = corrected[536];
assign input_data[537] = i_data   [526];
assign o_data    [526] = corrected[537];
assign input_data[538] = i_data   [527];
assign o_data    [527] = corrected[538];
assign input_data[539] = i_data   [528];
assign o_data    [528] = corrected[539];
assign input_data[540] = i_data   [529];
assign o_data    [529] = corrected[540];
assign input_data[541] = i_data   [530];
assign o_data    [530] = corrected[541];
assign input_data[542] = i_data   [531];
assign o_data    [531] = corrected[542];
assign input_data[543] = i_data   [532];
assign o_data    [532] = corrected[543];
assign input_data[544] = i_data   [533];
assign o_data    [533] = corrected[544];
assign input_data[545] = i_data   [534];
assign o_data    [534] = corrected[545];
assign input_data[546] = i_data   [535];
assign o_data    [535] = corrected[546];
assign input_data[547] = i_data   [536];
assign o_data    [536] = corrected[547];
assign input_data[548] = i_data   [537];
assign o_data    [537] = corrected[548];
assign input_data[549] = i_data   [538];
assign o_data    [538] = corrected[549];
assign input_data[550] = i_data   [539];
assign o_data    [539] = corrected[550];
assign input_data[551] = i_data   [540];
assign o_data    [540] = corrected[551];
assign input_data[552] = i_data   [541];
assign o_data    [541] = corrected[552];
assign input_data[553] = i_data   [542];
assign o_data    [542] = corrected[553];
assign input_data[554] = i_data   [543];
assign o_data    [543] = corrected[554];
assign input_data[555] = i_data   [544];
assign o_data    [544] = corrected[555];
assign input_data[556] = i_data   [545];
assign o_data    [545] = corrected[556];
assign input_data[557] = i_data   [546];
assign o_data    [546] = corrected[557];
assign input_data[558] = i_data   [547];
assign o_data    [547] = corrected[558];
assign input_data[559] = i_data   [548];
assign o_data    [548] = corrected[559];
assign input_data[560] = i_data   [549];
assign o_data    [549] = corrected[560];
assign input_data[561] = i_data   [550];
assign o_data    [550] = corrected[561];
assign input_data[562] = i_data   [551];
assign o_data    [551] = corrected[562];
assign input_data[563] = i_data   [552];
assign o_data    [552] = corrected[563];
assign input_data[564] = i_data   [553];
assign o_data    [553] = corrected[564];
assign input_data[565] = i_data   [554];
assign o_data    [554] = corrected[565];
assign input_data[566] = i_data   [555];
assign o_data    [555] = corrected[566];
assign input_data[567] = i_data   [556];
assign o_data    [556] = corrected[567];
assign input_data[568] = i_data   [557];
assign o_data    [557] = corrected[568];
assign input_data[569] = i_data   [558];
assign o_data    [558] = corrected[569];
assign input_data[570] = i_data   [559];
assign o_data    [559] = corrected[570];
assign input_data[571] = i_data   [560];
assign o_data    [560] = corrected[571];
assign input_data[572] = i_data   [561];
assign o_data    [561] = corrected[572];
assign input_data[573] = i_data   [562];
assign o_data    [562] = corrected[573];
assign input_data[574] = i_data   [563];
assign o_data    [563] = corrected[574];
assign input_data[575] = i_data   [564];
assign o_data    [564] = corrected[575];
assign input_data[576] = i_data   [565];
assign o_data    [565] = corrected[576];
assign input_data[577] = i_data   [566];
assign o_data    [566] = corrected[577];
assign input_data[578] = i_data   [567];
assign o_data    [567] = corrected[578];
assign input_data[579] = i_data   [568];
assign o_data    [568] = corrected[579];
assign input_data[580] = i_data   [569];
assign o_data    [569] = corrected[580];
assign input_data[581] = i_data   [570];
assign o_data    [570] = corrected[581];
assign input_data[582] = i_data   [571];
assign o_data    [571] = corrected[582];
assign input_data[583] = i_data   [572];
assign o_data    [572] = corrected[583];
assign input_data[584] = i_data   [573];
assign o_data    [573] = corrected[584];
assign input_data[585] = i_data   [574];
assign o_data    [574] = corrected[585];
assign input_data[586] = i_data   [575];
assign o_data    [575] = corrected[586];
assign input_data[587] = i_data   [576];
assign o_data    [576] = corrected[587];
assign input_data[588] = i_data   [577];
assign o_data    [577] = corrected[588];
assign input_data[589] = i_data   [578];
assign o_data    [578] = corrected[589];
assign input_data[590] = i_data   [579];
assign o_data    [579] = corrected[590];
assign input_data[591] = i_data   [580];
assign o_data    [580] = corrected[591];
assign input_data[592] = i_data   [581];
assign o_data    [581] = corrected[592];
assign input_data[593] = i_data   [582];
assign o_data    [582] = corrected[593];
assign input_data[594] = i_data   [583];
assign o_data    [583] = corrected[594];
assign input_data[595] = i_data   [584];
assign o_data    [584] = corrected[595];
assign input_data[596] = i_data   [585];
assign o_data    [585] = corrected[596];
assign input_data[597] = i_data   [586];
assign o_data    [586] = corrected[597];
assign input_data[598] = i_data   [587];
assign o_data    [587] = corrected[598];
assign input_data[599] = i_data   [588];
assign o_data    [588] = corrected[599];
assign input_data[600] = i_data   [589];
assign o_data    [589] = corrected[600];
assign input_data[601] = i_data   [590];
assign o_data    [590] = corrected[601];
assign input_data[602] = i_data   [591];
assign o_data    [591] = corrected[602];
assign input_data[603] = i_data   [592];
assign o_data    [592] = corrected[603];
assign input_data[604] = i_data   [593];
assign o_data    [593] = corrected[604];
assign input_data[605] = i_data   [594];
assign o_data    [594] = corrected[605];
assign input_data[606] = i_data   [595];
assign o_data    [595] = corrected[606];
assign input_data[607] = i_data   [596];
assign o_data    [596] = corrected[607];
assign input_data[608] = i_data   [597];
assign o_data    [597] = corrected[608];
assign input_data[609] = i_data   [598];
assign o_data    [598] = corrected[609];
assign input_data[610] = i_data   [599];
assign o_data    [599] = corrected[610];
assign input_data[611] = i_data   [600];
assign o_data    [600] = corrected[611];
assign input_data[612] = i_data   [601];
assign o_data    [601] = corrected[612];
assign input_data[613] = i_data   [602];
assign o_data    [602] = corrected[613];
assign input_data[614] = i_data   [603];
assign o_data    [603] = corrected[614];
assign input_data[615] = i_data   [604];
assign o_data    [604] = corrected[615];
assign input_data[616] = i_data   [605];
assign o_data    [605] = corrected[616];
assign input_data[617] = i_data   [606];
assign o_data    [606] = corrected[617];
assign input_data[618] = i_data   [607];
assign o_data    [607] = corrected[618];
assign input_data[619] = i_data   [608];
assign o_data    [608] = corrected[619];
assign input_data[620] = i_data   [609];
assign o_data    [609] = corrected[620];
assign input_data[621] = i_data   [610];
assign o_data    [610] = corrected[621];
assign input_data[622] = i_data   [611];
assign o_data    [611] = corrected[622];
assign input_data[623] = i_data   [612];
assign o_data    [612] = corrected[623];
assign input_data[624] = i_data   [613];
assign o_data    [613] = corrected[624];
assign input_data[625] = i_data   [614];
assign o_data    [614] = corrected[625];
assign input_data[626] = i_data   [615];
assign o_data    [615] = corrected[626];
assign input_data[627] = i_data   [616];
assign o_data    [616] = corrected[627];
assign input_data[628] = i_data   [617];
assign o_data    [617] = corrected[628];
assign input_data[629] = i_data   [618];
assign o_data    [618] = corrected[629];
assign input_data[630] = i_data   [619];
assign o_data    [619] = corrected[630];
assign input_data[631] = i_data   [620];
assign o_data    [620] = corrected[631];
assign input_data[632] = i_data   [621];
assign o_data    [621] = corrected[632];
assign input_data[633] = i_data   [622];
assign o_data    [622] = corrected[633];
assign input_data[634] = i_data   [623];
assign o_data    [623] = corrected[634];
assign input_data[635] = i_data   [624];
assign o_data    [624] = corrected[635];
assign input_data[636] = i_data   [625];
assign o_data    [625] = corrected[636];
assign input_data[637] = i_data   [626];
assign o_data    [626] = corrected[637];
assign input_data[638] = i_data   [627];
assign o_data    [627] = corrected[638];
assign input_data[639] = i_data   [628];
assign o_data    [628] = corrected[639];
assign input_data[640] = i_data   [629];
assign o_data    [629] = corrected[640];
assign input_data[641] = i_data   [630];
assign o_data    [630] = corrected[641];
assign input_data[642] = i_data   [631];
assign o_data    [631] = corrected[642];
assign input_data[643] = i_data   [632];
assign o_data    [632] = corrected[643];
assign input_data[644] = i_data   [633];
assign o_data    [633] = corrected[644];
assign input_data[645] = i_data   [634];
assign o_data    [634] = corrected[645];
assign input_data[646] = i_data   [635];
assign o_data    [635] = corrected[646];
assign input_data[647] = i_data   [636];
assign o_data    [636] = corrected[647];
assign input_data[648] = i_data   [637];
assign o_data    [637] = corrected[648];
assign input_data[649] = i_data   [638];
assign o_data    [638] = corrected[649];
assign input_data[650] = i_data   [639];
assign o_data    [639] = corrected[650];
assign input_data[651] = i_data   [640];
assign o_data    [640] = corrected[651];
assign input_data[652] = i_data   [641];
assign o_data    [641] = corrected[652];
assign input_data[653] = i_data   [642];
assign o_data    [642] = corrected[653];
assign input_data[654] = i_data   [643];
assign o_data    [643] = corrected[654];
assign input_data[655] = i_data   [644];
assign o_data    [644] = corrected[655];
assign input_data[656] = i_data   [645];
assign o_data    [645] = corrected[656];
assign input_data[657] = i_data   [646];
assign o_data    [646] = corrected[657];
assign input_data[658] = i_data   [647];
assign o_data    [647] = corrected[658];
assign input_data[659] = i_data   [648];
assign o_data    [648] = corrected[659];
assign input_data[660] = i_data   [649];
assign o_data    [649] = corrected[660];
assign input_data[661] = i_data   [650];
assign o_data    [650] = corrected[661];
assign input_data[662] = i_data   [651];
assign o_data    [651] = corrected[662];
assign input_data[663] = i_data   [652];
assign o_data    [652] = corrected[663];
assign input_data[664] = i_data   [653];
assign o_data    [653] = corrected[664];
assign input_data[665] = i_data   [654];
assign o_data    [654] = corrected[665];
assign input_data[666] = i_data   [655];
assign o_data    [655] = corrected[666];
assign input_data[667] = i_data   [656];
assign o_data    [656] = corrected[667];
assign input_data[668] = i_data   [657];
assign o_data    [657] = corrected[668];
assign input_data[669] = i_data   [658];
assign o_data    [658] = corrected[669];
assign input_data[670] = i_data   [659];
assign o_data    [659] = corrected[670];
assign input_data[671] = i_data   [660];
assign o_data    [660] = corrected[671];
assign input_data[672] = i_data   [661];
assign o_data    [661] = corrected[672];
assign input_data[673] = i_data   [662];
assign o_data    [662] = corrected[673];
assign input_data[674] = i_data   [663];
assign o_data    [663] = corrected[674];
assign input_data[675] = i_data   [664];
assign o_data    [664] = corrected[675];
assign input_data[676] = i_data   [665];
assign o_data    [665] = corrected[676];
assign input_data[677] = i_data   [666];
assign o_data    [666] = corrected[677];
assign input_data[678] = i_data   [667];
assign o_data    [667] = corrected[678];
assign input_data[679] = i_data   [668];
assign o_data    [668] = corrected[679];
assign input_data[680] = i_data   [669];
assign o_data    [669] = corrected[680];
assign input_data[681] = i_data   [670];
assign o_data    [670] = corrected[681];
assign input_data[682] = i_data   [671];
assign o_data    [671] = corrected[682];
assign input_data[683] = i_data   [672];
assign o_data    [672] = corrected[683];
assign input_data[684] = i_data   [673];
assign o_data    [673] = corrected[684];
assign input_data[685] = i_data   [674];
assign o_data    [674] = corrected[685];
assign input_data[686] = i_data   [675];
assign o_data    [675] = corrected[686];
assign input_data[687] = i_data   [676];
assign o_data    [676] = corrected[687];
assign input_data[688] = i_data   [677];
assign o_data    [677] = corrected[688];
assign input_data[689] = i_data   [678];
assign o_data    [678] = corrected[689];
assign input_data[690] = i_data   [679];
assign o_data    [679] = corrected[690];
assign input_data[691] = i_data   [680];
assign o_data    [680] = corrected[691];
assign input_data[692] = i_data   [681];
assign o_data    [681] = corrected[692];
assign input_data[693] = i_data   [682];
assign o_data    [682] = corrected[693];
assign input_data[694] = i_data   [683];
assign o_data    [683] = corrected[694];
assign input_data[695] = i_data   [684];
assign o_data    [684] = corrected[695];
assign input_data[696] = i_data   [685];
assign o_data    [685] = corrected[696];
assign input_data[697] = i_data   [686];
assign o_data    [686] = corrected[697];
assign input_data[698] = i_data   [687];
assign o_data    [687] = corrected[698];
assign input_data[699] = i_data   [688];
assign o_data    [688] = corrected[699];
assign input_data[700] = i_data   [689];
assign o_data    [689] = corrected[700];
assign input_data[701] = i_data   [690];
assign o_data    [690] = corrected[701];
assign input_data[702] = i_data   [691];
assign o_data    [691] = corrected[702];
assign input_data[703] = i_data   [692];
assign o_data    [692] = corrected[703];
assign input_data[704] = i_data   [693];
assign o_data    [693] = corrected[704];
assign input_data[705] = i_data   [694];
assign o_data    [694] = corrected[705];
assign input_data[706] = i_data   [695];
assign o_data    [695] = corrected[706];
assign input_data[707] = i_data   [696];
assign o_data    [696] = corrected[707];
assign input_data[708] = i_data   [697];
assign o_data    [697] = corrected[708];
assign input_data[709] = i_data   [698];
assign o_data    [698] = corrected[709];
assign input_data[710] = i_data   [699];
assign o_data    [699] = corrected[710];
assign input_data[711] = i_data   [700];
assign o_data    [700] = corrected[711];
assign input_data[712] = i_data   [701];
assign o_data    [701] = corrected[712];
assign input_data[713] = i_data   [702];
assign o_data    [702] = corrected[713];
assign input_data[714] = i_data   [703];
assign o_data    [703] = corrected[714];
assign input_data[715] = i_data   [704];
assign o_data    [704] = corrected[715];
assign input_data[716] = i_data   [705];
assign o_data    [705] = corrected[716];
assign input_data[717] = i_data   [706];
assign o_data    [706] = corrected[717];
assign input_data[718] = i_data   [707];
assign o_data    [707] = corrected[718];
assign input_data[719] = i_data   [708];
assign o_data    [708] = corrected[719];
assign input_data[720] = i_data   [709];
assign o_data    [709] = corrected[720];
assign input_data[721] = i_data   [710];
assign o_data    [710] = corrected[721];
assign input_data[722] = i_data   [711];
assign o_data    [711] = corrected[722];
assign input_data[723] = i_data   [712];
assign o_data    [712] = corrected[723];
assign input_data[724] = i_data   [713];
assign o_data    [713] = corrected[724];
assign input_data[725] = i_data   [714];
assign o_data    [714] = corrected[725];
assign input_data[726] = i_data   [715];
assign o_data    [715] = corrected[726];
assign input_data[727] = i_data   [716];
assign o_data    [716] = corrected[727];
assign input_data[728] = i_data   [717];
assign o_data    [717] = corrected[728];
assign input_data[729] = i_data   [718];
assign o_data    [718] = corrected[729];
assign input_data[730] = i_data   [719];
assign o_data    [719] = corrected[730];
assign input_data[731] = i_data   [720];
assign o_data    [720] = corrected[731];
assign input_data[732] = i_data   [721];
assign o_data    [721] = corrected[732];
assign input_data[733] = i_data   [722];
assign o_data    [722] = corrected[733];
assign input_data[734] = i_data   [723];
assign o_data    [723] = corrected[734];
assign input_data[735] = i_data   [724];
assign o_data    [724] = corrected[735];
assign input_data[736] = i_data   [725];
assign o_data    [725] = corrected[736];
assign input_data[737] = i_data   [726];
assign o_data    [726] = corrected[737];
assign input_data[738] = i_data   [727];
assign o_data    [727] = corrected[738];
assign input_data[739] = i_data   [728];
assign o_data    [728] = corrected[739];
assign input_data[740] = i_data   [729];
assign o_data    [729] = corrected[740];
assign input_data[741] = i_data   [730];
assign o_data    [730] = corrected[741];
assign input_data[742] = i_data   [731];
assign o_data    [731] = corrected[742];
assign input_data[743] = i_data   [732];
assign o_data    [732] = corrected[743];
assign input_data[744] = i_data   [733];
assign o_data    [733] = corrected[744];
assign input_data[745] = i_data   [734];
assign o_data    [734] = corrected[745];
assign input_data[746] = i_data   [735];
assign o_data    [735] = corrected[746];
assign input_data[747] = i_data   [736];
assign o_data    [736] = corrected[747];
assign input_data[748] = i_data   [737];
assign o_data    [737] = corrected[748];
assign input_data[749] = i_data   [738];
assign o_data    [738] = corrected[749];
assign input_data[750] = i_data   [739];
assign o_data    [739] = corrected[750];
assign input_data[751] = i_data   [740];
assign o_data    [740] = corrected[751];
assign input_data[752] = i_data   [741];
assign o_data    [741] = corrected[752];
assign input_data[753] = i_data   [742];
assign o_data    [742] = corrected[753];
assign input_data[754] = i_data   [743];
assign o_data    [743] = corrected[754];
assign input_data[755] = i_data   [744];
assign o_data    [744] = corrected[755];
assign input_data[756] = i_data   [745];
assign o_data    [745] = corrected[756];
assign input_data[757] = i_data   [746];
assign o_data    [746] = corrected[757];
assign input_data[758] = i_data   [747];
assign o_data    [747] = corrected[758];
assign input_data[759] = i_data   [748];
assign o_data    [748] = corrected[759];
assign input_data[760] = i_data   [749];
assign o_data    [749] = corrected[760];
assign input_data[761] = i_data   [750];
assign o_data    [750] = corrected[761];
assign input_data[762] = i_data   [751];
assign o_data    [751] = corrected[762];
assign input_data[763] = i_data   [752];
assign o_data    [752] = corrected[763];
assign input_data[764] = i_data   [753];
assign o_data    [753] = corrected[764];
assign input_data[765] = i_data   [754];
assign o_data    [754] = corrected[765];
assign input_data[766] = i_data   [755];
assign o_data    [755] = corrected[766];
assign input_data[767] = i_data   [756];
assign o_data    [756] = corrected[767];
assign input_data[768] = i_data   [757];
assign o_data    [757] = corrected[768];
assign input_data[769] = i_data   [758];
assign o_data    [758] = corrected[769];
assign input_data[770] = i_data   [759];
assign o_data    [759] = corrected[770];
assign input_data[771] = i_data   [760];
assign o_data    [760] = corrected[771];
assign input_data[772] = i_data   [761];
assign o_data    [761] = corrected[772];
assign input_data[773] = i_data   [762];
assign o_data    [762] = corrected[773];
assign input_data[774] = i_data   [763];
assign o_data    [763] = corrected[774];
assign input_data[775] = i_data   [764];
assign o_data    [764] = corrected[775];
assign input_data[776] = i_data   [765];
assign o_data    [765] = corrected[776];
assign input_data[777] = i_data   [766];
assign o_data    [766] = corrected[777];
assign input_data[778] = i_data   [767];
assign o_data    [767] = corrected[778];
assign input_data[779] = i_data   [768];
assign o_data    [768] = corrected[779];
assign input_data[780] = i_data   [769];
assign o_data    [769] = corrected[780];
assign input_data[781] = i_data   [770];
assign o_data    [770] = corrected[781];
assign input_data[782] = i_data   [771];
assign o_data    [771] = corrected[782];
assign input_data[783] = i_data   [772];
assign o_data    [772] = corrected[783];
assign input_data[784] = i_data   [773];
assign o_data    [773] = corrected[784];
assign input_data[785] = i_data   [774];
assign o_data    [774] = corrected[785];
assign input_data[786] = i_data   [775];
assign o_data    [775] = corrected[786];
assign input_data[787] = i_data   [776];
assign o_data    [776] = corrected[787];
assign input_data[788] = i_data   [777];
assign o_data    [777] = corrected[788];
assign input_data[789] = i_data   [778];
assign o_data    [778] = corrected[789];
assign input_data[790] = i_data   [779];
assign o_data    [779] = corrected[790];
assign input_data[791] = i_data   [780];
assign o_data    [780] = corrected[791];
assign input_data[792] = i_data   [781];
assign o_data    [781] = corrected[792];
assign input_data[793] = i_data   [782];
assign o_data    [782] = corrected[793];
assign input_data[794] = i_data   [783];
assign o_data    [783] = corrected[794];
assign input_data[795] = i_data   [784];
assign o_data    [784] = corrected[795];
assign input_data[796] = i_data   [785];
assign o_data    [785] = corrected[796];
assign input_data[797] = i_data   [786];
assign o_data    [786] = corrected[797];
assign input_data[798] = i_data   [787];
assign o_data    [787] = corrected[798];
assign input_data[799] = i_data   [788];
assign o_data    [788] = corrected[799];
assign input_data[800] = i_data   [789];
assign o_data    [789] = corrected[800];
assign input_data[801] = i_data   [790];
assign o_data    [790] = corrected[801];
assign input_data[802] = i_data   [791];
assign o_data    [791] = corrected[802];
assign input_data[803] = i_data   [792];
assign o_data    [792] = corrected[803];
assign input_data[804] = i_data   [793];
assign o_data    [793] = corrected[804];
assign input_data[805] = i_data   [794];
assign o_data    [794] = corrected[805];
assign input_data[806] = i_data   [795];
assign o_data    [795] = corrected[806];
assign input_data[807] = i_data   [796];
assign o_data    [796] = corrected[807];
assign input_data[808] = i_data   [797];
assign o_data    [797] = corrected[808];
assign input_data[809] = i_data   [798];
assign o_data    [798] = corrected[809];
assign input_data[810] = i_data   [799];
assign o_data    [799] = corrected[810];
assign input_data[811] = i_data   [800];
assign o_data    [800] = corrected[811];
assign input_data[812] = i_data   [801];
assign o_data    [801] = corrected[812];
assign input_data[813] = i_data   [802];
assign o_data    [802] = corrected[813];
assign input_data[814] = i_data   [803];
assign o_data    [803] = corrected[814];
assign input_data[815] = i_data   [804];
assign o_data    [804] = corrected[815];
assign input_data[816] = i_data   [805];
assign o_data    [805] = corrected[816];
assign input_data[817] = i_data   [806];
assign o_data    [806] = corrected[817];
assign input_data[818] = i_data   [807];
assign o_data    [807] = corrected[818];
assign input_data[819] = i_data   [808];
assign o_data    [808] = corrected[819];
assign input_data[820] = i_data   [809];
assign o_data    [809] = corrected[820];
assign input_data[821] = i_data   [810];
assign o_data    [810] = corrected[821];
assign input_data[822] = i_data   [811];
assign o_data    [811] = corrected[822];
assign input_data[823] = i_data   [812];
assign o_data    [812] = corrected[823];
assign input_data[824] = i_data   [813];
assign o_data    [813] = corrected[824];
assign input_data[825] = i_data   [814];
assign o_data    [814] = corrected[825];
assign input_data[826] = i_data   [815];
assign o_data    [815] = corrected[826];
assign input_data[827] = i_data   [816];
assign o_data    [816] = corrected[827];
assign input_data[828] = i_data   [817];
assign o_data    [817] = corrected[828];
assign input_data[829] = i_data   [818];
assign o_data    [818] = corrected[829];
assign input_data[830] = i_data   [819];
assign o_data    [819] = corrected[830];
assign input_data[831] = i_data   [820];
assign o_data    [820] = corrected[831];
assign input_data[832] = i_data   [821];
assign o_data    [821] = corrected[832];
assign input_data[833] = i_data   [822];
assign o_data    [822] = corrected[833];
assign input_data[834] = i_data   [823];
assign o_data    [823] = corrected[834];
assign input_data[835] = i_data   [824];
assign o_data    [824] = corrected[835];
assign input_data[836] = i_data   [825];
assign o_data    [825] = corrected[836];
assign input_data[837] = i_data   [826];
assign o_data    [826] = corrected[837];
assign input_data[838] = i_data   [827];
assign o_data    [827] = corrected[838];
assign input_data[839] = i_data   [828];
assign o_data    [828] = corrected[839];
assign input_data[840] = i_data   [829];
assign o_data    [829] = corrected[840];
assign input_data[841] = i_data   [830];
assign o_data    [830] = corrected[841];
assign input_data[842] = i_data   [831];
assign o_data    [831] = corrected[842];
assign input_data[843] = i_data   [832];
assign o_data    [832] = corrected[843];
assign input_data[844] = i_data   [833];
assign o_data    [833] = corrected[844];
assign input_data[845] = i_data   [834];
assign o_data    [834] = corrected[845];
assign input_data[846] = i_data   [835];
assign o_data    [835] = corrected[846];
assign input_data[847] = i_data   [836];
assign o_data    [836] = corrected[847];
assign input_data[848] = i_data   [837];
assign o_data    [837] = corrected[848];
assign input_data[849] = i_data   [838];
assign o_data    [838] = corrected[849];
assign input_data[850] = i_data   [839];
assign o_data    [839] = corrected[850];
assign input_data[851] = i_data   [840];
assign o_data    [840] = corrected[851];
assign input_data[852] = i_data   [841];
assign o_data    [841] = corrected[852];
assign input_data[853] = i_data   [842];
assign o_data    [842] = corrected[853];
assign input_data[854] = i_data   [843];
assign o_data    [843] = corrected[854];
assign input_data[855] = i_data   [844];
assign o_data    [844] = corrected[855];
assign input_data[856] = i_data   [845];
assign o_data    [845] = corrected[856];
assign input_data[857] = i_data   [846];
assign o_data    [846] = corrected[857];
assign input_data[858] = i_data   [847];
assign o_data    [847] = corrected[858];
assign input_data[859] = i_data   [848];
assign o_data    [848] = corrected[859];
assign input_data[860] = i_data   [849];
assign o_data    [849] = corrected[860];
assign input_data[861] = i_data   [850];
assign o_data    [850] = corrected[861];
assign input_data[862] = i_data   [851];
assign o_data    [851] = corrected[862];
assign input_data[863] = i_data   [852];
assign o_data    [852] = corrected[863];
assign input_data[864] = i_data   [853];
assign o_data    [853] = corrected[864];
assign input_data[865] = i_data   [854];
assign o_data    [854] = corrected[865];
assign input_data[866] = i_data   [855];
assign o_data    [855] = corrected[866];
assign input_data[867] = i_data   [856];
assign o_data    [856] = corrected[867];
assign input_data[868] = i_data   [857];
assign o_data    [857] = corrected[868];
assign input_data[869] = i_data   [858];
assign o_data    [858] = corrected[869];
assign input_data[870] = i_data   [859];
assign o_data    [859] = corrected[870];
assign input_data[871] = i_data   [860];
assign o_data    [860] = corrected[871];
assign input_data[872] = i_data   [861];
assign o_data    [861] = corrected[872];
assign input_data[873] = i_data   [862];
assign o_data    [862] = corrected[873];
assign input_data[874] = i_data   [863];
assign o_data    [863] = corrected[874];
assign input_data[875] = i_data   [864];
assign o_data    [864] = corrected[875];
assign input_data[876] = i_data   [865];
assign o_data    [865] = corrected[876];
assign input_data[877] = i_data   [866];
assign o_data    [866] = corrected[877];
assign input_data[878] = i_data   [867];
assign o_data    [867] = corrected[878];
assign input_data[879] = i_data   [868];
assign o_data    [868] = corrected[879];
assign input_data[880] = i_data   [869];
assign o_data    [869] = corrected[880];
assign input_data[881] = i_data   [870];
assign o_data    [870] = corrected[881];
assign input_data[882] = i_data   [871];
assign o_data    [871] = corrected[882];
assign input_data[883] = i_data   [872];
assign o_data    [872] = corrected[883];
assign input_data[884] = i_data   [873];
assign o_data    [873] = corrected[884];
assign input_data[885] = i_data   [874];
assign o_data    [874] = corrected[885];
assign input_data[886] = i_data   [875];
assign o_data    [875] = corrected[886];
assign input_data[887] = i_data   [876];
assign o_data    [876] = corrected[887];
assign input_data[888] = i_data   [877];
assign o_data    [877] = corrected[888];
assign input_data[889] = i_data   [878];
assign o_data    [878] = corrected[889];
assign input_data[890] = i_data   [879];
assign o_data    [879] = corrected[890];
assign input_data[891] = i_data   [880];
assign o_data    [880] = corrected[891];
assign input_data[892] = i_data   [881];
assign o_data    [881] = corrected[892];
assign input_data[893] = i_data   [882];
assign o_data    [882] = corrected[893];
assign input_data[894] = i_data   [883];
assign o_data    [883] = corrected[894];
assign input_data[895] = i_data   [884];
assign o_data    [884] = corrected[895];
assign input_data[896] = i_data   [885];
assign o_data    [885] = corrected[896];
assign input_data[897] = i_data   [886];
assign o_data    [886] = corrected[897];
assign input_data[898] = i_data   [887];
assign o_data    [887] = corrected[898];
assign input_data[899] = i_data   [888];
assign o_data    [888] = corrected[899];
assign input_data[900] = i_data   [889];
assign o_data    [889] = corrected[900];
assign input_data[901] = i_data   [890];
assign o_data    [890] = corrected[901];
assign input_data[902] = i_data   [891];
assign o_data    [891] = corrected[902];
assign input_data[903] = i_data   [892];
assign o_data    [892] = corrected[903];
assign input_data[904] = i_data   [893];
assign o_data    [893] = corrected[904];
assign input_data[905] = i_data   [894];
assign o_data    [894] = corrected[905];
assign input_data[906] = i_data   [895];
assign o_data    [895] = corrected[906];
assign input_data[907] = i_data   [896];
assign o_data    [896] = corrected[907];
assign input_data[908] = i_data   [897];
assign o_data    [897] = corrected[908];
assign input_data[909] = i_data   [898];
assign o_data    [898] = corrected[909];
assign input_data[910] = i_data   [899];
assign o_data    [899] = corrected[910];
assign input_data[911] = i_data   [900];
assign o_data    [900] = corrected[911];
assign input_data[912] = i_data   [901];
assign o_data    [901] = corrected[912];
assign input_data[913] = i_data   [902];
assign o_data    [902] = corrected[913];
assign input_data[914] = i_data   [903];
assign o_data    [903] = corrected[914];
assign input_data[915] = i_data   [904];
assign o_data    [904] = corrected[915];
assign input_data[916] = i_data   [905];
assign o_data    [905] = corrected[916];
assign input_data[917] = i_data   [906];
assign o_data    [906] = corrected[917];
assign input_data[918] = i_data   [907];
assign o_data    [907] = corrected[918];
assign input_data[919] = i_data   [908];
assign o_data    [908] = corrected[919];
assign input_data[920] = i_data   [909];
assign o_data    [909] = corrected[920];
assign input_data[921] = i_data   [910];
assign o_data    [910] = corrected[921];
assign input_data[922] = i_data   [911];
assign o_data    [911] = corrected[922];
assign input_data[923] = i_data   [912];
assign o_data    [912] = corrected[923];
assign input_data[924] = i_data   [913];
assign o_data    [913] = corrected[924];
assign input_data[925] = i_data   [914];
assign o_data    [914] = corrected[925];
assign input_data[926] = i_data   [915];
assign o_data    [915] = corrected[926];
assign input_data[927] = i_data   [916];
assign o_data    [916] = corrected[927];
assign input_data[928] = i_data   [917];
assign o_data    [917] = corrected[928];
assign input_data[929] = i_data   [918];
assign o_data    [918] = corrected[929];
assign input_data[930] = i_data   [919];
assign o_data    [919] = corrected[930];
assign input_data[931] = i_data   [920];
assign o_data    [920] = corrected[931];
assign input_data[932] = i_data   [921];
assign o_data    [921] = corrected[932];
assign input_data[933] = i_data   [922];
assign o_data    [922] = corrected[933];
assign input_data[934] = i_data   [923];
assign o_data    [923] = corrected[934];
assign input_data[935] = i_data   [924];
assign o_data    [924] = corrected[935];
assign input_data[936] = i_data   [925];
assign o_data    [925] = corrected[936];
assign input_data[937] = i_data   [926];
assign o_data    [926] = corrected[937];
assign input_data[938] = i_data   [927];
assign o_data    [927] = corrected[938];
assign input_data[939] = i_data   [928];
assign o_data    [928] = corrected[939];
assign input_data[940] = i_data   [929];
assign o_data    [929] = corrected[940];
assign input_data[941] = i_data   [930];
assign o_data    [930] = corrected[941];
assign input_data[942] = i_data   [931];
assign o_data    [931] = corrected[942];
assign input_data[943] = i_data   [932];
assign o_data    [932] = corrected[943];
assign input_data[944] = i_data   [933];
assign o_data    [933] = corrected[944];
assign input_data[945] = i_data   [934];
assign o_data    [934] = corrected[945];
assign input_data[946] = i_data   [935];
assign o_data    [935] = corrected[946];
assign input_data[947] = i_data   [936];
assign o_data    [936] = corrected[947];
assign input_data[948] = i_data   [937];
assign o_data    [937] = corrected[948];
assign input_data[949] = i_data   [938];
assign o_data    [938] = corrected[949];
assign input_data[950] = i_data   [939];
assign o_data    [939] = corrected[950];
assign input_data[951] = i_data   [940];
assign o_data    [940] = corrected[951];
assign input_data[952] = i_data   [941];
assign o_data    [941] = corrected[952];
assign input_data[953] = i_data   [942];
assign o_data    [942] = corrected[953];
assign input_data[954] = i_data   [943];
assign o_data    [943] = corrected[954];
assign input_data[955] = i_data   [944];
assign o_data    [944] = corrected[955];
assign input_data[956] = i_data   [945];
assign o_data    [945] = corrected[956];
assign input_data[957] = i_data   [946];
assign o_data    [946] = corrected[957];
assign input_data[958] = i_data   [947];
assign o_data    [947] = corrected[958];
assign input_data[959] = i_data   [948];
assign o_data    [948] = corrected[959];
assign input_data[960] = i_data   [949];
assign o_data    [949] = corrected[960];
assign input_data[961] = i_data   [950];
assign o_data    [950] = corrected[961];
assign input_data[962] = i_data   [951];
assign o_data    [951] = corrected[962];
assign input_data[963] = i_data   [952];
assign o_data    [952] = corrected[963];
assign input_data[964] = i_data   [953];
assign o_data    [953] = corrected[964];
assign input_data[965] = i_data   [954];
assign o_data    [954] = corrected[965];
assign input_data[966] = i_data   [955];
assign o_data    [955] = corrected[966];
assign input_data[967] = i_data   [956];
assign o_data    [956] = corrected[967];
assign input_data[968] = i_data   [957];
assign o_data    [957] = corrected[968];
assign input_data[969] = i_data   [958];
assign o_data    [958] = corrected[969];
assign input_data[970] = i_data   [959];
assign o_data    [959] = corrected[970];
assign input_data[971] = i_data   [960];
assign o_data    [960] = corrected[971];
assign input_data[972] = i_data   [961];
assign o_data    [961] = corrected[972];
assign input_data[973] = i_data   [962];
assign o_data    [962] = corrected[973];
assign input_data[974] = i_data   [963];
assign o_data    [963] = corrected[974];
assign input_data[975] = i_data   [964];
assign o_data    [964] = corrected[975];
assign input_data[976] = i_data   [965];
assign o_data    [965] = corrected[976];
assign input_data[977] = i_data   [966];
assign o_data    [966] = corrected[977];
assign input_data[978] = i_data   [967];
assign o_data    [967] = corrected[978];
assign input_data[979] = i_data   [968];
assign o_data    [968] = corrected[979];
assign input_data[980] = i_data   [969];
assign o_data    [969] = corrected[980];
assign input_data[981] = i_data   [970];
assign o_data    [970] = corrected[981];
assign input_data[982] = i_data   [971];
assign o_data    [971] = corrected[982];
assign input_data[983] = i_data   [972];
assign o_data    [972] = corrected[983];
assign input_data[984] = i_data   [973];
assign o_data    [973] = corrected[984];
assign input_data[985] = i_data   [974];
assign o_data    [974] = corrected[985];
assign input_data[986] = i_data   [975];
assign o_data    [975] = corrected[986];
assign input_data[987] = i_data   [976];
assign o_data    [976] = corrected[987];
assign input_data[988] = i_data   [977];
assign o_data    [977] = corrected[988];
assign input_data[989] = i_data   [978];
assign o_data    [978] = corrected[989];
assign input_data[990] = i_data   [979];
assign o_data    [979] = corrected[990];
assign input_data[991] = i_data   [980];
assign o_data    [980] = corrected[991];
assign input_data[992] = i_data   [981];
assign o_data    [981] = corrected[992];
assign input_data[993] = i_data   [982];
assign o_data    [982] = corrected[993];
assign input_data[994] = i_data   [983];
assign o_data    [983] = corrected[994];
assign input_data[995] = i_data   [984];
assign o_data    [984] = corrected[995];
assign input_data[996] = i_data   [985];
assign o_data    [985] = corrected[996];
assign input_data[997] = i_data   [986];
assign o_data    [986] = corrected[997];
assign input_data[998] = i_data   [987];
assign o_data    [987] = corrected[998];
assign input_data[999] = i_data   [988];
assign o_data    [988] = corrected[999];
assign input_data[1000] = i_data   [989];
assign o_data    [989] = corrected[1000];
assign input_data[1001] = i_data   [990];
assign o_data    [990] = corrected[1001];
assign input_data[1002] = i_data   [991];
assign o_data    [991] = corrected[1002];
assign input_data[1003] = i_data   [992];
assign o_data    [992] = corrected[1003];
assign input_data[1004] = i_data   [993];
assign o_data    [993] = corrected[1004];
assign input_data[1005] = i_data   [994];
assign o_data    [994] = corrected[1005];
assign input_data[1006] = i_data   [995];
assign o_data    [995] = corrected[1006];
assign input_data[1007] = i_data   [996];
assign o_data    [996] = corrected[1007];
assign input_data[1008] = i_data   [997];
assign o_data    [997] = corrected[1008];
assign input_data[1009] = i_data   [998];
assign o_data    [998] = corrected[1009];
assign input_data[1010] = i_data   [999];
assign o_data    [999] = corrected[1010];
assign input_data[1011] = i_data   [1000];
assign o_data    [1000] = corrected[1011];
assign input_data[1012] = i_data   [1001];
assign o_data    [1001] = corrected[1012];
assign input_data[1013] = i_data   [1002];
assign o_data    [1002] = corrected[1013];
assign input_data[1014] = i_data   [1003];
assign o_data    [1003] = corrected[1014];
assign input_data[1015] = i_data   [1004];
assign o_data    [1004] = corrected[1015];
assign input_data[1016] = i_data   [1005];
assign o_data    [1005] = corrected[1016];
assign input_data[1017] = i_data   [1006];
assign o_data    [1006] = corrected[1017];
assign input_data[1018] = i_data   [1007];
assign o_data    [1007] = corrected[1018];
assign input_data[1019] = i_data   [1008];
assign o_data    [1008] = corrected[1019];
assign input_data[1020] = i_data   [1009];
assign o_data    [1009] = corrected[1020];
assign input_data[1021] = i_data   [1010];
assign o_data    [1010] = corrected[1021];
assign input_data[1022] = i_data   [1011];
assign o_data    [1011] = corrected[1022];
assign input_data[1023] = i_data   [1012];
assign o_data    [1012] = corrected[1023];
assign syn_0000 = ecc_parity[0];
assign syn_0000_n = !(syn_0000); 
assign syn_0001 = ecc_parity[1];
assign syn_0001_n = !(syn_0001); 
assign syn_0002 = ecc_parity[2];
assign syn_0002_n = !(syn_0002); 
assign syn_0003 = ecc_parity[3];
assign syn_0003_n = !(syn_0003); 
assign syn_0004 = ecc_parity[4];
assign syn_0004_n = !(syn_0004); 
assign syn_0005 = ecc_parity[5];
assign syn_0005_n = !(syn_0005); 
assign syn_0006 = ecc_parity[6];
assign syn_0006_n = !(syn_0006); 
assign syn_0007 = ecc_parity[7];
assign syn_0007_n = !(syn_0007); 
assign syn_0008 = ecc_parity[8];
assign syn_0008_n = !(syn_0008); 
assign syn_0009 = ecc_parity[9];
assign syn_0009_n = !(syn_0009); 
assign nand0972 = !(syn_0002_n&syn_0001_n&syn_0000_n); 
assign nand0973 = !(syn_0002_n&syn_0001_n&syn_0000); 
assign nand0974 = !(syn_0002_n&syn_0001&syn_0000_n); 
assign nand0975 = !(syn_0002_n&syn_0001&syn_0000); 
assign nand0976 = !(syn_0002&syn_0001_n&syn_0000_n); 
assign nand0977 = !(syn_0002&syn_0001_n&syn_0000); 
assign nand0978 = !(syn_0002&syn_0001&syn_0000_n); 
assign nand0979 = !(syn_0002&syn_0001&syn_0000); 
assign nand0980 = !(syn_0003_n&syn_0005_n&syn_0004_n); 
assign nand0981 = !(syn_0003&syn_0005_n&syn_0004_n); 
assign nand0982 = !(syn_0003_n&syn_0004&syn_0005_n); 
assign nand0983 = !(syn_0004&syn_0003&syn_0005_n); 
assign nand0984 = !(syn_0003_n&syn_0005&syn_0004_n); 
assign nand0985 = !(syn_0003&syn_0005&syn_0004_n); 
assign nand0986 = !(syn_0003_n&syn_0004&syn_0005); 
assign nand0987 = !(syn_0004&syn_0003&syn_0005); 
assign nand0988 = !(syn_0008_n&syn_0007_n&syn_0006_n); 
assign nand0989 = !(syn_0008_n&syn_0006&syn_0007_n); 
assign nand0990 = !(syn_0007&syn_0008_n&syn_0006_n); 
assign nand0991 = !(syn_0007&syn_0008_n&syn_0006); 
assign nand0992 = !(syn_0007_n&syn_0006_n&syn_0008); 
assign nand0993 = !(syn_0006&syn_0007_n&syn_0008); 
assign nand0994 = !(syn_0007&syn_0006_n&syn_0008); 
assign nand0995 = !(syn_0007&syn_0006&syn_0008); 
assign nand0996 = !(syn_0009_n); 
assign nand0997 = !(syn_0009); 
assign nor0998 = !(nand0996|nand0980|nand0988|nand0972); 
assign invert0000 = nor0998;
assign nor0999 = !(nand0996|nand0980|nand0988|nand0973); 
assign invert0001 = nor0999;
assign nor1000 = !(nand0996|nand0974|nand0980|nand0988); 
assign invert0002 = nor1000;
assign nor1001 = !(nand0996|nand0980|nand0988|nand0975); 
assign invert0003 = nor1001;
assign nor1002 = !(nand0996|nand0980|nand0988|nand0976); 
assign invert0004 = nor1002;
assign nor1003 = !(nand0977|nand0996|nand0980|nand0988); 
assign invert0005 = nor1003;
assign nor1004 = !(nand0996|nand0980|nand0988|nand0978); 
assign invert0006 = nor1004;
assign nor1005 = !(nand0996|nand0979|nand0980|nand0988); 
assign invert0007 = nor1005;
assign nor1006 = !(nand0996|nand0988|nand0972|nand0981); 
assign invert0008 = nor1006;
assign nor1007 = !(nand0996|nand0988|nand0973|nand0981); 
assign invert0009 = nor1007;
assign nor1008 = !(nand0996|nand0974|nand0988|nand0981); 
assign invert0010 = nor1008;
assign nor1009 = !(nand0996|nand0988|nand0975|nand0981); 
assign invert0011 = nor1009;
assign nor1010 = !(nand0996|nand0988|nand0976|nand0981); 
assign invert0012 = nor1010;
assign nor1011 = !(nand0977|nand0996|nand0988|nand0981); 
assign invert0013 = nor1011;
assign nor1012 = !(nand0996|nand0988|nand0978|nand0981); 
assign invert0014 = nor1012;
assign nor1013 = !(nand0996|nand0979|nand0988|nand0981); 
assign invert0015 = nor1013;
assign nor1014 = !(nand0996|nand0988|nand0982|nand0972); 
assign invert0016 = nor1014;
assign nor1015 = !(nand0996|nand0988|nand0973|nand0982); 
assign invert0017 = nor1015;
assign nor1016 = !(nand0996|nand0974|nand0988|nand0982); 
assign invert0018 = nor1016;
assign nor1017 = !(nand0996|nand0988|nand0982|nand0975); 
assign invert0019 = nor1017;
assign nor1018 = !(nand0996|nand0988|nand0976|nand0982); 
assign invert0020 = nor1018;
assign nor1019 = !(nand0977|nand0996|nand0988|nand0982); 
assign invert0021 = nor1019;
assign nor1020 = !(nand0996|nand0988|nand0982|nand0978); 
assign invert0022 = nor1020;
assign nor1021 = !(nand0996|nand0979|nand0988|nand0982); 
assign invert0023 = nor1021;
assign nor1022 = !(nand0996|nand0983|nand0988|nand0972); 
assign invert0024 = nor1022;
assign nor1023 = !(nand0996|nand0983|nand0988|nand0973); 
assign invert0025 = nor1023;
assign nor1024 = !(nand0996|nand0974|nand0983|nand0988); 
assign invert0026 = nor1024;
assign nor1025 = !(nand0996|nand0983|nand0988|nand0975); 
assign invert0027 = nor1025;
assign nor1026 = !(nand0996|nand0983|nand0988|nand0976); 
assign invert0028 = nor1026;
assign nor1027 = !(nand0977|nand0996|nand0983|nand0988); 
assign invert0029 = nor1027;
assign nor1028 = !(nand0996|nand0983|nand0988|nand0978); 
assign invert0030 = nor1028;
assign nor1029 = !(nand0996|nand0983|nand0979|nand0988); 
assign invert0031 = nor1029;
assign nor1030 = !(nand0996|nand0988|nand0972|nand0984); 
assign invert0032 = nor1030;
assign nor1031 = !(nand0996|nand0988|nand0973|nand0984); 
assign invert0033 = nor1031;
assign nor1032 = !(nand0996|nand0974|nand0988|nand0984); 
assign invert0034 = nor1032;
assign nor1033 = !(nand0996|nand0988|nand0975|nand0984); 
assign invert0035 = nor1033;
assign nor1034 = !(nand0996|nand0988|nand0976|nand0984); 
assign invert0036 = nor1034;
assign nor1035 = !(nand0977|nand0996|nand0988|nand0984); 
assign invert0037 = nor1035;
assign nor1036 = !(nand0996|nand0988|nand0978|nand0984); 
assign invert0038 = nor1036;
assign nor1037 = !(nand0996|nand0979|nand0988|nand0984); 
assign invert0039 = nor1037;
assign nor1038 = !(nand0996|nand0988|nand0985|nand0972); 
assign invert0040 = nor1038;
assign nor1039 = !(nand0996|nand0988|nand0973|nand0985); 
assign invert0041 = nor1039;
assign nor1040 = !(nand0996|nand0974|nand0988|nand0985); 
assign invert0042 = nor1040;
assign nor1041 = !(nand0996|nand0988|nand0985|nand0975); 
assign invert0043 = nor1041;
assign nor1042 = !(nand0996|nand0988|nand0976|nand0985); 
assign invert0044 = nor1042;
assign nor1043 = !(nand0977|nand0996|nand0988|nand0985); 
assign invert0045 = nor1043;
assign nor1044 = !(nand0996|nand0988|nand0985|nand0978); 
assign invert0046 = nor1044;
assign nor1045 = !(nand0996|nand0979|nand0988|nand0985); 
assign invert0047 = nor1045;
assign nor1046 = !(nand0996|nand0986|nand0988|nand0972); 
assign invert0048 = nor1046;
assign nor1047 = !(nand0996|nand0986|nand0988|nand0973); 
assign invert0049 = nor1047;
assign nor1048 = !(nand0996|nand0986|nand0974|nand0988); 
assign invert0050 = nor1048;
assign nor1049 = !(nand0996|nand0986|nand0988|nand0975); 
assign invert0051 = nor1049;
assign nor1050 = !(nand0996|nand0986|nand0988|nand0976); 
assign invert0052 = nor1050;
assign nor1051 = !(nand0977|nand0996|nand0986|nand0988); 
assign invert0053 = nor1051;
assign nor1052 = !(nand0996|nand0986|nand0988|nand0978); 
assign invert0054 = nor1052;
assign nor1053 = !(nand0996|nand0986|nand0979|nand0988); 
assign invert0055 = nor1053;
assign nor1054 = !(nand0996|nand0988|nand0987|nand0972); 
assign invert0056 = nor1054;
assign nor1055 = !(nand0996|nand0988|nand0973|nand0987); 
assign invert0057 = nor1055;
assign nor1056 = !(nand0996|nand0974|nand0988|nand0987); 
assign invert0058 = nor1056;
assign nor1057 = !(nand0996|nand0988|nand0987|nand0975); 
assign invert0059 = nor1057;
assign nor1058 = !(nand0996|nand0988|nand0976|nand0987); 
assign invert0060 = nor1058;
assign nor1059 = !(nand0977|nand0996|nand0988|nand0987); 
assign invert0061 = nor1059;
assign nor1060 = !(nand0996|nand0988|nand0978|nand0987); 
assign invert0062 = nor1060;
assign nor1061 = !(nand0996|nand0979|nand0988|nand0987); 
assign invert0063 = nor1061;
assign nor1062 = !(nand0989|nand0996|nand0980|nand0972); 
assign invert0064 = nor1062;
assign nor1063 = !(nand0989|nand0996|nand0980|nand0973); 
assign invert0065 = nor1063;
assign nor1064 = !(nand0989|nand0996|nand0974|nand0980); 
assign invert0066 = nor1064;
assign nor1065 = !(nand0989|nand0996|nand0980|nand0975); 
assign invert0067 = nor1065;
assign nor1066 = !(nand0989|nand0996|nand0980|nand0976); 
assign invert0068 = nor1066;
assign nor1067 = !(nand0989|nand0977|nand0996|nand0980); 
assign invert0069 = nor1067;
assign nor1068 = !(nand0989|nand0996|nand0980|nand0978); 
assign invert0070 = nor1068;
assign nor1069 = !(nand0989|nand0996|nand0979|nand0980); 
assign invert0071 = nor1069;
assign nor1070 = !(nand0989|nand0996|nand0972|nand0981); 
assign invert0072 = nor1070;
assign nor1071 = !(nand0989|nand0996|nand0973|nand0981); 
assign invert0073 = nor1071;
assign nor1072 = !(nand0989|nand0996|nand0974|nand0981); 
assign invert0074 = nor1072;
assign nor1073 = !(nand0989|nand0996|nand0975|nand0981); 
assign invert0075 = nor1073;
assign nor1074 = !(nand0989|nand0996|nand0976|nand0981); 
assign invert0076 = nor1074;
assign nor1075 = !(nand0989|nand0977|nand0996|nand0981); 
assign invert0077 = nor1075;
assign nor1076 = !(nand0989|nand0996|nand0978|nand0981); 
assign invert0078 = nor1076;
assign nor1077 = !(nand0989|nand0996|nand0979|nand0981); 
assign invert0079 = nor1077;
assign nor1078 = !(nand0989|nand0996|nand0982|nand0972); 
assign invert0080 = nor1078;
assign nor1079 = !(nand0989|nand0996|nand0973|nand0982); 
assign invert0081 = nor1079;
assign nor1080 = !(nand0989|nand0996|nand0974|nand0982); 
assign invert0082 = nor1080;
assign nor1081 = !(nand0989|nand0996|nand0982|nand0975); 
assign invert0083 = nor1081;
assign nor1082 = !(nand0989|nand0996|nand0976|nand0982); 
assign invert0084 = nor1082;
assign nor1083 = !(nand0989|nand0977|nand0996|nand0982); 
assign invert0085 = nor1083;
assign nor1084 = !(nand0989|nand0996|nand0982|nand0978); 
assign invert0086 = nor1084;
assign nor1085 = !(nand0989|nand0996|nand0979|nand0982); 
assign invert0087 = nor1085;
assign nor1086 = !(nand0989|nand0996|nand0983|nand0972); 
assign invert0088 = nor1086;
assign nor1087 = !(nand0989|nand0996|nand0983|nand0973); 
assign invert0089 = nor1087;
assign nor1088 = !(nand0989|nand0996|nand0974|nand0983); 
assign invert0090 = nor1088;
assign nor1089 = !(nand0989|nand0996|nand0983|nand0975); 
assign invert0091 = nor1089;
assign nor1090 = !(nand0989|nand0996|nand0983|nand0976); 
assign invert0092 = nor1090;
assign nor1091 = !(nand0989|nand0977|nand0996|nand0983); 
assign invert0093 = nor1091;
assign nor1092 = !(nand0989|nand0996|nand0983|nand0978); 
assign invert0094 = nor1092;
assign nor1093 = !(nand0989|nand0996|nand0983|nand0979); 
assign invert0095 = nor1093;
assign nor1094 = !(nand0989|nand0996|nand0972|nand0984); 
assign invert0096 = nor1094;
assign nor1095 = !(nand0989|nand0996|nand0973|nand0984); 
assign invert0097 = nor1095;
assign nor1096 = !(nand0989|nand0996|nand0974|nand0984); 
assign invert0098 = nor1096;
assign nor1097 = !(nand0989|nand0996|nand0975|nand0984); 
assign invert0099 = nor1097;
assign nor1098 = !(nand0989|nand0996|nand0976|nand0984); 
assign invert0100 = nor1098;
assign nor1099 = !(nand0989|nand0977|nand0996|nand0984); 
assign invert0101 = nor1099;
assign nor1100 = !(nand0989|nand0996|nand0978|nand0984); 
assign invert0102 = nor1100;
assign nor1101 = !(nand0989|nand0996|nand0979|nand0984); 
assign invert0103 = nor1101;
assign nor1102 = !(nand0989|nand0996|nand0985|nand0972); 
assign invert0104 = nor1102;
assign nor1103 = !(nand0989|nand0996|nand0973|nand0985); 
assign invert0105 = nor1103;
assign nor1104 = !(nand0989|nand0996|nand0974|nand0985); 
assign invert0106 = nor1104;
assign nor1105 = !(nand0989|nand0996|nand0985|nand0975); 
assign invert0107 = nor1105;
assign nor1106 = !(nand0989|nand0996|nand0976|nand0985); 
assign invert0108 = nor1106;
assign nor1107 = !(nand0989|nand0977|nand0996|nand0985); 
assign invert0109 = nor1107;
assign nor1108 = !(nand0989|nand0996|nand0985|nand0978); 
assign invert0110 = nor1108;
assign nor1109 = !(nand0989|nand0996|nand0979|nand0985); 
assign invert0111 = nor1109;
assign nor1110 = !(nand0989|nand0996|nand0986|nand0972); 
assign invert0112 = nor1110;
assign nor1111 = !(nand0989|nand0996|nand0986|nand0973); 
assign invert0113 = nor1111;
assign nor1112 = !(nand0989|nand0996|nand0986|nand0974); 
assign invert0114 = nor1112;
assign nor1113 = !(nand0989|nand0996|nand0986|nand0975); 
assign invert0115 = nor1113;
assign nor1114 = !(nand0989|nand0996|nand0986|nand0976); 
assign invert0116 = nor1114;
assign nor1115 = !(nand0989|nand0977|nand0996|nand0986); 
assign invert0117 = nor1115;
assign nor1116 = !(nand0989|nand0996|nand0986|nand0978); 
assign invert0118 = nor1116;
assign nor1117 = !(nand0989|nand0996|nand0986|nand0979); 
assign invert0119 = nor1117;
assign nor1118 = !(nand0989|nand0996|nand0987|nand0972); 
assign invert0120 = nor1118;
assign nor1119 = !(nand0989|nand0996|nand0973|nand0987); 
assign invert0121 = nor1119;
assign nor1120 = !(nand0989|nand0996|nand0974|nand0987); 
assign invert0122 = nor1120;
assign nor1121 = !(nand0989|nand0996|nand0987|nand0975); 
assign invert0123 = nor1121;
assign nor1122 = !(nand0989|nand0996|nand0976|nand0987); 
assign invert0124 = nor1122;
assign nor1123 = !(nand0989|nand0977|nand0996|nand0987); 
assign invert0125 = nor1123;
assign nor1124 = !(nand0989|nand0996|nand0978|nand0987); 
assign invert0126 = nor1124;
assign nor1125 = !(nand0989|nand0996|nand0979|nand0987); 
assign invert0127 = nor1125;
assign nor1126 = !(nand0996|nand0990|nand0980|nand0972); 
assign invert0128 = nor1126;
assign nor1127 = !(nand0996|nand0990|nand0980|nand0973); 
assign invert0129 = nor1127;
assign nor1128 = !(nand0996|nand0974|nand0990|nand0980); 
assign invert0130 = nor1128;
assign nor1129 = !(nand0996|nand0990|nand0980|nand0975); 
assign invert0131 = nor1129;
assign nor1130 = !(nand0996|nand0990|nand0980|nand0976); 
assign invert0132 = nor1130;
assign nor1131 = !(nand0977|nand0996|nand0990|nand0980); 
assign invert0133 = nor1131;
assign nor1132 = !(nand0996|nand0990|nand0980|nand0978); 
assign invert0134 = nor1132;
assign nor1133 = !(nand0996|nand0990|nand0979|nand0980); 
assign invert0135 = nor1133;
assign nor1134 = !(nand0996|nand0990|nand0972|nand0981); 
assign invert0136 = nor1134;
assign nor1135 = !(nand0996|nand0990|nand0973|nand0981); 
assign invert0137 = nor1135;
assign nor1136 = !(nand0996|nand0974|nand0990|nand0981); 
assign invert0138 = nor1136;
assign nor1137 = !(nand0996|nand0990|nand0975|nand0981); 
assign invert0139 = nor1137;
assign nor1138 = !(nand0996|nand0990|nand0976|nand0981); 
assign invert0140 = nor1138;
assign nor1139 = !(nand0977|nand0996|nand0990|nand0981); 
assign invert0141 = nor1139;
assign nor1140 = !(nand0996|nand0990|nand0978|nand0981); 
assign invert0142 = nor1140;
assign nor1141 = !(nand0996|nand0990|nand0979|nand0981); 
assign invert0143 = nor1141;
assign nor1142 = !(nand0996|nand0990|nand0982|nand0972); 
assign invert0144 = nor1142;
assign nor1143 = !(nand0996|nand0990|nand0973|nand0982); 
assign invert0145 = nor1143;
assign nor1144 = !(nand0996|nand0974|nand0990|nand0982); 
assign invert0146 = nor1144;
assign nor1145 = !(nand0996|nand0990|nand0982|nand0975); 
assign invert0147 = nor1145;
assign nor1146 = !(nand0996|nand0990|nand0976|nand0982); 
assign invert0148 = nor1146;
assign nor1147 = !(nand0977|nand0996|nand0990|nand0982); 
assign invert0149 = nor1147;
assign nor1148 = !(nand0996|nand0990|nand0982|nand0978); 
assign invert0150 = nor1148;
assign nor1149 = !(nand0996|nand0990|nand0979|nand0982); 
assign invert0151 = nor1149;
assign nor1150 = !(nand0996|nand0983|nand0990|nand0972); 
assign invert0152 = nor1150;
assign nor1151 = !(nand0996|nand0983|nand0990|nand0973); 
assign invert0153 = nor1151;
assign nor1152 = !(nand0996|nand0974|nand0983|nand0990); 
assign invert0154 = nor1152;
assign nor1153 = !(nand0996|nand0983|nand0990|nand0975); 
assign invert0155 = nor1153;
assign nor1154 = !(nand0996|nand0983|nand0990|nand0976); 
assign invert0156 = nor1154;
assign nor1155 = !(nand0977|nand0996|nand0983|nand0990); 
assign invert0157 = nor1155;
assign nor1156 = !(nand0996|nand0983|nand0990|nand0978); 
assign invert0158 = nor1156;
assign nor1157 = !(nand0996|nand0983|nand0990|nand0979); 
assign invert0159 = nor1157;
assign nor1158 = !(nand0996|nand0990|nand0972|nand0984); 
assign invert0160 = nor1158;
assign nor1159 = !(nand0996|nand0990|nand0973|nand0984); 
assign invert0161 = nor1159;
assign nor1160 = !(nand0996|nand0974|nand0990|nand0984); 
assign invert0162 = nor1160;
assign nor1161 = !(nand0996|nand0990|nand0975|nand0984); 
assign invert0163 = nor1161;
assign nor1162 = !(nand0996|nand0990|nand0976|nand0984); 
assign invert0164 = nor1162;
assign nor1163 = !(nand0977|nand0996|nand0990|nand0984); 
assign invert0165 = nor1163;
assign nor1164 = !(nand0996|nand0990|nand0978|nand0984); 
assign invert0166 = nor1164;
assign nor1165 = !(nand0996|nand0990|nand0979|nand0984); 
assign invert0167 = nor1165;
assign nor1166 = !(nand0996|nand0990|nand0985|nand0972); 
assign invert0168 = nor1166;
assign nor1167 = !(nand0996|nand0990|nand0973|nand0985); 
assign invert0169 = nor1167;
assign nor1168 = !(nand0996|nand0974|nand0990|nand0985); 
assign invert0170 = nor1168;
assign nor1169 = !(nand0996|nand0990|nand0985|nand0975); 
assign invert0171 = nor1169;
assign nor1170 = !(nand0996|nand0990|nand0976|nand0985); 
assign invert0172 = nor1170;
assign nor1171 = !(nand0977|nand0996|nand0990|nand0985); 
assign invert0173 = nor1171;
assign nor1172 = !(nand0996|nand0990|nand0985|nand0978); 
assign invert0174 = nor1172;
assign nor1173 = !(nand0996|nand0990|nand0979|nand0985); 
assign invert0175 = nor1173;
assign nor1174 = !(nand0996|nand0986|nand0990|nand0972); 
assign invert0176 = nor1174;
assign nor1175 = !(nand0996|nand0986|nand0990|nand0973); 
assign invert0177 = nor1175;
assign nor1176 = !(nand0996|nand0986|nand0974|nand0990); 
assign invert0178 = nor1176;
assign nor1177 = !(nand0996|nand0986|nand0990|nand0975); 
assign invert0179 = nor1177;
assign nor1178 = !(nand0996|nand0986|nand0990|nand0976); 
assign invert0180 = nor1178;
assign nor1179 = !(nand0977|nand0996|nand0986|nand0990); 
assign invert0181 = nor1179;
assign nor1180 = !(nand0996|nand0986|nand0990|nand0978); 
assign invert0182 = nor1180;
assign nor1181 = !(nand0996|nand0986|nand0990|nand0979); 
assign invert0183 = nor1181;
assign nor1182 = !(nand0996|nand0990|nand0987|nand0972); 
assign invert0184 = nor1182;
assign nor1183 = !(nand0996|nand0990|nand0973|nand0987); 
assign invert0185 = nor1183;
assign nor1184 = !(nand0996|nand0974|nand0990|nand0987); 
assign invert0186 = nor1184;
assign nor1185 = !(nand0996|nand0990|nand0987|nand0975); 
assign invert0187 = nor1185;
assign nor1186 = !(nand0996|nand0990|nand0976|nand0987); 
assign invert0188 = nor1186;
assign nor1187 = !(nand0977|nand0996|nand0990|nand0987); 
assign invert0189 = nor1187;
assign nor1188 = !(nand0996|nand0990|nand0978|nand0987); 
assign invert0190 = nor1188;
assign nor1189 = !(nand0996|nand0990|nand0979|nand0987); 
assign invert0191 = nor1189;
assign nor1190 = !(nand0996|nand0980|nand0972|nand0991); 
assign invert0192 = nor1190;
assign nor1191 = !(nand0996|nand0980|nand0973|nand0991); 
assign invert0193 = nor1191;
assign nor1192 = !(nand0996|nand0974|nand0980|nand0991); 
assign invert0194 = nor1192;
assign nor1193 = !(nand0996|nand0980|nand0975|nand0991); 
assign invert0195 = nor1193;
assign nor1194 = !(nand0996|nand0980|nand0976|nand0991); 
assign invert0196 = nor1194;
assign nor1195 = !(nand0977|nand0996|nand0980|nand0991); 
assign invert0197 = nor1195;
assign nor1196 = !(nand0996|nand0980|nand0978|nand0991); 
assign invert0198 = nor1196;
assign nor1197 = !(nand0996|nand0979|nand0980|nand0991); 
assign invert0199 = nor1197;
assign nor1198 = !(nand0996|nand0972|nand0991|nand0981); 
assign invert0200 = nor1198;
assign nor1199 = !(nand0996|nand0973|nand0991|nand0981); 
assign invert0201 = nor1199;
assign nor1200 = !(nand0996|nand0974|nand0991|nand0981); 
assign invert0202 = nor1200;
assign nor1201 = !(nand0996|nand0975|nand0991|nand0981); 
assign invert0203 = nor1201;
assign nor1202 = !(nand0996|nand0976|nand0991|nand0981); 
assign invert0204 = nor1202;
assign nor1203 = !(nand0977|nand0996|nand0991|nand0981); 
assign invert0205 = nor1203;
assign nor1204 = !(nand0996|nand0978|nand0991|nand0981); 
assign invert0206 = nor1204;
assign nor1205 = !(nand0996|nand0979|nand0991|nand0981); 
assign invert0207 = nor1205;
assign nor1206 = !(nand0996|nand0982|nand0972|nand0991); 
assign invert0208 = nor1206;
assign nor1207 = !(nand0996|nand0973|nand0982|nand0991); 
assign invert0209 = nor1207;
assign nor1208 = !(nand0996|nand0974|nand0982|nand0991); 
assign invert0210 = nor1208;
assign nor1209 = !(nand0996|nand0982|nand0975|nand0991); 
assign invert0211 = nor1209;
assign nor1210 = !(nand0996|nand0976|nand0982|nand0991); 
assign invert0212 = nor1210;
assign nor1211 = !(nand0977|nand0996|nand0982|nand0991); 
assign invert0213 = nor1211;
assign nor1212 = !(nand0996|nand0982|nand0978|nand0991); 
assign invert0214 = nor1212;
assign nor1213 = !(nand0996|nand0979|nand0982|nand0991); 
assign invert0215 = nor1213;
assign nor1214 = !(nand0996|nand0983|nand0972|nand0991); 
assign invert0216 = nor1214;
assign nor1215 = !(nand0996|nand0983|nand0973|nand0991); 
assign invert0217 = nor1215;
assign nor1216 = !(nand0996|nand0974|nand0983|nand0991); 
assign invert0218 = nor1216;
assign nor1217 = !(nand0996|nand0983|nand0975|nand0991); 
assign invert0219 = nor1217;
assign nor1218 = !(nand0996|nand0983|nand0976|nand0991); 
assign invert0220 = nor1218;
assign nor1219 = !(nand0977|nand0996|nand0983|nand0991); 
assign invert0221 = nor1219;
assign nor1220 = !(nand0996|nand0983|nand0978|nand0991); 
assign invert0222 = nor1220;
assign nor1221 = !(nand0996|nand0983|nand0979|nand0991); 
assign invert0223 = nor1221;
assign nor1222 = !(nand0996|nand0972|nand0984|nand0991); 
assign invert0224 = nor1222;
assign nor1223 = !(nand0996|nand0973|nand0984|nand0991); 
assign invert0225 = nor1223;
assign nor1224 = !(nand0996|nand0974|nand0984|nand0991); 
assign invert0226 = nor1224;
assign nor1225 = !(nand0996|nand0975|nand0984|nand0991); 
assign invert0227 = nor1225;
assign nor1226 = !(nand0996|nand0976|nand0984|nand0991); 
assign invert0228 = nor1226;
assign nor1227 = !(nand0977|nand0996|nand0984|nand0991); 
assign invert0229 = nor1227;
assign nor1228 = !(nand0996|nand0978|nand0984|nand0991); 
assign invert0230 = nor1228;
assign nor1229 = !(nand0996|nand0979|nand0984|nand0991); 
assign invert0231 = nor1229;
assign nor1230 = !(nand0996|nand0985|nand0972|nand0991); 
assign invert0232 = nor1230;
assign nor1231 = !(nand0996|nand0973|nand0985|nand0991); 
assign invert0233 = nor1231;
assign nor1232 = !(nand0996|nand0974|nand0985|nand0991); 
assign invert0234 = nor1232;
assign nor1233 = !(nand0996|nand0985|nand0975|nand0991); 
assign invert0235 = nor1233;
assign nor1234 = !(nand0996|nand0976|nand0985|nand0991); 
assign invert0236 = nor1234;
assign nor1235 = !(nand0977|nand0996|nand0985|nand0991); 
assign invert0237 = nor1235;
assign nor1236 = !(nand0996|nand0985|nand0978|nand0991); 
assign invert0238 = nor1236;
assign nor1237 = !(nand0996|nand0979|nand0985|nand0991); 
assign invert0239 = nor1237;
assign nor1238 = !(nand0996|nand0986|nand0972|nand0991); 
assign invert0240 = nor1238;
assign nor1239 = !(nand0996|nand0986|nand0973|nand0991); 
assign invert0241 = nor1239;
assign nor1240 = !(nand0996|nand0986|nand0974|nand0991); 
assign invert0242 = nor1240;
assign nor1241 = !(nand0996|nand0986|nand0975|nand0991); 
assign invert0243 = nor1241;
assign nor1242 = !(nand0996|nand0986|nand0976|nand0991); 
assign invert0244 = nor1242;
assign nor1243 = !(nand0977|nand0996|nand0986|nand0991); 
assign invert0245 = nor1243;
assign nor1244 = !(nand0996|nand0986|nand0978|nand0991); 
assign invert0246 = nor1244;
assign nor1245 = !(nand0996|nand0986|nand0979|nand0991); 
assign invert0247 = nor1245;
assign nor1246 = !(nand0996|nand0987|nand0972|nand0991); 
assign invert0248 = nor1246;
assign nor1247 = !(nand0996|nand0973|nand0987|nand0991); 
assign invert0249 = nor1247;
assign nor1248 = !(nand0996|nand0974|nand0987|nand0991); 
assign invert0250 = nor1248;
assign nor1249 = !(nand0996|nand0987|nand0975|nand0991); 
assign invert0251 = nor1249;
assign nor1250 = !(nand0996|nand0976|nand0987|nand0991); 
assign invert0252 = nor1250;
assign nor1251 = !(nand0977|nand0996|nand0987|nand0991); 
assign invert0253 = nor1251;
assign nor1252 = !(nand0996|nand0978|nand0987|nand0991); 
assign invert0254 = nor1252;
assign nor1253 = !(nand0996|nand0979|nand0987|nand0991); 
assign invert0255 = nor1253;
assign nor1254 = !(nand0996|nand0980|nand0992|nand0972); 
assign invert0256 = nor1254;
assign nor1255 = !(nand0996|nand0980|nand0973|nand0992); 
assign invert0257 = nor1255;
assign nor1256 = !(nand0996|nand0974|nand0980|nand0992); 
assign invert0258 = nor1256;
assign nor1257 = !(nand0996|nand0980|nand0992|nand0975); 
assign invert0259 = nor1257;
assign nor1258 = !(nand0996|nand0980|nand0976|nand0992); 
assign invert0260 = nor1258;
assign nor1259 = !(nand0977|nand0996|nand0980|nand0992); 
assign invert0261 = nor1259;
assign nor1260 = !(nand0996|nand0980|nand0992|nand0978); 
assign invert0262 = nor1260;
assign nor1261 = !(nand0996|nand0979|nand0980|nand0992); 
assign invert0263 = nor1261;
assign nor1262 = !(nand0996|nand0992|nand0972|nand0981); 
assign invert0264 = nor1262;
assign nor1263 = !(nand0996|nand0973|nand0992|nand0981); 
assign invert0265 = nor1263;
assign nor1264 = !(nand0996|nand0974|nand0992|nand0981); 
assign invert0266 = nor1264;
assign nor1265 = !(nand0996|nand0992|nand0975|nand0981); 
assign invert0267 = nor1265;
assign nor1266 = !(nand0996|nand0976|nand0992|nand0981); 
assign invert0268 = nor1266;
assign nor1267 = !(nand0977|nand0996|nand0992|nand0981); 
assign invert0269 = nor1267;
assign nor1268 = !(nand0996|nand0992|nand0978|nand0981); 
assign invert0270 = nor1268;
assign nor1269 = !(nand0996|nand0979|nand0992|nand0981); 
assign invert0271 = nor1269;
assign nor1270 = !(nand0996|nand0992|nand0982|nand0972); 
assign invert0272 = nor1270;
assign nor1271 = !(nand0996|nand0973|nand0992|nand0982); 
assign invert0273 = nor1271;
assign nor1272 = !(nand0996|nand0974|nand0992|nand0982); 
assign invert0274 = nor1272;
assign nor1273 = !(nand0996|nand0992|nand0982|nand0975); 
assign invert0275 = nor1273;
assign nor1274 = !(nand0996|nand0976|nand0992|nand0982); 
assign invert0276 = nor1274;
assign nor1275 = !(nand0977|nand0996|nand0992|nand0982); 
assign invert0277 = nor1275;
assign nor1276 = !(nand0996|nand0992|nand0982|nand0978); 
assign invert0278 = nor1276;
assign nor1277 = !(nand0996|nand0979|nand0992|nand0982); 
assign invert0279 = nor1277;
assign nor1278 = !(nand0996|nand0983|nand0992|nand0972); 
assign invert0280 = nor1278;
assign nor1279 = !(nand0996|nand0983|nand0973|nand0992); 
assign invert0281 = nor1279;
assign nor1280 = !(nand0996|nand0974|nand0983|nand0992); 
assign invert0282 = nor1280;
assign nor1281 = !(nand0996|nand0983|nand0992|nand0975); 
assign invert0283 = nor1281;
assign nor1282 = !(nand0996|nand0983|nand0976|nand0992); 
assign invert0284 = nor1282;
assign nor1283 = !(nand0977|nand0996|nand0983|nand0992); 
assign invert0285 = nor1283;
assign nor1284 = !(nand0996|nand0983|nand0992|nand0978); 
assign invert0286 = nor1284;
assign nor1285 = !(nand0996|nand0983|nand0979|nand0992); 
assign invert0287 = nor1285;
assign nor1286 = !(nand0996|nand0992|nand0972|nand0984); 
assign invert0288 = nor1286;
assign nor1287 = !(nand0996|nand0973|nand0992|nand0984); 
assign invert0289 = nor1287;
assign nor1288 = !(nand0996|nand0974|nand0992|nand0984); 
assign invert0290 = nor1288;
assign nor1289 = !(nand0996|nand0992|nand0975|nand0984); 
assign invert0291 = nor1289;
assign nor1290 = !(nand0996|nand0976|nand0992|nand0984); 
assign invert0292 = nor1290;
assign nor1291 = !(nand0977|nand0996|nand0992|nand0984); 
assign invert0293 = nor1291;
assign nor1292 = !(nand0996|nand0992|nand0978|nand0984); 
assign invert0294 = nor1292;
assign nor1293 = !(nand0996|nand0979|nand0992|nand0984); 
assign invert0295 = nor1293;
assign nor1294 = !(nand0996|nand0985|nand0992|nand0972); 
assign invert0296 = nor1294;
assign nor1295 = !(nand0996|nand0973|nand0985|nand0992); 
assign invert0297 = nor1295;
assign nor1296 = !(nand0996|nand0974|nand0985|nand0992); 
assign invert0298 = nor1296;
assign nor1297 = !(nand0996|nand0985|nand0992|nand0975); 
assign invert0299 = nor1297;
assign nor1298 = !(nand0996|nand0976|nand0985|nand0992); 
assign invert0300 = nor1298;
assign nor1299 = !(nand0977|nand0996|nand0985|nand0992); 
assign invert0301 = nor1299;
assign nor1300 = !(nand0996|nand0985|nand0992|nand0978); 
assign invert0302 = nor1300;
assign nor1301 = !(nand0996|nand0979|nand0985|nand0992); 
assign invert0303 = nor1301;
assign nor1302 = !(nand0996|nand0986|nand0992|nand0972); 
assign invert0304 = nor1302;
assign nor1303 = !(nand0996|nand0986|nand0973|nand0992); 
assign invert0305 = nor1303;
assign nor1304 = !(nand0996|nand0986|nand0974|nand0992); 
assign invert0306 = nor1304;
assign nor1305 = !(nand0996|nand0986|nand0992|nand0975); 
assign invert0307 = nor1305;
assign nor1306 = !(nand0996|nand0986|nand0976|nand0992); 
assign invert0308 = nor1306;
assign nor1307 = !(nand0977|nand0996|nand0986|nand0992); 
assign invert0309 = nor1307;
assign nor1308 = !(nand0996|nand0986|nand0992|nand0978); 
assign invert0310 = nor1308;
assign nor1309 = !(nand0996|nand0986|nand0979|nand0992); 
assign invert0311 = nor1309;
assign nor1310 = !(nand0996|nand0992|nand0987|nand0972); 
assign invert0312 = nor1310;
assign nor1311 = !(nand0996|nand0973|nand0992|nand0987); 
assign invert0313 = nor1311;
assign nor1312 = !(nand0996|nand0974|nand0992|nand0987); 
assign invert0314 = nor1312;
assign nor1313 = !(nand0996|nand0992|nand0987|nand0975); 
assign invert0315 = nor1313;
assign nor1314 = !(nand0996|nand0976|nand0992|nand0987); 
assign invert0316 = nor1314;
assign nor1315 = !(nand0977|nand0996|nand0992|nand0987); 
assign invert0317 = nor1315;
assign nor1316 = !(nand0996|nand0992|nand0978|nand0987); 
assign invert0318 = nor1316;
assign nor1317 = !(nand0996|nand0979|nand0992|nand0987); 
assign invert0319 = nor1317;
assign nor1318 = !(nand0996|nand0993|nand0980|nand0972); 
assign invert0320 = nor1318;
assign nor1319 = !(nand0996|nand0993|nand0980|nand0973); 
assign invert0321 = nor1319;
assign nor1320 = !(nand0996|nand0993|nand0974|nand0980); 
assign invert0322 = nor1320;
assign nor1321 = !(nand0996|nand0993|nand0980|nand0975); 
assign invert0323 = nor1321;
assign nor1322 = !(nand0996|nand0993|nand0980|nand0976); 
assign invert0324 = nor1322;
assign nor1323 = !(nand0977|nand0996|nand0993|nand0980); 
assign invert0325 = nor1323;
assign nor1324 = !(nand0996|nand0993|nand0980|nand0978); 
assign invert0326 = nor1324;
assign nor1325 = !(nand0996|nand0993|nand0979|nand0980); 
assign invert0327 = nor1325;
assign nor1326 = !(nand0996|nand0993|nand0972|nand0981); 
assign invert0328 = nor1326;
assign nor1327 = !(nand0996|nand0993|nand0973|nand0981); 
assign invert0329 = nor1327;
assign nor1328 = !(nand0996|nand0993|nand0974|nand0981); 
assign invert0330 = nor1328;
assign nor1329 = !(nand0996|nand0993|nand0975|nand0981); 
assign invert0331 = nor1329;
assign nor1330 = !(nand0996|nand0993|nand0976|nand0981); 
assign invert0332 = nor1330;
assign nor1331 = !(nand0977|nand0996|nand0993|nand0981); 
assign invert0333 = nor1331;
assign nor1332 = !(nand0996|nand0993|nand0978|nand0981); 
assign invert0334 = nor1332;
assign nor1333 = !(nand0996|nand0993|nand0979|nand0981); 
assign invert0335 = nor1333;
assign nor1334 = !(nand0996|nand0993|nand0982|nand0972); 
assign invert0336 = nor1334;
assign nor1335 = !(nand0996|nand0993|nand0973|nand0982); 
assign invert0337 = nor1335;
assign nor1336 = !(nand0996|nand0993|nand0974|nand0982); 
assign invert0338 = nor1336;
assign nor1337 = !(nand0996|nand0993|nand0982|nand0975); 
assign invert0339 = nor1337;
assign nor1338 = !(nand0996|nand0993|nand0976|nand0982); 
assign invert0340 = nor1338;
assign nor1339 = !(nand0977|nand0996|nand0993|nand0982); 
assign invert0341 = nor1339;
assign nor1340 = !(nand0996|nand0993|nand0982|nand0978); 
assign invert0342 = nor1340;
assign nor1341 = !(nand0996|nand0993|nand0979|nand0982); 
assign invert0343 = nor1341;
assign nor1342 = !(nand0996|nand0993|nand0983|nand0972); 
assign invert0344 = nor1342;
assign nor1343 = !(nand0996|nand0993|nand0983|nand0973); 
assign invert0345 = nor1343;
assign nor1344 = !(nand0996|nand0993|nand0974|nand0983); 
assign invert0346 = nor1344;
assign nor1345 = !(nand0996|nand0993|nand0983|nand0975); 
assign invert0347 = nor1345;
assign nor1346 = !(nand0996|nand0993|nand0983|nand0976); 
assign invert0348 = nor1346;
assign nor1347 = !(nand0977|nand0996|nand0993|nand0983); 
assign invert0349 = nor1347;
assign nor1348 = !(nand0996|nand0993|nand0983|nand0978); 
assign invert0350 = nor1348;
assign nor1349 = !(nand0996|nand0993|nand0983|nand0979); 
assign invert0351 = nor1349;
assign nor1350 = !(nand0996|nand0993|nand0972|nand0984); 
assign invert0352 = nor1350;
assign nor1351 = !(nand0996|nand0993|nand0973|nand0984); 
assign invert0353 = nor1351;
assign nor1352 = !(nand0996|nand0993|nand0974|nand0984); 
assign invert0354 = nor1352;
assign nor1353 = !(nand0996|nand0993|nand0975|nand0984); 
assign invert0355 = nor1353;
assign nor1354 = !(nand0996|nand0993|nand0976|nand0984); 
assign invert0356 = nor1354;
assign nor1355 = !(nand0977|nand0996|nand0993|nand0984); 
assign invert0357 = nor1355;
assign nor1356 = !(nand0996|nand0993|nand0978|nand0984); 
assign invert0358 = nor1356;
assign nor1357 = !(nand0996|nand0993|nand0979|nand0984); 
assign invert0359 = nor1357;
assign nor1358 = !(nand0996|nand0993|nand0985|nand0972); 
assign invert0360 = nor1358;
assign nor1359 = !(nand0996|nand0993|nand0973|nand0985); 
assign invert0361 = nor1359;
assign nor1360 = !(nand0996|nand0993|nand0974|nand0985); 
assign invert0362 = nor1360;
assign nor1361 = !(nand0996|nand0993|nand0985|nand0975); 
assign invert0363 = nor1361;
assign nor1362 = !(nand0996|nand0993|nand0976|nand0985); 
assign invert0364 = nor1362;
assign nor1363 = !(nand0977|nand0996|nand0993|nand0985); 
assign invert0365 = nor1363;
assign nor1364 = !(nand0996|nand0993|nand0985|nand0978); 
assign invert0366 = nor1364;
assign nor1365 = !(nand0996|nand0993|nand0979|nand0985); 
assign invert0367 = nor1365;
assign nor1366 = !(nand0996|nand0986|nand0993|nand0972); 
assign invert0368 = nor1366;
assign nor1367 = !(nand0996|nand0986|nand0993|nand0973); 
assign invert0369 = nor1367;
assign nor1368 = !(nand0996|nand0986|nand0993|nand0974); 
assign invert0370 = nor1368;
assign nor1369 = !(nand0996|nand0986|nand0993|nand0975); 
assign invert0371 = nor1369;
assign nor1370 = !(nand0996|nand0986|nand0993|nand0976); 
assign invert0372 = nor1370;
assign nor1371 = !(nand0977|nand0996|nand0986|nand0993); 
assign invert0373 = nor1371;
assign nor1372 = !(nand0996|nand0986|nand0993|nand0978); 
assign invert0374 = nor1372;
assign nor1373 = !(nand0996|nand0986|nand0993|nand0979); 
assign invert0375 = nor1373;
assign nor1374 = !(nand0996|nand0993|nand0987|nand0972); 
assign invert0376 = nor1374;
assign nor1375 = !(nand0996|nand0993|nand0973|nand0987); 
assign invert0377 = nor1375;
assign nor1376 = !(nand0996|nand0993|nand0974|nand0987); 
assign invert0378 = nor1376;
assign nor1377 = !(nand0996|nand0993|nand0987|nand0975); 
assign invert0379 = nor1377;
assign nor1378 = !(nand0996|nand0993|nand0976|nand0987); 
assign invert0380 = nor1378;
assign nor1379 = !(nand0977|nand0996|nand0993|nand0987); 
assign invert0381 = nor1379;
assign nor1380 = !(nand0996|nand0993|nand0978|nand0987); 
assign invert0382 = nor1380;
assign nor1381 = !(nand0996|nand0993|nand0979|nand0987); 
assign invert0383 = nor1381;
assign nor1382 = !(nand0996|nand0980|nand0994|nand0972); 
assign invert0384 = nor1382;
assign nor1383 = !(nand0996|nand0980|nand0973|nand0994); 
assign invert0385 = nor1383;
assign nor1384 = !(nand0996|nand0974|nand0980|nand0994); 
assign invert0386 = nor1384;
assign nor1385 = !(nand0996|nand0980|nand0975|nand0994); 
assign invert0387 = nor1385;
assign nor1386 = !(nand0996|nand0980|nand0976|nand0994); 
assign invert0388 = nor1386;
assign nor1387 = !(nand0977|nand0996|nand0980|nand0994); 
assign invert0389 = nor1387;
assign nor1388 = !(nand0996|nand0980|nand0978|nand0994); 
assign invert0390 = nor1388;
assign nor1389 = !(nand0996|nand0979|nand0980|nand0994); 
assign invert0391 = nor1389;
assign nor1390 = !(nand0996|nand0994|nand0972|nand0981); 
assign invert0392 = nor1390;
assign nor1391 = !(nand0996|nand0973|nand0994|nand0981); 
assign invert0393 = nor1391;
assign nor1392 = !(nand0996|nand0974|nand0994|nand0981); 
assign invert0394 = nor1392;
assign nor1393 = !(nand0996|nand0975|nand0994|nand0981); 
assign invert0395 = nor1393;
assign nor1394 = !(nand0996|nand0976|nand0994|nand0981); 
assign invert0396 = nor1394;
assign nor1395 = !(nand0977|nand0996|nand0994|nand0981); 
assign invert0397 = nor1395;
assign nor1396 = !(nand0996|nand0978|nand0994|nand0981); 
assign invert0398 = nor1396;
assign nor1397 = !(nand0996|nand0979|nand0994|nand0981); 
assign invert0399 = nor1397;
assign nor1398 = !(nand0996|nand0982|nand0994|nand0972); 
assign invert0400 = nor1398;
assign nor1399 = !(nand0996|nand0973|nand0982|nand0994); 
assign invert0401 = nor1399;
assign nor1400 = !(nand0996|nand0974|nand0982|nand0994); 
assign invert0402 = nor1400;
assign nor1401 = !(nand0996|nand0982|nand0975|nand0994); 
assign invert0403 = nor1401;
assign nor1402 = !(nand0996|nand0976|nand0982|nand0994); 
assign invert0404 = nor1402;
assign nor1403 = !(nand0977|nand0996|nand0982|nand0994); 
assign invert0405 = nor1403;
assign nor1404 = !(nand0996|nand0982|nand0978|nand0994); 
assign invert0406 = nor1404;
assign nor1405 = !(nand0996|nand0979|nand0982|nand0994); 
assign invert0407 = nor1405;
assign nor1406 = !(nand0996|nand0983|nand0994|nand0972); 
assign invert0408 = nor1406;
assign nor1407 = !(nand0996|nand0983|nand0973|nand0994); 
assign invert0409 = nor1407;
assign nor1408 = !(nand0996|nand0974|nand0983|nand0994); 
assign invert0410 = nor1408;
assign nor1409 = !(nand0996|nand0983|nand0975|nand0994); 
assign invert0411 = nor1409;
assign nor1410 = !(nand0996|nand0983|nand0976|nand0994); 
assign invert0412 = nor1410;
assign nor1411 = !(nand0977|nand0996|nand0983|nand0994); 
assign invert0413 = nor1411;
assign nor1412 = !(nand0996|nand0983|nand0978|nand0994); 
assign invert0414 = nor1412;
assign nor1413 = !(nand0996|nand0983|nand0979|nand0994); 
assign invert0415 = nor1413;
assign nor1414 = !(nand0996|nand0994|nand0972|nand0984); 
assign invert0416 = nor1414;
assign nor1415 = !(nand0996|nand0973|nand0994|nand0984); 
assign invert0417 = nor1415;
assign nor1416 = !(nand0996|nand0974|nand0994|nand0984); 
assign invert0418 = nor1416;
assign nor1417 = !(nand0996|nand0975|nand0994|nand0984); 
assign invert0419 = nor1417;
assign nor1418 = !(nand0996|nand0976|nand0994|nand0984); 
assign invert0420 = nor1418;
assign nor1419 = !(nand0977|nand0996|nand0994|nand0984); 
assign invert0421 = nor1419;
assign nor1420 = !(nand0996|nand0978|nand0994|nand0984); 
assign invert0422 = nor1420;
assign nor1421 = !(nand0996|nand0979|nand0994|nand0984); 
assign invert0423 = nor1421;
assign nor1422 = !(nand0996|nand0985|nand0994|nand0972); 
assign invert0424 = nor1422;
assign nor1423 = !(nand0996|nand0973|nand0985|nand0994); 
assign invert0425 = nor1423;
assign nor1424 = !(nand0996|nand0974|nand0985|nand0994); 
assign invert0426 = nor1424;
assign nor1425 = !(nand0996|nand0985|nand0975|nand0994); 
assign invert0427 = nor1425;
assign nor1426 = !(nand0996|nand0976|nand0985|nand0994); 
assign invert0428 = nor1426;
assign nor1427 = !(nand0977|nand0996|nand0985|nand0994); 
assign invert0429 = nor1427;
assign nor1428 = !(nand0996|nand0985|nand0978|nand0994); 
assign invert0430 = nor1428;
assign nor1429 = !(nand0996|nand0979|nand0985|nand0994); 
assign invert0431 = nor1429;
assign nor1430 = !(nand0996|nand0986|nand0994|nand0972); 
assign invert0432 = nor1430;
assign nor1431 = !(nand0996|nand0986|nand0973|nand0994); 
assign invert0433 = nor1431;
assign nor1432 = !(nand0996|nand0986|nand0974|nand0994); 
assign invert0434 = nor1432;
assign nor1433 = !(nand0996|nand0986|nand0975|nand0994); 
assign invert0435 = nor1433;
assign nor1434 = !(nand0996|nand0986|nand0976|nand0994); 
assign invert0436 = nor1434;
assign nor1435 = !(nand0977|nand0996|nand0986|nand0994); 
assign invert0437 = nor1435;
assign nor1436 = !(nand0996|nand0986|nand0978|nand0994); 
assign invert0438 = nor1436;
assign nor1437 = !(nand0996|nand0986|nand0979|nand0994); 
assign invert0439 = nor1437;
assign nor1438 = !(nand0996|nand0987|nand0994|nand0972); 
assign invert0440 = nor1438;
assign nor1439 = !(nand0996|nand0973|nand0987|nand0994); 
assign invert0441 = nor1439;
assign nor1440 = !(nand0996|nand0974|nand0987|nand0994); 
assign invert0442 = nor1440;
assign nor1441 = !(nand0996|nand0987|nand0975|nand0994); 
assign invert0443 = nor1441;
assign nor1442 = !(nand0996|nand0976|nand0987|nand0994); 
assign invert0444 = nor1442;
assign nor1443 = !(nand0977|nand0996|nand0987|nand0994); 
assign invert0445 = nor1443;
assign nor1444 = !(nand0996|nand0978|nand0987|nand0994); 
assign invert0446 = nor1444;
assign nor1445 = !(nand0996|nand0979|nand0987|nand0994); 
assign invert0447 = nor1445;
assign nor1446 = !(nand0996|nand0980|nand0995|nand0972); 
assign invert0448 = nor1446;
assign nor1447 = !(nand0996|nand0980|nand0995|nand0973); 
assign invert0449 = nor1447;
assign nor1448 = !(nand0996|nand0974|nand0980|nand0995); 
assign invert0450 = nor1448;
assign nor1449 = !(nand0996|nand0980|nand0995|nand0975); 
assign invert0451 = nor1449;
assign nor1450 = !(nand0996|nand0980|nand0976|nand0995); 
assign invert0452 = nor1450;
assign nor1451 = !(nand0977|nand0996|nand0980|nand0995); 
assign invert0453 = nor1451;
assign nor1452 = !(nand0996|nand0980|nand0995|nand0978); 
assign invert0454 = nor1452;
assign nor1453 = !(nand0996|nand0979|nand0980|nand0995); 
assign invert0455 = nor1453;
assign nor1454 = !(nand0996|nand0995|nand0972|nand0981); 
assign invert0456 = nor1454;
assign nor1455 = !(nand0996|nand0995|nand0973|nand0981); 
assign invert0457 = nor1455;
assign nor1456 = !(nand0996|nand0974|nand0995|nand0981); 
assign invert0458 = nor1456;
assign nor1457 = !(nand0996|nand0995|nand0975|nand0981); 
assign invert0459 = nor1457;
assign nor1458 = !(nand0996|nand0976|nand0995|nand0981); 
assign invert0460 = nor1458;
assign nor1459 = !(nand0977|nand0996|nand0995|nand0981); 
assign invert0461 = nor1459;
assign nor1460 = !(nand0996|nand0995|nand0978|nand0981); 
assign invert0462 = nor1460;
assign nor1461 = !(nand0996|nand0979|nand0995|nand0981); 
assign invert0463 = nor1461;
assign nor1462 = !(nand0996|nand0995|nand0982|nand0972); 
assign invert0464 = nor1462;
assign nor1463 = !(nand0996|nand0995|nand0973|nand0982); 
assign invert0465 = nor1463;
assign nor1464 = !(nand0996|nand0974|nand0995|nand0982); 
assign invert0466 = nor1464;
assign nor1465 = !(nand0996|nand0995|nand0982|nand0975); 
assign invert0467 = nor1465;
assign nor1466 = !(nand0996|nand0976|nand0995|nand0982); 
assign invert0468 = nor1466;
assign nor1467 = !(nand0977|nand0996|nand0995|nand0982); 
assign invert0469 = nor1467;
assign nor1468 = !(nand0996|nand0995|nand0982|nand0978); 
assign invert0470 = nor1468;
assign nor1469 = !(nand0996|nand0979|nand0995|nand0982); 
assign invert0471 = nor1469;
assign nor1470 = !(nand0996|nand0983|nand0995|nand0972); 
assign invert0472 = nor1470;
assign nor1471 = !(nand0996|nand0983|nand0995|nand0973); 
assign invert0473 = nor1471;
assign nor1472 = !(nand0996|nand0974|nand0983|nand0995); 
assign invert0474 = nor1472;
assign nor1473 = !(nand0996|nand0983|nand0995|nand0975); 
assign invert0475 = nor1473;
assign nor1474 = !(nand0996|nand0983|nand0976|nand0995); 
assign invert0476 = nor1474;
assign nor1475 = !(nand0977|nand0996|nand0983|nand0995); 
assign invert0477 = nor1475;
assign nor1476 = !(nand0996|nand0983|nand0995|nand0978); 
assign invert0478 = nor1476;
assign nor1477 = !(nand0996|nand0983|nand0979|nand0995); 
assign invert0479 = nor1477;
assign nor1478 = !(nand0996|nand0995|nand0972|nand0984); 
assign invert0480 = nor1478;
assign nor1479 = !(nand0996|nand0995|nand0973|nand0984); 
assign invert0481 = nor1479;
assign nor1480 = !(nand0996|nand0974|nand0995|nand0984); 
assign invert0482 = nor1480;
assign nor1481 = !(nand0996|nand0995|nand0975|nand0984); 
assign invert0483 = nor1481;
assign nor1482 = !(nand0996|nand0976|nand0995|nand0984); 
assign invert0484 = nor1482;
assign nor1483 = !(nand0977|nand0996|nand0995|nand0984); 
assign invert0485 = nor1483;
assign nor1484 = !(nand0996|nand0995|nand0978|nand0984); 
assign invert0486 = nor1484;
assign nor1485 = !(nand0996|nand0979|nand0995|nand0984); 
assign invert0487 = nor1485;
assign nor1486 = !(nand0996|nand0995|nand0985|nand0972); 
assign invert0488 = nor1486;
assign nor1487 = !(nand0996|nand0995|nand0973|nand0985); 
assign invert0489 = nor1487;
assign nor1488 = !(nand0996|nand0974|nand0995|nand0985); 
assign invert0490 = nor1488;
assign nor1489 = !(nand0996|nand0995|nand0985|nand0975); 
assign invert0491 = nor1489;
assign nor1490 = !(nand0996|nand0976|nand0995|nand0985); 
assign invert0492 = nor1490;
assign nor1491 = !(nand0977|nand0996|nand0995|nand0985); 
assign invert0493 = nor1491;
assign nor1492 = !(nand0996|nand0995|nand0985|nand0978); 
assign invert0494 = nor1492;
assign nor1493 = !(nand0996|nand0979|nand0995|nand0985); 
assign invert0495 = nor1493;
assign nor1494 = !(nand0996|nand0986|nand0995|nand0972); 
assign invert0496 = nor1494;
assign nor1495 = !(nand0996|nand0986|nand0995|nand0973); 
assign invert0497 = nor1495;
assign nor1496 = !(nand0996|nand0986|nand0974|nand0995); 
assign invert0498 = nor1496;
assign nor1497 = !(nand0996|nand0986|nand0995|nand0975); 
assign invert0499 = nor1497;
assign nor1498 = !(nand0996|nand0986|nand0976|nand0995); 
assign invert0500 = nor1498;
assign nor1499 = !(nand0977|nand0996|nand0986|nand0995); 
assign invert0501 = nor1499;
assign nor1500 = !(nand0996|nand0986|nand0995|nand0978); 
assign invert0502 = nor1500;
assign nor1501 = !(nand0996|nand0986|nand0979|nand0995); 
assign invert0503 = nor1501;
assign nor1502 = !(nand0996|nand0995|nand0987|nand0972); 
assign invert0504 = nor1502;
assign nor1503 = !(nand0996|nand0995|nand0973|nand0987); 
assign invert0505 = nor1503;
assign nor1504 = !(nand0996|nand0974|nand0995|nand0987); 
assign invert0506 = nor1504;
assign nor1505 = !(nand0996|nand0995|nand0987|nand0975); 
assign invert0507 = nor1505;
assign nor1506 = !(nand0996|nand0976|nand0995|nand0987); 
assign invert0508 = nor1506;
assign nor1507 = !(nand0977|nand0996|nand0995|nand0987); 
assign invert0509 = nor1507;
assign nor1508 = !(nand0996|nand0995|nand0978|nand0987); 
assign invert0510 = nor1508;
assign nor1509 = !(nand0996|nand0979|nand0995|nand0987); 
assign invert0511 = nor1509;
assign nor1510 = !(nand0980|nand0988|nand0997|nand0972); 
assign invert0512 = nor1510;
assign nor1511 = !(nand0980|nand0988|nand0973|nand0997); 
assign invert0513 = nor1511;
assign nor1512 = !(nand0974|nand0980|nand0988|nand0997); 
assign invert0514 = nor1512;
assign nor1513 = !(nand0980|nand0988|nand0997|nand0975); 
assign invert0515 = nor1513;
assign nor1514 = !(nand0980|nand0988|nand0976|nand0997); 
assign invert0516 = nor1514;
assign nor1515 = !(nand0977|nand0980|nand0988|nand0997); 
assign invert0517 = nor1515;
assign nor1516 = !(nand0980|nand0988|nand0997|nand0978); 
assign invert0518 = nor1516;
assign nor1517 = !(nand0979|nand0980|nand0988|nand0997); 
assign invert0519 = nor1517;
assign nor1518 = !(nand0988|nand0997|nand0972|nand0981); 
assign invert0520 = nor1518;
assign nor1519 = !(nand0988|nand0973|nand0997|nand0981); 
assign invert0521 = nor1519;
assign nor1520 = !(nand0974|nand0988|nand0997|nand0981); 
assign invert0522 = nor1520;
assign nor1521 = !(nand0988|nand0997|nand0975|nand0981); 
assign invert0523 = nor1521;
assign nor1522 = !(nand0988|nand0976|nand0997|nand0981); 
assign invert0524 = nor1522;
assign nor1523 = !(nand0977|nand0988|nand0997|nand0981); 
assign invert0525 = nor1523;
assign nor1524 = !(nand0988|nand0997|nand0978|nand0981); 
assign invert0526 = nor1524;
assign nor1525 = !(nand0979|nand0988|nand0997|nand0981); 
assign invert0527 = nor1525;
assign nor1526 = !(nand0988|nand0982|nand0997|nand0972); 
assign invert0528 = nor1526;
assign nor1527 = !(nand0988|nand0973|nand0982|nand0997); 
assign invert0529 = nor1527;
assign nor1528 = !(nand0974|nand0988|nand0982|nand0997); 
assign invert0530 = nor1528;
assign nor1529 = !(nand0988|nand0982|nand0997|nand0975); 
assign invert0531 = nor1529;
assign nor1530 = !(nand0988|nand0976|nand0982|nand0997); 
assign invert0532 = nor1530;
assign nor1531 = !(nand0977|nand0988|nand0982|nand0997); 
assign invert0533 = nor1531;
assign nor1532 = !(nand0988|nand0982|nand0997|nand0978); 
assign invert0534 = nor1532;
assign nor1533 = !(nand0979|nand0988|nand0982|nand0997); 
assign invert0535 = nor1533;
assign nor1534 = !(nand0983|nand0988|nand0997|nand0972); 
assign invert0536 = nor1534;
assign nor1535 = !(nand0983|nand0988|nand0973|nand0997); 
assign invert0537 = nor1535;
assign nor1536 = !(nand0974|nand0983|nand0988|nand0997); 
assign invert0538 = nor1536;
assign nor1537 = !(nand0983|nand0988|nand0997|nand0975); 
assign invert0539 = nor1537;
assign nor1538 = !(nand0983|nand0988|nand0976|nand0997); 
assign invert0540 = nor1538;
assign nor1539 = !(nand0977|nand0983|nand0988|nand0997); 
assign invert0541 = nor1539;
assign nor1540 = !(nand0983|nand0988|nand0997|nand0978); 
assign invert0542 = nor1540;
assign nor1541 = !(nand0983|nand0979|nand0988|nand0997); 
assign invert0543 = nor1541;
assign nor1542 = !(nand0988|nand0997|nand0972|nand0984); 
assign invert0544 = nor1542;
assign nor1543 = !(nand0988|nand0973|nand0997|nand0984); 
assign invert0545 = nor1543;
assign nor1544 = !(nand0974|nand0988|nand0997|nand0984); 
assign invert0546 = nor1544;
assign nor1545 = !(nand0988|nand0997|nand0975|nand0984); 
assign invert0547 = nor1545;
assign nor1546 = !(nand0988|nand0976|nand0997|nand0984); 
assign invert0548 = nor1546;
assign nor1547 = !(nand0977|nand0988|nand0997|nand0984); 
assign invert0549 = nor1547;
assign nor1548 = !(nand0988|nand0997|nand0978|nand0984); 
assign invert0550 = nor1548;
assign nor1549 = !(nand0979|nand0988|nand0997|nand0984); 
assign invert0551 = nor1549;
assign nor1550 = !(nand0988|nand0985|nand0997|nand0972); 
assign invert0552 = nor1550;
assign nor1551 = !(nand0988|nand0973|nand0985|nand0997); 
assign invert0553 = nor1551;
assign nor1552 = !(nand0974|nand0988|nand0985|nand0997); 
assign invert0554 = nor1552;
assign nor1553 = !(nand0988|nand0985|nand0997|nand0975); 
assign invert0555 = nor1553;
assign nor1554 = !(nand0988|nand0976|nand0985|nand0997); 
assign invert0556 = nor1554;
assign nor1555 = !(nand0977|nand0988|nand0985|nand0997); 
assign invert0557 = nor1555;
assign nor1556 = !(nand0988|nand0985|nand0997|nand0978); 
assign invert0558 = nor1556;
assign nor1557 = !(nand0979|nand0988|nand0985|nand0997); 
assign invert0559 = nor1557;
assign nor1558 = !(nand0986|nand0988|nand0997|nand0972); 
assign invert0560 = nor1558;
assign nor1559 = !(nand0986|nand0988|nand0973|nand0997); 
assign invert0561 = nor1559;
assign nor1560 = !(nand0986|nand0974|nand0988|nand0997); 
assign invert0562 = nor1560;
assign nor1561 = !(nand0986|nand0988|nand0997|nand0975); 
assign invert0563 = nor1561;
assign nor1562 = !(nand0986|nand0988|nand0976|nand0997); 
assign invert0564 = nor1562;
assign nor1563 = !(nand0977|nand0986|nand0988|nand0997); 
assign invert0565 = nor1563;
assign nor1564 = !(nand0986|nand0988|nand0997|nand0978); 
assign invert0566 = nor1564;
assign nor1565 = !(nand0986|nand0979|nand0988|nand0997); 
assign invert0567 = nor1565;
assign nor1566 = !(nand0988|nand0997|nand0987|nand0972); 
assign invert0568 = nor1566;
assign nor1567 = !(nand0988|nand0973|nand0997|nand0987); 
assign invert0569 = nor1567;
assign nor1568 = !(nand0974|nand0988|nand0997|nand0987); 
assign invert0570 = nor1568;
assign nor1569 = !(nand0988|nand0997|nand0987|nand0975); 
assign invert0571 = nor1569;
assign nor1570 = !(nand0988|nand0976|nand0997|nand0987); 
assign invert0572 = nor1570;
assign nor1571 = !(nand0977|nand0988|nand0997|nand0987); 
assign invert0573 = nor1571;
assign nor1572 = !(nand0988|nand0997|nand0978|nand0987); 
assign invert0574 = nor1572;
assign nor1573 = !(nand0979|nand0988|nand0997|nand0987); 
assign invert0575 = nor1573;
assign nor1574 = !(nand0989|nand0980|nand0997|nand0972); 
assign invert0576 = nor1574;
assign nor1575 = !(nand0989|nand0980|nand0973|nand0997); 
assign invert0577 = nor1575;
assign nor1576 = !(nand0989|nand0974|nand0980|nand0997); 
assign invert0578 = nor1576;
assign nor1577 = !(nand0989|nand0980|nand0997|nand0975); 
assign invert0579 = nor1577;
assign nor1578 = !(nand0989|nand0980|nand0976|nand0997); 
assign invert0580 = nor1578;
assign nor1579 = !(nand0989|nand0977|nand0980|nand0997); 
assign invert0581 = nor1579;
assign nor1580 = !(nand0989|nand0980|nand0997|nand0978); 
assign invert0582 = nor1580;
assign nor1581 = !(nand0989|nand0979|nand0980|nand0997); 
assign invert0583 = nor1581;
assign nor1582 = !(nand0989|nand0997|nand0972|nand0981); 
assign invert0584 = nor1582;
assign nor1583 = !(nand0989|nand0973|nand0997|nand0981); 
assign invert0585 = nor1583;
assign nor1584 = !(nand0989|nand0974|nand0997|nand0981); 
assign invert0586 = nor1584;
assign nor1585 = !(nand0989|nand0997|nand0975|nand0981); 
assign invert0587 = nor1585;
assign nor1586 = !(nand0989|nand0976|nand0997|nand0981); 
assign invert0588 = nor1586;
assign nor1587 = !(nand0989|nand0977|nand0997|nand0981); 
assign invert0589 = nor1587;
assign nor1588 = !(nand0989|nand0997|nand0978|nand0981); 
assign invert0590 = nor1588;
assign nor1589 = !(nand0989|nand0979|nand0997|nand0981); 
assign invert0591 = nor1589;
assign nor1590 = !(nand0989|nand0982|nand0997|nand0972); 
assign invert0592 = nor1590;
assign nor1591 = !(nand0989|nand0973|nand0982|nand0997); 
assign invert0593 = nor1591;
assign nor1592 = !(nand0989|nand0974|nand0982|nand0997); 
assign invert0594 = nor1592;
assign nor1593 = !(nand0989|nand0982|nand0997|nand0975); 
assign invert0595 = nor1593;
assign nor1594 = !(nand0989|nand0976|nand0982|nand0997); 
assign invert0596 = nor1594;
assign nor1595 = !(nand0989|nand0977|nand0982|nand0997); 
assign invert0597 = nor1595;
assign nor1596 = !(nand0989|nand0982|nand0997|nand0978); 
assign invert0598 = nor1596;
assign nor1597 = !(nand0989|nand0979|nand0982|nand0997); 
assign invert0599 = nor1597;
assign nor1598 = !(nand0989|nand0983|nand0997|nand0972); 
assign invert0600 = nor1598;
assign nor1599 = !(nand0989|nand0983|nand0973|nand0997); 
assign invert0601 = nor1599;
assign nor1600 = !(nand0989|nand0974|nand0983|nand0997); 
assign invert0602 = nor1600;
assign nor1601 = !(nand0989|nand0983|nand0997|nand0975); 
assign invert0603 = nor1601;
assign nor1602 = !(nand0989|nand0983|nand0976|nand0997); 
assign invert0604 = nor1602;
assign nor1603 = !(nand0989|nand0977|nand0983|nand0997); 
assign invert0605 = nor1603;
assign nor1604 = !(nand0989|nand0983|nand0997|nand0978); 
assign invert0606 = nor1604;
assign nor1605 = !(nand0989|nand0983|nand0979|nand0997); 
assign invert0607 = nor1605;
assign nor1606 = !(nand0989|nand0997|nand0972|nand0984); 
assign invert0608 = nor1606;
assign nor1607 = !(nand0989|nand0973|nand0997|nand0984); 
assign invert0609 = nor1607;
assign nor1608 = !(nand0989|nand0974|nand0997|nand0984); 
assign invert0610 = nor1608;
assign nor1609 = !(nand0989|nand0997|nand0975|nand0984); 
assign invert0611 = nor1609;
assign nor1610 = !(nand0989|nand0976|nand0997|nand0984); 
assign invert0612 = nor1610;
assign nor1611 = !(nand0989|nand0977|nand0997|nand0984); 
assign invert0613 = nor1611;
assign nor1612 = !(nand0989|nand0997|nand0978|nand0984); 
assign invert0614 = nor1612;
assign nor1613 = !(nand0989|nand0979|nand0997|nand0984); 
assign invert0615 = nor1613;
assign nor1614 = !(nand0989|nand0985|nand0997|nand0972); 
assign invert0616 = nor1614;
assign nor1615 = !(nand0989|nand0973|nand0985|nand0997); 
assign invert0617 = nor1615;
assign nor1616 = !(nand0989|nand0974|nand0985|nand0997); 
assign invert0618 = nor1616;
assign nor1617 = !(nand0989|nand0985|nand0997|nand0975); 
assign invert0619 = nor1617;
assign nor1618 = !(nand0989|nand0976|nand0985|nand0997); 
assign invert0620 = nor1618;
assign nor1619 = !(nand0989|nand0977|nand0985|nand0997); 
assign invert0621 = nor1619;
assign nor1620 = !(nand0989|nand0985|nand0997|nand0978); 
assign invert0622 = nor1620;
assign nor1621 = !(nand0989|nand0979|nand0985|nand0997); 
assign invert0623 = nor1621;
assign nor1622 = !(nand0989|nand0986|nand0997|nand0972); 
assign invert0624 = nor1622;
assign nor1623 = !(nand0989|nand0986|nand0973|nand0997); 
assign invert0625 = nor1623;
assign nor1624 = !(nand0989|nand0986|nand0974|nand0997); 
assign invert0626 = nor1624;
assign nor1625 = !(nand0989|nand0986|nand0997|nand0975); 
assign invert0627 = nor1625;
assign nor1626 = !(nand0989|nand0986|nand0976|nand0997); 
assign invert0628 = nor1626;
assign nor1627 = !(nand0989|nand0977|nand0986|nand0997); 
assign invert0629 = nor1627;
assign nor1628 = !(nand0989|nand0986|nand0997|nand0978); 
assign invert0630 = nor1628;
assign nor1629 = !(nand0989|nand0986|nand0979|nand0997); 
assign invert0631 = nor1629;
assign nor1630 = !(nand0989|nand0997|nand0987|nand0972); 
assign invert0632 = nor1630;
assign nor1631 = !(nand0989|nand0973|nand0997|nand0987); 
assign invert0633 = nor1631;
assign nor1632 = !(nand0989|nand0974|nand0997|nand0987); 
assign invert0634 = nor1632;
assign nor1633 = !(nand0989|nand0997|nand0987|nand0975); 
assign invert0635 = nor1633;
assign nor1634 = !(nand0989|nand0976|nand0997|nand0987); 
assign invert0636 = nor1634;
assign nor1635 = !(nand0989|nand0977|nand0997|nand0987); 
assign invert0637 = nor1635;
assign nor1636 = !(nand0989|nand0997|nand0978|nand0987); 
assign invert0638 = nor1636;
assign nor1637 = !(nand0989|nand0979|nand0997|nand0987); 
assign invert0639 = nor1637;
assign nor1638 = !(nand0990|nand0980|nand0997|nand0972); 
assign invert0640 = nor1638;
assign nor1639 = !(nand0990|nand0980|nand0973|nand0997); 
assign invert0641 = nor1639;
assign nor1640 = !(nand0974|nand0990|nand0980|nand0997); 
assign invert0642 = nor1640;
assign nor1641 = !(nand0990|nand0980|nand0997|nand0975); 
assign invert0643 = nor1641;
assign nor1642 = !(nand0990|nand0980|nand0976|nand0997); 
assign invert0644 = nor1642;
assign nor1643 = !(nand0977|nand0990|nand0980|nand0997); 
assign invert0645 = nor1643;
assign nor1644 = !(nand0990|nand0980|nand0997|nand0978); 
assign invert0646 = nor1644;
assign nor1645 = !(nand0990|nand0979|nand0980|nand0997); 
assign invert0647 = nor1645;
assign nor1646 = !(nand0990|nand0997|nand0972|nand0981); 
assign invert0648 = nor1646;
assign nor1647 = !(nand0990|nand0973|nand0997|nand0981); 
assign invert0649 = nor1647;
assign nor1648 = !(nand0974|nand0990|nand0997|nand0981); 
assign invert0650 = nor1648;
assign nor1649 = !(nand0990|nand0997|nand0975|nand0981); 
assign invert0651 = nor1649;
assign nor1650 = !(nand0990|nand0976|nand0997|nand0981); 
assign invert0652 = nor1650;
assign nor1651 = !(nand0977|nand0990|nand0997|nand0981); 
assign invert0653 = nor1651;
assign nor1652 = !(nand0990|nand0997|nand0978|nand0981); 
assign invert0654 = nor1652;
assign nor1653 = !(nand0990|nand0979|nand0997|nand0981); 
assign invert0655 = nor1653;
assign nor1654 = !(nand0990|nand0982|nand0997|nand0972); 
assign invert0656 = nor1654;
assign nor1655 = !(nand0990|nand0973|nand0982|nand0997); 
assign invert0657 = nor1655;
assign nor1656 = !(nand0974|nand0990|nand0982|nand0997); 
assign invert0658 = nor1656;
assign nor1657 = !(nand0990|nand0982|nand0997|nand0975); 
assign invert0659 = nor1657;
assign nor1658 = !(nand0990|nand0976|nand0982|nand0997); 
assign invert0660 = nor1658;
assign nor1659 = !(nand0977|nand0990|nand0982|nand0997); 
assign invert0661 = nor1659;
assign nor1660 = !(nand0990|nand0982|nand0997|nand0978); 
assign invert0662 = nor1660;
assign nor1661 = !(nand0990|nand0979|nand0982|nand0997); 
assign invert0663 = nor1661;
assign nor1662 = !(nand0983|nand0990|nand0997|nand0972); 
assign invert0664 = nor1662;
assign nor1663 = !(nand0983|nand0990|nand0973|nand0997); 
assign invert0665 = nor1663;
assign nor1664 = !(nand0974|nand0983|nand0990|nand0997); 
assign invert0666 = nor1664;
assign nor1665 = !(nand0983|nand0990|nand0997|nand0975); 
assign invert0667 = nor1665;
assign nor1666 = !(nand0983|nand0990|nand0976|nand0997); 
assign invert0668 = nor1666;
assign nor1667 = !(nand0977|nand0983|nand0990|nand0997); 
assign invert0669 = nor1667;
assign nor1668 = !(nand0983|nand0990|nand0997|nand0978); 
assign invert0670 = nor1668;
assign nor1669 = !(nand0983|nand0990|nand0979|nand0997); 
assign invert0671 = nor1669;
assign nor1670 = !(nand0990|nand0997|nand0972|nand0984); 
assign invert0672 = nor1670;
assign nor1671 = !(nand0990|nand0973|nand0997|nand0984); 
assign invert0673 = nor1671;
assign nor1672 = !(nand0974|nand0990|nand0997|nand0984); 
assign invert0674 = nor1672;
assign nor1673 = !(nand0990|nand0997|nand0975|nand0984); 
assign invert0675 = nor1673;
assign nor1674 = !(nand0990|nand0976|nand0997|nand0984); 
assign invert0676 = nor1674;
assign nor1675 = !(nand0977|nand0990|nand0997|nand0984); 
assign invert0677 = nor1675;
assign nor1676 = !(nand0990|nand0997|nand0978|nand0984); 
assign invert0678 = nor1676;
assign nor1677 = !(nand0990|nand0979|nand0997|nand0984); 
assign invert0679 = nor1677;
assign nor1678 = !(nand0990|nand0985|nand0997|nand0972); 
assign invert0680 = nor1678;
assign nor1679 = !(nand0990|nand0973|nand0985|nand0997); 
assign invert0681 = nor1679;
assign nor1680 = !(nand0974|nand0990|nand0985|nand0997); 
assign invert0682 = nor1680;
assign nor1681 = !(nand0990|nand0985|nand0997|nand0975); 
assign invert0683 = nor1681;
assign nor1682 = !(nand0990|nand0976|nand0985|nand0997); 
assign invert0684 = nor1682;
assign nor1683 = !(nand0977|nand0990|nand0985|nand0997); 
assign invert0685 = nor1683;
assign nor1684 = !(nand0990|nand0985|nand0997|nand0978); 
assign invert0686 = nor1684;
assign nor1685 = !(nand0990|nand0979|nand0985|nand0997); 
assign invert0687 = nor1685;
assign nor1686 = !(nand0986|nand0990|nand0997|nand0972); 
assign invert0688 = nor1686;
assign nor1687 = !(nand0986|nand0990|nand0973|nand0997); 
assign invert0689 = nor1687;
assign nor1688 = !(nand0986|nand0974|nand0990|nand0997); 
assign invert0690 = nor1688;
assign nor1689 = !(nand0986|nand0990|nand0997|nand0975); 
assign invert0691 = nor1689;
assign nor1690 = !(nand0986|nand0990|nand0976|nand0997); 
assign invert0692 = nor1690;
assign nor1691 = !(nand0977|nand0986|nand0990|nand0997); 
assign invert0693 = nor1691;
assign nor1692 = !(nand0986|nand0990|nand0997|nand0978); 
assign invert0694 = nor1692;
assign nor1693 = !(nand0986|nand0990|nand0979|nand0997); 
assign invert0695 = nor1693;
assign nor1694 = !(nand0990|nand0997|nand0987|nand0972); 
assign invert0696 = nor1694;
assign nor1695 = !(nand0990|nand0973|nand0997|nand0987); 
assign invert0697 = nor1695;
assign nor1696 = !(nand0974|nand0990|nand0997|nand0987); 
assign invert0698 = nor1696;
assign nor1697 = !(nand0990|nand0997|nand0987|nand0975); 
assign invert0699 = nor1697;
assign nor1698 = !(nand0990|nand0976|nand0997|nand0987); 
assign invert0700 = nor1698;
assign nor1699 = !(nand0977|nand0990|nand0997|nand0987); 
assign invert0701 = nor1699;
assign nor1700 = !(nand0990|nand0997|nand0978|nand0987); 
assign invert0702 = nor1700;
assign nor1701 = !(nand0990|nand0979|nand0997|nand0987); 
assign invert0703 = nor1701;
assign nor1702 = !(nand0980|nand0997|nand0972|nand0991); 
assign invert0704 = nor1702;
assign nor1703 = !(nand0980|nand0973|nand0997|nand0991); 
assign invert0705 = nor1703;
assign nor1704 = !(nand0974|nand0980|nand0997|nand0991); 
assign invert0706 = nor1704;
assign nor1705 = !(nand0980|nand0997|nand0975|nand0991); 
assign invert0707 = nor1705;
assign nor1706 = !(nand0980|nand0976|nand0997|nand0991); 
assign invert0708 = nor1706;
assign nor1707 = !(nand0977|nand0980|nand0997|nand0991); 
assign invert0709 = nor1707;
assign nor1708 = !(nand0980|nand0997|nand0978|nand0991); 
assign invert0710 = nor1708;
assign nor1709 = !(nand0979|nand0980|nand0997|nand0991); 
assign invert0711 = nor1709;
assign nor1710 = !(nand0997|nand0972|nand0991|nand0981); 
assign invert0712 = nor1710;
assign nor1711 = !(nand0973|nand0997|nand0991|nand0981); 
assign invert0713 = nor1711;
assign nor1712 = !(nand0974|nand0997|nand0991|nand0981); 
assign invert0714 = nor1712;
assign nor1713 = !(nand0997|nand0975|nand0991|nand0981); 
assign invert0715 = nor1713;
assign nor1714 = !(nand0976|nand0997|nand0991|nand0981); 
assign invert0716 = nor1714;
assign nor1715 = !(nand0977|nand0997|nand0991|nand0981); 
assign invert0717 = nor1715;
assign nor1716 = !(nand0997|nand0978|nand0991|nand0981); 
assign invert0718 = nor1716;
assign nor1717 = !(nand0979|nand0997|nand0991|nand0981); 
assign invert0719 = nor1717;
assign nor1718 = !(nand0982|nand0997|nand0972|nand0991); 
assign invert0720 = nor1718;
assign nor1719 = !(nand0973|nand0982|nand0997|nand0991); 
assign invert0721 = nor1719;
assign nor1720 = !(nand0974|nand0982|nand0997|nand0991); 
assign invert0722 = nor1720;
assign nor1721 = !(nand0982|nand0997|nand0975|nand0991); 
assign invert0723 = nor1721;
assign nor1722 = !(nand0976|nand0982|nand0997|nand0991); 
assign invert0724 = nor1722;
assign nor1723 = !(nand0977|nand0982|nand0997|nand0991); 
assign invert0725 = nor1723;
assign nor1724 = !(nand0982|nand0997|nand0978|nand0991); 
assign invert0726 = nor1724;
assign nor1725 = !(nand0979|nand0982|nand0997|nand0991); 
assign invert0727 = nor1725;
assign nor1726 = !(nand0983|nand0997|nand0972|nand0991); 
assign invert0728 = nor1726;
assign nor1727 = !(nand0983|nand0973|nand0997|nand0991); 
assign invert0729 = nor1727;
assign nor1728 = !(nand0974|nand0983|nand0997|nand0991); 
assign invert0730 = nor1728;
assign nor1729 = !(nand0983|nand0997|nand0975|nand0991); 
assign invert0731 = nor1729;
assign nor1730 = !(nand0983|nand0976|nand0997|nand0991); 
assign invert0732 = nor1730;
assign nor1731 = !(nand0977|nand0983|nand0997|nand0991); 
assign invert0733 = nor1731;
assign nor1732 = !(nand0983|nand0997|nand0978|nand0991); 
assign invert0734 = nor1732;
assign nor1733 = !(nand0983|nand0979|nand0997|nand0991); 
assign invert0735 = nor1733;
assign nor1734 = !(nand0997|nand0972|nand0984|nand0991); 
assign invert0736 = nor1734;
assign nor1735 = !(nand0973|nand0997|nand0984|nand0991); 
assign invert0737 = nor1735;
assign nor1736 = !(nand0974|nand0997|nand0984|nand0991); 
assign invert0738 = nor1736;
assign nor1737 = !(nand0997|nand0975|nand0984|nand0991); 
assign invert0739 = nor1737;
assign nor1738 = !(nand0976|nand0997|nand0984|nand0991); 
assign invert0740 = nor1738;
assign nor1739 = !(nand0977|nand0997|nand0984|nand0991); 
assign invert0741 = nor1739;
assign nor1740 = !(nand0997|nand0978|nand0984|nand0991); 
assign invert0742 = nor1740;
assign nor1741 = !(nand0979|nand0997|nand0984|nand0991); 
assign invert0743 = nor1741;
assign nor1742 = !(nand0985|nand0997|nand0972|nand0991); 
assign invert0744 = nor1742;
assign nor1743 = !(nand0973|nand0985|nand0997|nand0991); 
assign invert0745 = nor1743;
assign nor1744 = !(nand0974|nand0985|nand0997|nand0991); 
assign invert0746 = nor1744;
assign nor1745 = !(nand0985|nand0997|nand0975|nand0991); 
assign invert0747 = nor1745;
assign nor1746 = !(nand0976|nand0985|nand0997|nand0991); 
assign invert0748 = nor1746;
assign nor1747 = !(nand0977|nand0985|nand0997|nand0991); 
assign invert0749 = nor1747;
assign nor1748 = !(nand0985|nand0997|nand0978|nand0991); 
assign invert0750 = nor1748;
assign nor1749 = !(nand0979|nand0985|nand0997|nand0991); 
assign invert0751 = nor1749;
assign nor1750 = !(nand0986|nand0997|nand0972|nand0991); 
assign invert0752 = nor1750;
assign nor1751 = !(nand0986|nand0973|nand0997|nand0991); 
assign invert0753 = nor1751;
assign nor1752 = !(nand0986|nand0974|nand0997|nand0991); 
assign invert0754 = nor1752;
assign nor1753 = !(nand0986|nand0997|nand0975|nand0991); 
assign invert0755 = nor1753;
assign nor1754 = !(nand0986|nand0976|nand0997|nand0991); 
assign invert0756 = nor1754;
assign nor1755 = !(nand0977|nand0986|nand0997|nand0991); 
assign invert0757 = nor1755;
assign nor1756 = !(nand0986|nand0997|nand0978|nand0991); 
assign invert0758 = nor1756;
assign nor1757 = !(nand0986|nand0979|nand0997|nand0991); 
assign invert0759 = nor1757;
assign nor1758 = !(nand0997|nand0987|nand0972|nand0991); 
assign invert0760 = nor1758;
assign nor1759 = !(nand0973|nand0997|nand0987|nand0991); 
assign invert0761 = nor1759;
assign nor1760 = !(nand0974|nand0997|nand0987|nand0991); 
assign invert0762 = nor1760;
assign nor1761 = !(nand0997|nand0987|nand0975|nand0991); 
assign invert0763 = nor1761;
assign nor1762 = !(nand0976|nand0997|nand0987|nand0991); 
assign invert0764 = nor1762;
assign nor1763 = !(nand0977|nand0997|nand0987|nand0991); 
assign invert0765 = nor1763;
assign nor1764 = !(nand0997|nand0978|nand0987|nand0991); 
assign invert0766 = nor1764;
assign nor1765 = !(nand0979|nand0997|nand0987|nand0991); 
assign invert0767 = nor1765;
assign nor1766 = !(nand0980|nand0992|nand0997|nand0972); 
assign invert0768 = nor1766;
assign nor1767 = !(nand0980|nand0973|nand0992|nand0997); 
assign invert0769 = nor1767;
assign nor1768 = !(nand0974|nand0980|nand0992|nand0997); 
assign invert0770 = nor1768;
assign nor1769 = !(nand0980|nand0992|nand0997|nand0975); 
assign invert0771 = nor1769;
assign nor1770 = !(nand0980|nand0976|nand0992|nand0997); 
assign invert0772 = nor1770;
assign nor1771 = !(nand0977|nand0980|nand0992|nand0997); 
assign invert0773 = nor1771;
assign nor1772 = !(nand0980|nand0992|nand0997|nand0978); 
assign invert0774 = nor1772;
assign nor1773 = !(nand0979|nand0980|nand0992|nand0997); 
assign invert0775 = nor1773;
assign nor1774 = !(nand0992|nand0997|nand0972|nand0981); 
assign invert0776 = nor1774;
assign nor1775 = !(nand0973|nand0992|nand0997|nand0981); 
assign invert0777 = nor1775;
assign nor1776 = !(nand0974|nand0992|nand0997|nand0981); 
assign invert0778 = nor1776;
assign nor1777 = !(nand0992|nand0997|nand0975|nand0981); 
assign invert0779 = nor1777;
assign nor1778 = !(nand0976|nand0992|nand0997|nand0981); 
assign invert0780 = nor1778;
assign nor1779 = !(nand0977|nand0992|nand0997|nand0981); 
assign invert0781 = nor1779;
assign nor1780 = !(nand0992|nand0997|nand0978|nand0981); 
assign invert0782 = nor1780;
assign nor1781 = !(nand0979|nand0992|nand0997|nand0981); 
assign invert0783 = nor1781;
assign nor1782 = !(nand0992|nand0982|nand0997|nand0972); 
assign invert0784 = nor1782;
assign nor1783 = !(nand0973|nand0992|nand0982|nand0997); 
assign invert0785 = nor1783;
assign nor1784 = !(nand0974|nand0992|nand0982|nand0997); 
assign invert0786 = nor1784;
assign nor1785 = !(nand0992|nand0982|nand0997|nand0975); 
assign invert0787 = nor1785;
assign nor1786 = !(nand0976|nand0992|nand0982|nand0997); 
assign invert0788 = nor1786;
assign nor1787 = !(nand0977|nand0992|nand0982|nand0997); 
assign invert0789 = nor1787;
assign nor1788 = !(nand0992|nand0982|nand0997|nand0978); 
assign invert0790 = nor1788;
assign nor1789 = !(nand0979|nand0992|nand0982|nand0997); 
assign invert0791 = nor1789;
assign nor1790 = !(nand0983|nand0992|nand0997|nand0972); 
assign invert0792 = nor1790;
assign nor1791 = !(nand0983|nand0973|nand0992|nand0997); 
assign invert0793 = nor1791;
assign nor1792 = !(nand0974|nand0983|nand0992|nand0997); 
assign invert0794 = nor1792;
assign nor1793 = !(nand0983|nand0992|nand0997|nand0975); 
assign invert0795 = nor1793;
assign nor1794 = !(nand0983|nand0976|nand0992|nand0997); 
assign invert0796 = nor1794;
assign nor1795 = !(nand0977|nand0983|nand0992|nand0997); 
assign invert0797 = nor1795;
assign nor1796 = !(nand0983|nand0992|nand0997|nand0978); 
assign invert0798 = nor1796;
assign nor1797 = !(nand0983|nand0979|nand0992|nand0997); 
assign invert0799 = nor1797;
assign nor1798 = !(nand0992|nand0997|nand0972|nand0984); 
assign invert0800 = nor1798;
assign nor1799 = !(nand0973|nand0992|nand0997|nand0984); 
assign invert0801 = nor1799;
assign nor1800 = !(nand0974|nand0992|nand0997|nand0984); 
assign invert0802 = nor1800;
assign nor1801 = !(nand0992|nand0997|nand0975|nand0984); 
assign invert0803 = nor1801;
assign nor1802 = !(nand0976|nand0992|nand0997|nand0984); 
assign invert0804 = nor1802;
assign nor1803 = !(nand0977|nand0992|nand0997|nand0984); 
assign invert0805 = nor1803;
assign nor1804 = !(nand0992|nand0997|nand0978|nand0984); 
assign invert0806 = nor1804;
assign nor1805 = !(nand0979|nand0992|nand0997|nand0984); 
assign invert0807 = nor1805;
assign nor1806 = !(nand0985|nand0992|nand0997|nand0972); 
assign invert0808 = nor1806;
assign nor1807 = !(nand0973|nand0985|nand0992|nand0997); 
assign invert0809 = nor1807;
assign nor1808 = !(nand0974|nand0985|nand0992|nand0997); 
assign invert0810 = nor1808;
assign nor1809 = !(nand0985|nand0992|nand0997|nand0975); 
assign invert0811 = nor1809;
assign nor1810 = !(nand0976|nand0985|nand0992|nand0997); 
assign invert0812 = nor1810;
assign nor1811 = !(nand0977|nand0985|nand0992|nand0997); 
assign invert0813 = nor1811;
assign nor1812 = !(nand0985|nand0992|nand0997|nand0978); 
assign invert0814 = nor1812;
assign nor1813 = !(nand0979|nand0985|nand0992|nand0997); 
assign invert0815 = nor1813;
assign nor1814 = !(nand0986|nand0992|nand0997|nand0972); 
assign invert0816 = nor1814;
assign nor1815 = !(nand0986|nand0973|nand0992|nand0997); 
assign invert0817 = nor1815;
assign nor1816 = !(nand0986|nand0974|nand0992|nand0997); 
assign invert0818 = nor1816;
assign nor1817 = !(nand0986|nand0992|nand0997|nand0975); 
assign invert0819 = nor1817;
assign nor1818 = !(nand0986|nand0976|nand0992|nand0997); 
assign invert0820 = nor1818;
assign nor1819 = !(nand0977|nand0986|nand0992|nand0997); 
assign invert0821 = nor1819;
assign nor1820 = !(nand0986|nand0992|nand0997|nand0978); 
assign invert0822 = nor1820;
assign nor1821 = !(nand0986|nand0979|nand0992|nand0997); 
assign invert0823 = nor1821;
assign nor1822 = !(nand0992|nand0997|nand0987|nand0972); 
assign invert0824 = nor1822;
assign nor1823 = !(nand0973|nand0992|nand0997|nand0987); 
assign invert0825 = nor1823;
assign nor1824 = !(nand0974|nand0992|nand0997|nand0987); 
assign invert0826 = nor1824;
assign nor1825 = !(nand0992|nand0997|nand0987|nand0975); 
assign invert0827 = nor1825;
assign nor1826 = !(nand0976|nand0992|nand0997|nand0987); 
assign invert0828 = nor1826;
assign nor1827 = !(nand0977|nand0992|nand0997|nand0987); 
assign invert0829 = nor1827;
assign nor1828 = !(nand0992|nand0997|nand0978|nand0987); 
assign invert0830 = nor1828;
assign nor1829 = !(nand0979|nand0992|nand0997|nand0987); 
assign invert0831 = nor1829;
assign nor1830 = !(nand0993|nand0980|nand0997|nand0972); 
assign invert0832 = nor1830;
assign nor1831 = !(nand0993|nand0980|nand0973|nand0997); 
assign invert0833 = nor1831;
assign nor1832 = !(nand0993|nand0974|nand0980|nand0997); 
assign invert0834 = nor1832;
assign nor1833 = !(nand0993|nand0980|nand0997|nand0975); 
assign invert0835 = nor1833;
assign nor1834 = !(nand0993|nand0980|nand0976|nand0997); 
assign invert0836 = nor1834;
assign nor1835 = !(nand0977|nand0993|nand0980|nand0997); 
assign invert0837 = nor1835;
assign nor1836 = !(nand0993|nand0980|nand0997|nand0978); 
assign invert0838 = nor1836;
assign nor1837 = !(nand0993|nand0979|nand0980|nand0997); 
assign invert0839 = nor1837;
assign nor1838 = !(nand0993|nand0997|nand0972|nand0981); 
assign invert0840 = nor1838;
assign nor1839 = !(nand0993|nand0973|nand0997|nand0981); 
assign invert0841 = nor1839;
assign nor1840 = !(nand0993|nand0974|nand0997|nand0981); 
assign invert0842 = nor1840;
assign nor1841 = !(nand0993|nand0997|nand0975|nand0981); 
assign invert0843 = nor1841;
assign nor1842 = !(nand0993|nand0976|nand0997|nand0981); 
assign invert0844 = nor1842;
assign nor1843 = !(nand0977|nand0993|nand0997|nand0981); 
assign invert0845 = nor1843;
assign nor1844 = !(nand0993|nand0997|nand0978|nand0981); 
assign invert0846 = nor1844;
assign nor1845 = !(nand0993|nand0979|nand0997|nand0981); 
assign invert0847 = nor1845;
assign nor1846 = !(nand0993|nand0982|nand0997|nand0972); 
assign invert0848 = nor1846;
assign nor1847 = !(nand0993|nand0973|nand0982|nand0997); 
assign invert0849 = nor1847;
assign nor1848 = !(nand0993|nand0974|nand0982|nand0997); 
assign invert0850 = nor1848;
assign nor1849 = !(nand0993|nand0982|nand0997|nand0975); 
assign invert0851 = nor1849;
assign nor1850 = !(nand0993|nand0976|nand0982|nand0997); 
assign invert0852 = nor1850;
assign nor1851 = !(nand0977|nand0993|nand0982|nand0997); 
assign invert0853 = nor1851;
assign nor1852 = !(nand0993|nand0982|nand0997|nand0978); 
assign invert0854 = nor1852;
assign nor1853 = !(nand0993|nand0979|nand0982|nand0997); 
assign invert0855 = nor1853;
assign nor1854 = !(nand0993|nand0983|nand0997|nand0972); 
assign invert0856 = nor1854;
assign nor1855 = !(nand0993|nand0983|nand0973|nand0997); 
assign invert0857 = nor1855;
assign nor1856 = !(nand0993|nand0974|nand0983|nand0997); 
assign invert0858 = nor1856;
assign nor1857 = !(nand0993|nand0983|nand0997|nand0975); 
assign invert0859 = nor1857;
assign nor1858 = !(nand0993|nand0983|nand0976|nand0997); 
assign invert0860 = nor1858;
assign nor1859 = !(nand0977|nand0993|nand0983|nand0997); 
assign invert0861 = nor1859;
assign nor1860 = !(nand0993|nand0983|nand0997|nand0978); 
assign invert0862 = nor1860;
assign nor1861 = !(nand0993|nand0983|nand0979|nand0997); 
assign invert0863 = nor1861;
assign nor1862 = !(nand0993|nand0997|nand0972|nand0984); 
assign invert0864 = nor1862;
assign nor1863 = !(nand0993|nand0973|nand0997|nand0984); 
assign invert0865 = nor1863;
assign nor1864 = !(nand0993|nand0974|nand0997|nand0984); 
assign invert0866 = nor1864;
assign nor1865 = !(nand0993|nand0997|nand0975|nand0984); 
assign invert0867 = nor1865;
assign nor1866 = !(nand0993|nand0976|nand0997|nand0984); 
assign invert0868 = nor1866;
assign nor1867 = !(nand0977|nand0993|nand0997|nand0984); 
assign invert0869 = nor1867;
assign nor1868 = !(nand0993|nand0997|nand0978|nand0984); 
assign invert0870 = nor1868;
assign nor1869 = !(nand0993|nand0979|nand0997|nand0984); 
assign invert0871 = nor1869;
assign nor1870 = !(nand0993|nand0985|nand0997|nand0972); 
assign invert0872 = nor1870;
assign nor1871 = !(nand0993|nand0973|nand0985|nand0997); 
assign invert0873 = nor1871;
assign nor1872 = !(nand0993|nand0974|nand0985|nand0997); 
assign invert0874 = nor1872;
assign nor1873 = !(nand0993|nand0985|nand0997|nand0975); 
assign invert0875 = nor1873;
assign nor1874 = !(nand0993|nand0976|nand0985|nand0997); 
assign invert0876 = nor1874;
assign nor1875 = !(nand0977|nand0993|nand0985|nand0997); 
assign invert0877 = nor1875;
assign nor1876 = !(nand0993|nand0985|nand0997|nand0978); 
assign invert0878 = nor1876;
assign nor1877 = !(nand0993|nand0979|nand0985|nand0997); 
assign invert0879 = nor1877;
assign nor1878 = !(nand0986|nand0993|nand0997|nand0972); 
assign invert0880 = nor1878;
assign nor1879 = !(nand0986|nand0993|nand0973|nand0997); 
assign invert0881 = nor1879;
assign nor1880 = !(nand0986|nand0993|nand0974|nand0997); 
assign invert0882 = nor1880;
assign nor1881 = !(nand0986|nand0993|nand0997|nand0975); 
assign invert0883 = nor1881;
assign nor1882 = !(nand0986|nand0993|nand0976|nand0997); 
assign invert0884 = nor1882;
assign nor1883 = !(nand0977|nand0986|nand0993|nand0997); 
assign invert0885 = nor1883;
assign nor1884 = !(nand0986|nand0993|nand0997|nand0978); 
assign invert0886 = nor1884;
assign nor1885 = !(nand0986|nand0993|nand0979|nand0997); 
assign invert0887 = nor1885;
assign nor1886 = !(nand0993|nand0997|nand0987|nand0972); 
assign invert0888 = nor1886;
assign nor1887 = !(nand0993|nand0973|nand0997|nand0987); 
assign invert0889 = nor1887;
assign nor1888 = !(nand0993|nand0974|nand0997|nand0987); 
assign invert0890 = nor1888;
assign nor1889 = !(nand0993|nand0997|nand0987|nand0975); 
assign invert0891 = nor1889;
assign nor1890 = !(nand0993|nand0976|nand0997|nand0987); 
assign invert0892 = nor1890;
assign nor1891 = !(nand0977|nand0993|nand0997|nand0987); 
assign invert0893 = nor1891;
assign nor1892 = !(nand0993|nand0997|nand0978|nand0987); 
assign invert0894 = nor1892;
assign nor1893 = !(nand0993|nand0979|nand0997|nand0987); 
assign invert0895 = nor1893;
assign nor1894 = !(nand0980|nand0997|nand0994|nand0972); 
assign invert0896 = nor1894;
assign nor1895 = !(nand0980|nand0973|nand0997|nand0994); 
assign invert0897 = nor1895;
assign nor1896 = !(nand0974|nand0980|nand0997|nand0994); 
assign invert0898 = nor1896;
assign nor1897 = !(nand0980|nand0997|nand0975|nand0994); 
assign invert0899 = nor1897;
assign nor1898 = !(nand0980|nand0976|nand0997|nand0994); 
assign invert0900 = nor1898;
assign nor1899 = !(nand0977|nand0980|nand0997|nand0994); 
assign invert0901 = nor1899;
assign nor1900 = !(nand0980|nand0997|nand0978|nand0994); 
assign invert0902 = nor1900;
assign nor1901 = !(nand0979|nand0980|nand0997|nand0994); 
assign invert0903 = nor1901;
assign nor1902 = !(nand0997|nand0994|nand0972|nand0981); 
assign invert0904 = nor1902;
assign nor1903 = !(nand0973|nand0997|nand0994|nand0981); 
assign invert0905 = nor1903;
assign nor1904 = !(nand0974|nand0997|nand0994|nand0981); 
assign invert0906 = nor1904;
assign nor1905 = !(nand0997|nand0975|nand0994|nand0981); 
assign invert0907 = nor1905;
assign nor1906 = !(nand0976|nand0997|nand0994|nand0981); 
assign invert0908 = nor1906;
assign nor1907 = !(nand0977|nand0997|nand0994|nand0981); 
assign invert0909 = nor1907;
assign nor1908 = !(nand0997|nand0978|nand0994|nand0981); 
assign invert0910 = nor1908;
assign nor1909 = !(nand0979|nand0997|nand0994|nand0981); 
assign invert0911 = nor1909;
assign nor1910 = !(nand0982|nand0997|nand0994|nand0972); 
assign invert0912 = nor1910;
assign nor1911 = !(nand0973|nand0982|nand0997|nand0994); 
assign invert0913 = nor1911;
assign nor1912 = !(nand0974|nand0982|nand0997|nand0994); 
assign invert0914 = nor1912;
assign nor1913 = !(nand0982|nand0997|nand0975|nand0994); 
assign invert0915 = nor1913;
assign nor1914 = !(nand0976|nand0982|nand0997|nand0994); 
assign invert0916 = nor1914;
assign nor1915 = !(nand0977|nand0982|nand0997|nand0994); 
assign invert0917 = nor1915;
assign nor1916 = !(nand0982|nand0997|nand0978|nand0994); 
assign invert0918 = nor1916;
assign nor1917 = !(nand0979|nand0982|nand0997|nand0994); 
assign invert0919 = nor1917;
assign nor1918 = !(nand0983|nand0997|nand0994|nand0972); 
assign invert0920 = nor1918;
assign nor1919 = !(nand0983|nand0973|nand0997|nand0994); 
assign invert0921 = nor1919;
assign nor1920 = !(nand0974|nand0983|nand0997|nand0994); 
assign invert0922 = nor1920;
assign nor1921 = !(nand0983|nand0997|nand0975|nand0994); 
assign invert0923 = nor1921;
assign nor1922 = !(nand0983|nand0976|nand0997|nand0994); 
assign invert0924 = nor1922;
assign nor1923 = !(nand0977|nand0983|nand0997|nand0994); 
assign invert0925 = nor1923;
assign nor1924 = !(nand0983|nand0997|nand0978|nand0994); 
assign invert0926 = nor1924;
assign nor1925 = !(nand0983|nand0979|nand0997|nand0994); 
assign invert0927 = nor1925;
assign nor1926 = !(nand0997|nand0994|nand0972|nand0984); 
assign invert0928 = nor1926;
assign nor1927 = !(nand0973|nand0997|nand0994|nand0984); 
assign invert0929 = nor1927;
assign nor1928 = !(nand0974|nand0997|nand0994|nand0984); 
assign invert0930 = nor1928;
assign nor1929 = !(nand0997|nand0975|nand0994|nand0984); 
assign invert0931 = nor1929;
assign nor1930 = !(nand0976|nand0997|nand0994|nand0984); 
assign invert0932 = nor1930;
assign nor1931 = !(nand0977|nand0997|nand0994|nand0984); 
assign invert0933 = nor1931;
assign nor1932 = !(nand0997|nand0978|nand0994|nand0984); 
assign invert0934 = nor1932;
assign nor1933 = !(nand0979|nand0997|nand0994|nand0984); 
assign invert0935 = nor1933;
assign nor1934 = !(nand0985|nand0997|nand0994|nand0972); 
assign invert0936 = nor1934;
assign nor1935 = !(nand0973|nand0985|nand0997|nand0994); 
assign invert0937 = nor1935;
assign nor1936 = !(nand0974|nand0985|nand0997|nand0994); 
assign invert0938 = nor1936;
assign nor1937 = !(nand0985|nand0997|nand0975|nand0994); 
assign invert0939 = nor1937;
assign nor1938 = !(nand0976|nand0985|nand0997|nand0994); 
assign invert0940 = nor1938;
assign nor1939 = !(nand0977|nand0985|nand0997|nand0994); 
assign invert0941 = nor1939;
assign nor1940 = !(nand0985|nand0997|nand0978|nand0994); 
assign invert0942 = nor1940;
assign nor1941 = !(nand0979|nand0985|nand0997|nand0994); 
assign invert0943 = nor1941;
assign nor1942 = !(nand0986|nand0997|nand0994|nand0972); 
assign invert0944 = nor1942;
assign nor1943 = !(nand0986|nand0973|nand0997|nand0994); 
assign invert0945 = nor1943;
assign nor1944 = !(nand0986|nand0974|nand0997|nand0994); 
assign invert0946 = nor1944;
assign nor1945 = !(nand0986|nand0997|nand0975|nand0994); 
assign invert0947 = nor1945;
assign nor1946 = !(nand0986|nand0976|nand0997|nand0994); 
assign invert0948 = nor1946;
assign nor1947 = !(nand0977|nand0986|nand0997|nand0994); 
assign invert0949 = nor1947;
assign nor1948 = !(nand0986|nand0997|nand0978|nand0994); 
assign invert0950 = nor1948;
assign nor1949 = !(nand0986|nand0979|nand0997|nand0994); 
assign invert0951 = nor1949;
assign nor1950 = !(nand0997|nand0987|nand0994|nand0972); 
assign invert0952 = nor1950;
assign nor1951 = !(nand0973|nand0997|nand0987|nand0994); 
assign invert0953 = nor1951;
assign nor1952 = !(nand0974|nand0997|nand0987|nand0994); 
assign invert0954 = nor1952;
assign nor1953 = !(nand0997|nand0987|nand0975|nand0994); 
assign invert0955 = nor1953;
assign nor1954 = !(nand0976|nand0997|nand0987|nand0994); 
assign invert0956 = nor1954;
assign nor1955 = !(nand0977|nand0997|nand0987|nand0994); 
assign invert0957 = nor1955;
assign nor1956 = !(nand0997|nand0978|nand0987|nand0994); 
assign invert0958 = nor1956;
assign nor1957 = !(nand0979|nand0997|nand0987|nand0994); 
assign invert0959 = nor1957;
assign nor1958 = !(nand0980|nand0995|nand0997|nand0972); 
assign invert0960 = nor1958;
assign nor1959 = !(nand0980|nand0995|nand0973|nand0997); 
assign invert0961 = nor1959;
assign nor1960 = !(nand0974|nand0980|nand0995|nand0997); 
assign invert0962 = nor1960;
assign nor1961 = !(nand0980|nand0995|nand0997|nand0975); 
assign invert0963 = nor1961;
assign nor1962 = !(nand0980|nand0976|nand0995|nand0997); 
assign invert0964 = nor1962;
assign nor1963 = !(nand0977|nand0980|nand0995|nand0997); 
assign invert0965 = nor1963;
assign nor1964 = !(nand0980|nand0995|nand0997|nand0978); 
assign invert0966 = nor1964;
assign nor1965 = !(nand0979|nand0980|nand0995|nand0997); 
assign invert0967 = nor1965;
assign nor1966 = !(nand0995|nand0997|nand0972|nand0981); 
assign invert0968 = nor1966;
assign nor1967 = !(nand0995|nand0973|nand0997|nand0981); 
assign invert0969 = nor1967;
assign nor1968 = !(nand0974|nand0995|nand0997|nand0981); 
assign invert0970 = nor1968;
assign nor1969 = !(nand0995|nand0997|nand0975|nand0981); 
assign invert0971 = nor1969;
assign nor1970 = !(nand0976|nand0995|nand0997|nand0981); 
assign invert0972 = nor1970;
assign nor1971 = !(nand0977|nand0995|nand0997|nand0981); 
assign invert0973 = nor1971;
assign nor1972 = !(nand0995|nand0997|nand0978|nand0981); 
assign invert0974 = nor1972;
assign nor1973 = !(nand0979|nand0995|nand0997|nand0981); 
assign invert0975 = nor1973;
assign nor1974 = !(nand0995|nand0982|nand0997|nand0972); 
assign invert0976 = nor1974;
assign nor1975 = !(nand0995|nand0973|nand0982|nand0997); 
assign invert0977 = nor1975;
assign nor1976 = !(nand0974|nand0995|nand0982|nand0997); 
assign invert0978 = nor1976;
assign nor1977 = !(nand0995|nand0982|nand0997|nand0975); 
assign invert0979 = nor1977;
assign nor1978 = !(nand0976|nand0995|nand0982|nand0997); 
assign invert0980 = nor1978;
assign nor1979 = !(nand0977|nand0995|nand0982|nand0997); 
assign invert0981 = nor1979;
assign nor1980 = !(nand0995|nand0982|nand0997|nand0978); 
assign invert0982 = nor1980;
assign nor1981 = !(nand0979|nand0995|nand0982|nand0997); 
assign invert0983 = nor1981;
assign nor1982 = !(nand0983|nand0995|nand0997|nand0972); 
assign invert0984 = nor1982;
assign nor1983 = !(nand0983|nand0995|nand0973|nand0997); 
assign invert0985 = nor1983;
assign nor1984 = !(nand0974|nand0983|nand0995|nand0997); 
assign invert0986 = nor1984;
assign nor1985 = !(nand0983|nand0995|nand0997|nand0975); 
assign invert0987 = nor1985;
assign nor1986 = !(nand0983|nand0976|nand0995|nand0997); 
assign invert0988 = nor1986;
assign nor1987 = !(nand0977|nand0983|nand0995|nand0997); 
assign invert0989 = nor1987;
assign nor1988 = !(nand0983|nand0995|nand0997|nand0978); 
assign invert0990 = nor1988;
assign nor1989 = !(nand0983|nand0979|nand0995|nand0997); 
assign invert0991 = nor1989;
assign nor1990 = !(nand0995|nand0997|nand0972|nand0984); 
assign invert0992 = nor1990;
assign nor1991 = !(nand0995|nand0973|nand0997|nand0984); 
assign invert0993 = nor1991;
assign nor1992 = !(nand0974|nand0995|nand0997|nand0984); 
assign invert0994 = nor1992;
assign nor1993 = !(nand0995|nand0997|nand0975|nand0984); 
assign invert0995 = nor1993;
assign nor1994 = !(nand0976|nand0995|nand0997|nand0984); 
assign invert0996 = nor1994;
assign nor1995 = !(nand0977|nand0995|nand0997|nand0984); 
assign invert0997 = nor1995;
assign nor1996 = !(nand0995|nand0997|nand0978|nand0984); 
assign invert0998 = nor1996;
assign nor1997 = !(nand0979|nand0995|nand0997|nand0984); 
assign invert0999 = nor1997;
assign nor1998 = !(nand0995|nand0985|nand0997|nand0972); 
assign invert1000 = nor1998;
assign nor1999 = !(nand0995|nand0973|nand0985|nand0997); 
assign invert1001 = nor1999;
assign nor2000 = !(nand0974|nand0995|nand0985|nand0997); 
assign invert1002 = nor2000;
assign nor2001 = !(nand0995|nand0985|nand0997|nand0975); 
assign invert1003 = nor2001;
assign nor2002 = !(nand0976|nand0995|nand0985|nand0997); 
assign invert1004 = nor2002;
assign nor2003 = !(nand0977|nand0995|nand0985|nand0997); 
assign invert1005 = nor2003;
assign nor2004 = !(nand0995|nand0985|nand0997|nand0978); 
assign invert1006 = nor2004;
assign nor2005 = !(nand0979|nand0995|nand0985|nand0997); 
assign invert1007 = nor2005;
assign nor2006 = !(nand0986|nand0995|nand0997|nand0972); 
assign invert1008 = nor2006;
assign nor2007 = !(nand0986|nand0995|nand0973|nand0997); 
assign invert1009 = nor2007;
assign nor2008 = !(nand0986|nand0974|nand0995|nand0997); 
assign invert1010 = nor2008;
assign nor2009 = !(nand0986|nand0995|nand0997|nand0975); 
assign invert1011 = nor2009;
assign nor2010 = !(nand0986|nand0976|nand0995|nand0997); 
assign invert1012 = nor2010;
assign nor2011 = !(nand0977|nand0986|nand0995|nand0997); 
assign invert1013 = nor2011;
assign nor2012 = !(nand0986|nand0995|nand0997|nand0978); 
assign invert1014 = nor2012;
assign nor2013 = !(nand0986|nand0979|nand0995|nand0997); 
assign invert1015 = nor2013;
assign nor2014 = !(nand0995|nand0997|nand0987|nand0972); 
assign invert1016 = nor2014;
assign nor2015 = !(nand0995|nand0973|nand0997|nand0987); 
assign invert1017 = nor2015;
assign nor2016 = !(nand0974|nand0995|nand0997|nand0987); 
assign invert1018 = nor2016;
assign nor2017 = !(nand0995|nand0997|nand0987|nand0975); 
assign invert1019 = nor2017;
assign nor2018 = !(nand0976|nand0995|nand0997|nand0987); 
assign invert1020 = nor2018;
assign nor2019 = !(nand0977|nand0995|nand0997|nand0987); 
assign invert1021 = nor2019;
assign nor2020 = !(nand0995|nand0997|nand0978|nand0987); 
assign invert1022 = nor2020;
assign nor2021 = !(nand0979|nand0995|nand0997|nand0987); 
assign invert1023 = nor2021;
assign corrected[0] = (invert0000^input_data[0]); 
assign corrected[1] = (invert0001^input_data[1]); 
assign corrected[2] = (input_data[2]^invert0002); 
assign corrected[3] = (input_data[3]^invert0003); 
assign corrected[4] = (invert0004^input_data[4]); 
assign corrected[5] = (input_data[5]^invert0005); 
assign corrected[6] = (input_data[6]^invert0006); 
assign corrected[7] = (invert0007^input_data[7]); 
assign corrected[8] = (input_data[8]^invert0008); 
assign corrected[9] = (input_data[9]^invert0009); 
assign corrected[10] = (input_data[10]^invert0010); 
assign corrected[11] = (invert0011^input_data[11]); 
assign corrected[12] = (input_data[12]^invert0012); 
assign corrected[13] = (input_data[13]^invert0013); 
assign corrected[14] = (input_data[14]^invert0014); 
assign corrected[15] = (input_data[15]^invert0015); 
assign corrected[16] = (input_data[16]^invert0016); 
assign corrected[17] = (invert0017^input_data[17]); 
assign corrected[18] = (invert0018^input_data[18]); 
assign corrected[19] = (invert0019^input_data[19]); 
assign corrected[20] = (input_data[20]^invert0020); 
assign corrected[21] = (input_data[21]^invert0021); 
assign corrected[22] = (invert0022^input_data[22]); 
assign corrected[23] = (input_data[23]^invert0023); 
assign corrected[24] = (invert0024^input_data[24]); 
assign corrected[25] = (input_data[25]^invert0025); 
assign corrected[26] = (input_data[26]^invert0026); 
assign corrected[27] = (input_data[27]^invert0027); 
assign corrected[28] = (input_data[28]^invert0028); 
assign corrected[29] = (invert0029^input_data[29]); 
assign corrected[30] = (input_data[30]^invert0030); 
assign corrected[31] = (input_data[31]^invert0031); 
assign corrected[32] = (input_data[32]^invert0032); 
assign corrected[33] = (input_data[33]^invert0033); 
assign corrected[34] = (invert0034^input_data[34]); 
assign corrected[35] = (input_data[35]^invert0035); 
assign corrected[36] = (input_data[36]^invert0036); 
assign corrected[37] = (invert0037^input_data[37]); 
assign corrected[38] = (input_data[38]^invert0038); 
assign corrected[39] = (invert0039^input_data[39]); 
assign corrected[40] = (input_data[40]^invert0040); 
assign corrected[41] = (invert0041^input_data[41]); 
assign corrected[42] = (input_data[42]^invert0042); 
assign corrected[43] = (input_data[43]^invert0043); 
assign corrected[44] = (input_data[44]^invert0044); 
assign corrected[45] = (invert0045^input_data[45]); 
assign corrected[46] = (invert0046^input_data[46]); 
assign corrected[47] = (invert0047^input_data[47]); 
assign corrected[48] = (invert0048^input_data[48]); 
assign corrected[49] = (invert0049^input_data[49]); 
assign corrected[50] = (invert0050^input_data[50]); 
assign corrected[51] = (input_data[51]^invert0051); 
assign corrected[52] = (input_data[52]^invert0052); 
assign corrected[53] = (input_data[53]^invert0053); 
assign corrected[54] = (input_data[54]^invert0054); 
assign corrected[55] = (invert0055^input_data[55]); 
assign corrected[56] = (invert0056^input_data[56]); 
assign corrected[57] = (invert0057^input_data[57]); 
assign corrected[58] = (invert0058^input_data[58]); 
assign corrected[59] = (invert0059^input_data[59]); 
assign corrected[60] = (invert0060^input_data[60]); 
assign corrected[61] = (invert0061^input_data[61]); 
assign corrected[62] = (invert0062^input_data[62]); 
assign corrected[63] = (invert0063^input_data[63]); 
assign corrected[64] = (invert0064^input_data[64]); 
assign corrected[65] = (input_data[65]^invert0065); 
assign corrected[66] = (invert0066^input_data[66]); 
assign corrected[67] = (input_data[67]^invert0067); 
assign corrected[68] = (input_data[68]^invert0068); 
assign corrected[69] = (invert0069^input_data[69]); 
assign corrected[70] = (invert0070^input_data[70]); 
assign corrected[71] = (invert0071^input_data[71]); 
assign corrected[72] = (invert0072^input_data[72]); 
assign corrected[73] = (invert0073^input_data[73]); 
assign corrected[74] = (invert0074^input_data[74]); 
assign corrected[75] = (input_data[75]^invert0075); 
assign corrected[76] = (invert0076^input_data[76]); 
assign corrected[77] = (input_data[77]^invert0077); 
assign corrected[78] = (input_data[78]^invert0078); 
assign corrected[79] = (invert0079^input_data[79]); 
assign corrected[80] = (invert0080^input_data[80]); 
assign corrected[81] = (input_data[81]^invert0081); 
assign corrected[82] = (invert0082^input_data[82]); 
assign corrected[83] = (invert0083^input_data[83]); 
assign corrected[84] = (input_data[84]^invert0084); 
assign corrected[85] = (input_data[85]^invert0085); 
assign corrected[86] = (input_data[86]^invert0086); 
assign corrected[87] = (input_data[87]^invert0087); 
assign corrected[88] = (input_data[88]^invert0088); 
assign corrected[89] = (input_data[89]^invert0089); 
assign corrected[90] = (invert0090^input_data[90]); 
assign corrected[91] = (input_data[91]^invert0091); 
assign corrected[92] = (invert0092^input_data[92]); 
assign corrected[93] = (input_data[93]^invert0093); 
assign corrected[94] = (input_data[94]^invert0094); 
assign corrected[95] = (input_data[95]^invert0095); 
assign corrected[96] = (input_data[96]^invert0096); 
assign corrected[97] = (input_data[97]^invert0097); 
assign corrected[98] = (input_data[98]^invert0098); 
assign corrected[99] = (invert0099^input_data[99]); 
assign corrected[100] = (input_data[100]^invert0100); 
assign corrected[101] = (input_data[101]^invert0101); 
assign corrected[102] = (input_data[102]^invert0102); 
assign corrected[103] = (invert0103^input_data[103]); 
assign corrected[104] = (invert0104^input_data[104]); 
assign corrected[105] = (input_data[105]^invert0105); 
assign corrected[106] = (input_data[106]^invert0106); 
assign corrected[107] = (input_data[107]^invert0107); 
assign corrected[108] = (invert0108^input_data[108]); 
assign corrected[109] = (invert0109^input_data[109]); 
assign corrected[110] = (input_data[110]^invert0110); 
assign corrected[111] = (invert0111^input_data[111]); 
assign corrected[112] = (invert0112^input_data[112]); 
assign corrected[113] = (invert0113^input_data[113]); 
assign corrected[114] = (invert0114^input_data[114]); 
assign corrected[115] = (input_data[115]^invert0115); 
assign corrected[116] = (input_data[116]^invert0116); 
assign corrected[117] = (input_data[117]^invert0117); 
assign corrected[118] = (invert0118^input_data[118]); 
assign corrected[119] = (invert0119^input_data[119]); 
assign corrected[120] = (input_data[120]^invert0120); 
assign corrected[121] = (input_data[121]^invert0121); 
assign corrected[122] = (input_data[122]^invert0122); 
assign corrected[123] = (input_data[123]^invert0123); 
assign corrected[124] = (invert0124^input_data[124]); 
assign corrected[125] = (input_data[125]^invert0125); 
assign corrected[126] = (invert0126^input_data[126]); 
assign corrected[127] = (invert0127^input_data[127]); 
assign corrected[128] = (invert0128^input_data[128]); 
assign corrected[129] = (invert0129^input_data[129]); 
assign corrected[130] = (input_data[130]^invert0130); 
assign corrected[131] = (input_data[131]^invert0131); 
assign corrected[132] = (input_data[132]^invert0132); 
assign corrected[133] = (input_data[133]^invert0133); 
assign corrected[134] = (invert0134^input_data[134]); 
assign corrected[135] = (input_data[135]^invert0135); 
assign corrected[136] = (input_data[136]^invert0136); 
assign corrected[137] = (invert0137^input_data[137]); 
assign corrected[138] = (invert0138^input_data[138]); 
assign corrected[139] = (invert0139^input_data[139]); 
assign corrected[140] = (invert0140^input_data[140]); 
assign corrected[141] = (input_data[141]^invert0141); 
assign corrected[142] = (invert0142^input_data[142]); 
assign corrected[143] = (invert0143^input_data[143]); 
assign corrected[144] = (invert0144^input_data[144]); 
assign corrected[145] = (invert0145^input_data[145]); 
assign corrected[146] = (invert0146^input_data[146]); 
assign corrected[147] = (invert0147^input_data[147]); 
assign corrected[148] = (input_data[148]^invert0148); 
assign corrected[149] = (input_data[149]^invert0149); 
assign corrected[150] = (invert0150^input_data[150]); 
assign corrected[151] = (input_data[151]^invert0151); 
assign corrected[152] = (invert0152^input_data[152]); 
assign corrected[153] = (invert0153^input_data[153]); 
assign corrected[154] = (invert0154^input_data[154]); 
assign corrected[155] = (invert0155^input_data[155]); 
assign corrected[156] = (invert0156^input_data[156]); 
assign corrected[157] = (invert0157^input_data[157]); 
assign corrected[158] = (input_data[158]^invert0158); 
assign corrected[159] = (input_data[159]^invert0159); 
assign corrected[160] = (invert0160^input_data[160]); 
assign corrected[161] = (invert0161^input_data[161]); 
assign corrected[162] = (invert0162^input_data[162]); 
assign corrected[163] = (invert0163^input_data[163]); 
assign corrected[164] = (input_data[164]^invert0164); 
assign corrected[165] = (input_data[165]^invert0165); 
assign corrected[166] = (input_data[166]^invert0166); 
assign corrected[167] = (input_data[167]^invert0167); 
assign corrected[168] = (input_data[168]^invert0168); 
assign corrected[169] = (invert0169^input_data[169]); 
assign corrected[170] = (invert0170^input_data[170]); 
assign corrected[171] = (invert0171^input_data[171]); 
assign corrected[172] = (invert0172^input_data[172]); 
assign corrected[173] = (invert0173^input_data[173]); 
assign corrected[174] = (input_data[174]^invert0174); 
assign corrected[175] = (input_data[175]^invert0175); 
assign corrected[176] = (invert0176^input_data[176]); 
assign corrected[177] = (invert0177^input_data[177]); 
assign corrected[178] = (input_data[178]^invert0178); 
assign corrected[179] = (invert0179^input_data[179]); 
assign corrected[180] = (invert0180^input_data[180]); 
assign corrected[181] = (input_data[181]^invert0181); 
assign corrected[182] = (input_data[182]^invert0182); 
assign corrected[183] = (input_data[183]^invert0183); 
assign corrected[184] = (input_data[184]^invert0184); 
assign corrected[185] = (invert0185^input_data[185]); 
assign corrected[186] = (input_data[186]^invert0186); 
assign corrected[187] = (input_data[187]^invert0187); 
assign corrected[188] = (invert0188^input_data[188]); 
assign corrected[189] = (invert0189^input_data[189]); 
assign corrected[190] = (invert0190^input_data[190]); 
assign corrected[191] = (input_data[191]^invert0191); 
assign corrected[192] = (input_data[192]^invert0192); 
assign corrected[193] = (input_data[193]^invert0193); 
assign corrected[194] = (input_data[194]^invert0194); 
assign corrected[195] = (invert0195^input_data[195]); 
assign corrected[196] = (input_data[196]^invert0196); 
assign corrected[197] = (input_data[197]^invert0197); 
assign corrected[198] = (invert0198^input_data[198]); 
assign corrected[199] = (input_data[199]^invert0199); 
assign corrected[200] = (invert0200^input_data[200]); 
assign corrected[201] = (invert0201^input_data[201]); 
assign corrected[202] = (input_data[202]^invert0202); 
assign corrected[203] = (invert0203^input_data[203]); 
assign corrected[204] = (invert0204^input_data[204]); 
assign corrected[205] = (invert0205^input_data[205]); 
assign corrected[206] = (invert0206^input_data[206]); 
assign corrected[207] = (invert0207^input_data[207]); 
assign corrected[208] = (input_data[208]^invert0208); 
assign corrected[209] = (invert0209^input_data[209]); 
assign corrected[210] = (invert0210^input_data[210]); 
assign corrected[211] = (invert0211^input_data[211]); 
assign corrected[212] = (input_data[212]^invert0212); 
assign corrected[213] = (invert0213^input_data[213]); 
assign corrected[214] = (invert0214^input_data[214]); 
assign corrected[215] = (invert0215^input_data[215]); 
assign corrected[216] = (invert0216^input_data[216]); 
assign corrected[217] = (input_data[217]^invert0217); 
assign corrected[218] = (input_data[218]^invert0218); 
assign corrected[219] = (invert0219^input_data[219]); 
assign corrected[220] = (invert0220^input_data[220]); 
assign corrected[221] = (invert0221^input_data[221]); 
assign corrected[222] = (invert0222^input_data[222]); 
assign corrected[223] = (invert0223^input_data[223]); 
assign corrected[224] = (invert0224^input_data[224]); 
assign corrected[225] = (input_data[225]^invert0225); 
assign corrected[226] = (input_data[226]^invert0226); 
assign corrected[227] = (input_data[227]^invert0227); 
assign corrected[228] = (input_data[228]^invert0228); 
assign corrected[229] = (invert0229^input_data[229]); 
assign corrected[230] = (invert0230^input_data[230]); 
assign corrected[231] = (invert0231^input_data[231]); 
assign corrected[232] = (invert0232^input_data[232]); 
assign corrected[233] = (invert0233^input_data[233]); 
assign corrected[234] = (invert0234^input_data[234]); 
assign corrected[235] = (input_data[235]^invert0235); 
assign corrected[236] = (input_data[236]^invert0236); 
assign corrected[237] = (invert0237^input_data[237]); 
assign corrected[238] = (input_data[238]^invert0238); 
assign corrected[239] = (invert0239^input_data[239]); 
assign corrected[240] = (invert0240^input_data[240]); 
assign corrected[241] = (input_data[241]^invert0241); 
assign corrected[242] = (input_data[242]^invert0242); 
assign corrected[243] = (invert0243^input_data[243]); 
assign corrected[244] = (input_data[244]^invert0244); 
assign corrected[245] = (invert0245^input_data[245]); 
assign corrected[246] = (input_data[246]^invert0246); 
assign corrected[247] = (input_data[247]^invert0247); 
assign corrected[248] = (invert0248^input_data[248]); 
assign corrected[249] = (input_data[249]^invert0249); 
assign corrected[250] = (invert0250^input_data[250]); 
assign corrected[251] = (input_data[251]^invert0251); 
assign corrected[252] = (input_data[252]^invert0252); 
assign corrected[253] = (invert0253^input_data[253]); 
assign corrected[254] = (input_data[254]^invert0254); 
assign corrected[255] = (invert0255^input_data[255]); 
assign corrected[256] = (input_data[256]^invert0256); 
assign corrected[257] = (input_data[257]^invert0257); 
assign corrected[258] = (invert0258^input_data[258]); 
assign corrected[259] = (input_data[259]^invert0259); 
assign corrected[260] = (invert0260^input_data[260]); 
assign corrected[261] = (input_data[261]^invert0261); 
assign corrected[262] = (input_data[262]^invert0262); 
assign corrected[263] = (invert0263^input_data[263]); 
assign corrected[264] = (input_data[264]^invert0264); 
assign corrected[265] = (invert0265^input_data[265]); 
assign corrected[266] = (invert0266^input_data[266]); 
assign corrected[267] = (input_data[267]^invert0267); 
assign corrected[268] = (input_data[268]^invert0268); 
assign corrected[269] = (invert0269^input_data[269]); 
assign corrected[270] = (invert0270^input_data[270]); 
assign corrected[271] = (input_data[271]^invert0271); 
assign corrected[272] = (input_data[272]^invert0272); 
assign corrected[273] = (invert0273^input_data[273]); 
assign corrected[274] = (input_data[274]^invert0274); 
assign corrected[275] = (invert0275^input_data[275]); 
assign corrected[276] = (invert0276^input_data[276]); 
assign corrected[277] = (input_data[277]^invert0277); 
assign corrected[278] = (input_data[278]^invert0278); 
assign corrected[279] = (invert0279^input_data[279]); 
assign corrected[280] = (invert0280^input_data[280]); 
assign corrected[281] = (invert0281^input_data[281]); 
assign corrected[282] = (invert0282^input_data[282]); 
assign corrected[283] = (input_data[283]^invert0283); 
assign corrected[284] = (input_data[284]^invert0284); 
assign corrected[285] = (invert0285^input_data[285]); 
assign corrected[286] = (input_data[286]^invert0286); 
assign corrected[287] = (input_data[287]^invert0287); 
assign corrected[288] = (invert0288^input_data[288]); 
assign corrected[289] = (input_data[289]^invert0289); 
assign corrected[290] = (input_data[290]^invert0290); 
assign corrected[291] = (invert0291^input_data[291]); 
assign corrected[292] = (invert0292^input_data[292]); 
assign corrected[293] = (input_data[293]^invert0293); 
assign corrected[294] = (input_data[294]^invert0294); 
assign corrected[295] = (invert0295^input_data[295]); 
assign corrected[296] = (input_data[296]^invert0296); 
assign corrected[297] = (invert0297^input_data[297]); 
assign corrected[298] = (input_data[298]^invert0298); 
assign corrected[299] = (input_data[299]^invert0299); 
assign corrected[300] = (invert0300^input_data[300]); 
assign corrected[301] = (input_data[301]^invert0301); 
assign corrected[302] = (input_data[302]^invert0302); 
assign corrected[303] = (invert0303^input_data[303]); 
assign corrected[304] = (input_data[304]^invert0304); 
assign corrected[305] = (invert0305^input_data[305]); 
assign corrected[306] = (invert0306^input_data[306]); 
assign corrected[307] = (input_data[307]^invert0307); 
assign corrected[308] = (invert0308^input_data[308]); 
assign corrected[309] = (invert0309^input_data[309]); 
assign corrected[310] = (invert0310^input_data[310]); 
assign corrected[311] = (input_data[311]^invert0311); 
assign corrected[312] = (input_data[312]^invert0312); 
assign corrected[313] = (invert0313^input_data[313]); 
assign corrected[314] = (input_data[314]^invert0314); 
assign corrected[315] = (invert0315^input_data[315]); 
assign corrected[316] = (invert0316^input_data[316]); 
assign corrected[317] = (input_data[317]^invert0317); 
assign corrected[318] = (invert0318^input_data[318]); 
assign corrected[319] = (input_data[319]^invert0319); 
assign corrected[320] = (invert0320^input_data[320]); 
assign corrected[321] = (invert0321^input_data[321]); 
assign corrected[322] = (input_data[322]^invert0322); 
assign corrected[323] = (invert0323^input_data[323]); 
assign corrected[324] = (invert0324^input_data[324]); 
assign corrected[325] = (invert0325^input_data[325]); 
assign corrected[326] = (invert0326^input_data[326]); 
assign corrected[327] = (input_data[327]^invert0327); 
assign corrected[328] = (input_data[328]^invert0328); 
assign corrected[329] = (input_data[329]^invert0329); 
assign corrected[330] = (invert0330^input_data[330]); 
assign corrected[331] = (invert0331^input_data[331]); 
assign corrected[332] = (input_data[332]^invert0332); 
assign corrected[333] = (invert0333^input_data[333]); 
assign corrected[334] = (input_data[334]^invert0334); 
assign corrected[335] = (invert0335^input_data[335]); 
assign corrected[336] = (invert0336^input_data[336]); 
assign corrected[337] = (input_data[337]^invert0337); 
assign corrected[338] = (input_data[338]^invert0338); 
assign corrected[339] = (invert0339^input_data[339]); 
assign corrected[340] = (input_data[340]^invert0340); 
assign corrected[341] = (invert0341^input_data[341]); 
assign corrected[342] = (invert0342^input_data[342]); 
assign corrected[343] = (input_data[343]^invert0343); 
assign corrected[344] = (input_data[344]^invert0344); 
assign corrected[345] = (input_data[345]^invert0345); 
assign corrected[346] = (input_data[346]^invert0346); 
assign corrected[347] = (input_data[347]^invert0347); 
assign corrected[348] = (invert0348^input_data[348]); 
assign corrected[349] = (input_data[349]^invert0349); 
assign corrected[350] = (invert0350^input_data[350]); 
assign corrected[351] = (invert0351^input_data[351]); 
assign corrected[352] = (invert0352^input_data[352]); 
assign corrected[353] = (input_data[353]^invert0353); 
assign corrected[354] = (input_data[354]^invert0354); 
assign corrected[355] = (input_data[355]^invert0355); 
assign corrected[356] = (input_data[356]^invert0356); 
assign corrected[357] = (invert0357^input_data[357]); 
assign corrected[358] = (invert0358^input_data[358]); 
assign corrected[359] = (input_data[359]^invert0359); 
assign corrected[360] = (invert0360^input_data[360]); 
assign corrected[361] = (input_data[361]^invert0361); 
assign corrected[362] = (input_data[362]^invert0362); 
assign corrected[363] = (input_data[363]^invert0363); 
assign corrected[364] = (input_data[364]^invert0364); 
assign corrected[365] = (invert0365^input_data[365]); 
assign corrected[366] = (invert0366^input_data[366]); 
assign corrected[367] = (input_data[367]^invert0367); 
assign corrected[368] = (invert0368^input_data[368]); 
assign corrected[369] = (input_data[369]^invert0369); 
assign corrected[370] = (invert0370^input_data[370]); 
assign corrected[371] = (input_data[371]^invert0371); 
assign corrected[372] = (invert0372^input_data[372]); 
assign corrected[373] = (invert0373^input_data[373]); 
assign corrected[374] = (input_data[374]^invert0374); 
assign corrected[375] = (invert0375^input_data[375]); 
assign corrected[376] = (input_data[376]^invert0376); 
assign corrected[377] = (input_data[377]^invert0377); 
assign corrected[378] = (invert0378^input_data[378]); 
assign corrected[379] = (input_data[379]^invert0379); 
assign corrected[380] = (input_data[380]^invert0380); 
assign corrected[381] = (invert0381^input_data[381]); 
assign corrected[382] = (invert0382^input_data[382]); 
assign corrected[383] = (input_data[383]^invert0383); 
assign corrected[384] = (invert0384^input_data[384]); 
assign corrected[385] = (invert0385^input_data[385]); 
assign corrected[386] = (invert0386^input_data[386]); 
assign corrected[387] = (invert0387^input_data[387]); 
assign corrected[388] = (input_data[388]^invert0388); 
assign corrected[389] = (input_data[389]^invert0389); 
assign corrected[390] = (input_data[390]^invert0390); 
assign corrected[391] = (invert0391^input_data[391]); 
assign corrected[392] = (invert0392^input_data[392]); 
assign corrected[393] = (input_data[393]^invert0393); 
assign corrected[394] = (invert0394^input_data[394]); 
assign corrected[395] = (input_data[395]^invert0395); 
assign corrected[396] = (invert0396^input_data[396]); 
assign corrected[397] = (invert0397^input_data[397]); 
assign corrected[398] = (input_data[398]^invert0398); 
assign corrected[399] = (invert0399^input_data[399]); 
assign corrected[400] = (invert0400^input_data[400]); 
assign corrected[401] = (input_data[401]^invert0401); 
assign corrected[402] = (invert0402^input_data[402]); 
assign corrected[403] = (input_data[403]^invert0403); 
assign corrected[404] = (input_data[404]^invert0404); 
assign corrected[405] = (invert0405^input_data[405]); 
assign corrected[406] = (input_data[406]^invert0406); 
assign corrected[407] = (input_data[407]^invert0407); 
assign corrected[408] = (invert0408^input_data[408]); 
assign corrected[409] = (input_data[409]^invert0409); 
assign corrected[410] = (invert0410^input_data[410]); 
assign corrected[411] = (invert0411^input_data[411]); 
assign corrected[412] = (invert0412^input_data[412]); 
assign corrected[413] = (input_data[413]^invert0413); 
assign corrected[414] = (input_data[414]^invert0414); 
assign corrected[415] = (invert0415^input_data[415]); 
assign corrected[416] = (input_data[416]^invert0416); 
assign corrected[417] = (input_data[417]^invert0417); 
assign corrected[418] = (invert0418^input_data[418]); 
assign corrected[419] = (input_data[419]^invert0419); 
assign corrected[420] = (invert0420^input_data[420]); 
assign corrected[421] = (input_data[421]^invert0421); 
assign corrected[422] = (input_data[422]^invert0422); 
assign corrected[423] = (invert0423^input_data[423]); 
assign corrected[424] = (input_data[424]^invert0424); 
assign corrected[425] = (invert0425^input_data[425]); 
assign corrected[426] = (input_data[426]^invert0426); 
assign corrected[427] = (input_data[427]^invert0427); 
assign corrected[428] = (invert0428^input_data[428]); 
assign corrected[429] = (input_data[429]^invert0429); 
assign corrected[430] = (invert0430^input_data[430]); 
assign corrected[431] = (input_data[431]^invert0431); 
assign corrected[432] = (input_data[432]^invert0432); 
assign corrected[433] = (invert0433^input_data[433]); 
assign corrected[434] = (input_data[434]^invert0434); 
assign corrected[435] = (invert0435^input_data[435]); 
assign corrected[436] = (input_data[436]^invert0436); 
assign corrected[437] = (input_data[437]^invert0437); 
assign corrected[438] = (invert0438^input_data[438]); 
assign corrected[439] = (input_data[439]^invert0439); 
assign corrected[440] = (input_data[440]^invert0440); 
assign corrected[441] = (invert0441^input_data[441]); 
assign corrected[442] = (invert0442^input_data[442]); 
assign corrected[443] = (input_data[443]^invert0443); 
assign corrected[444] = (invert0444^input_data[444]); 
assign corrected[445] = (input_data[445]^invert0445); 
assign corrected[446] = (invert0446^input_data[446]); 
assign corrected[447] = (invert0447^input_data[447]); 
assign corrected[448] = (input_data[448]^invert0448); 
assign corrected[449] = (input_data[449]^invert0449); 
assign corrected[450] = (input_data[450]^invert0450); 
assign corrected[451] = (invert0451^input_data[451]); 
assign corrected[452] = (input_data[452]^invert0452); 
assign corrected[453] = (input_data[453]^invert0453); 
assign corrected[454] = (invert0454^input_data[454]); 
assign corrected[455] = (input_data[455]^invert0455); 
assign corrected[456] = (invert0456^input_data[456]); 
assign corrected[457] = (invert0457^input_data[457]); 
assign corrected[458] = (input_data[458]^invert0458); 
assign corrected[459] = (input_data[459]^invert0459); 
assign corrected[460] = (input_data[460]^invert0460); 
assign corrected[461] = (invert0461^input_data[461]); 
assign corrected[462] = (invert0462^input_data[462]); 
assign corrected[463] = (input_data[463]^invert0463); 
assign corrected[464] = (input_data[464]^invert0464); 
assign corrected[465] = (invert0465^input_data[465]); 
assign corrected[466] = (input_data[466]^invert0466); 
assign corrected[467] = (invert0467^input_data[467]); 
assign corrected[468] = (invert0468^input_data[468]); 
assign corrected[469] = (input_data[469]^invert0469); 
assign corrected[470] = (input_data[470]^invert0470); 
assign corrected[471] = (invert0471^input_data[471]); 
assign corrected[472] = (invert0472^input_data[472]); 
assign corrected[473] = (input_data[473]^invert0473); 
assign corrected[474] = (input_data[474]^invert0474); 
assign corrected[475] = (invert0475^input_data[475]); 
assign corrected[476] = (invert0476^input_data[476]); 
assign corrected[477] = (invert0477^input_data[477]); 
assign corrected[478] = (input_data[478]^invert0478); 
assign corrected[479] = (input_data[479]^invert0479); 
assign corrected[480] = (input_data[480]^invert0480); 
assign corrected[481] = (invert0481^input_data[481]); 
assign corrected[482] = (input_data[482]^invert0482); 
assign corrected[483] = (input_data[483]^invert0483); 
assign corrected[484] = (invert0484^input_data[484]); 
assign corrected[485] = (input_data[485]^invert0485); 
assign corrected[486] = (invert0486^input_data[486]); 
assign corrected[487] = (input_data[487]^invert0487); 
assign corrected[488] = (invert0488^input_data[488]); 
assign corrected[489] = (invert0489^input_data[489]); 
assign corrected[490] = (input_data[490]^invert0490); 
assign corrected[491] = (input_data[491]^invert0491); 
assign corrected[492] = (input_data[492]^invert0492); 
assign corrected[493] = (invert0493^input_data[493]); 
assign corrected[494] = (invert0494^input_data[494]); 
assign corrected[495] = (input_data[495]^invert0495); 
assign corrected[496] = (input_data[496]^invert0496); 
assign corrected[497] = (input_data[497]^invert0497); 
assign corrected[498] = (invert0498^input_data[498]); 
assign corrected[499] = (invert0499^input_data[499]); 
assign corrected[500] = (input_data[500]^invert0500); 
assign corrected[501] = (invert0501^input_data[501]); 
assign corrected[502] = (invert0502^input_data[502]); 
assign corrected[503] = (input_data[503]^invert0503); 
assign corrected[504] = (invert0504^input_data[504]); 
assign corrected[505] = (invert0505^input_data[505]); 
assign corrected[506] = (invert0506^input_data[506]); 
assign corrected[507] = (invert0507^input_data[507]); 
assign corrected[508] = (invert0508^input_data[508]); 
assign corrected[509] = (input_data[509]^invert0509); 
assign corrected[510] = (input_data[510]^invert0510); 
assign corrected[511] = (invert0511^input_data[511]); 
assign corrected[512] = (invert0512^input_data[512]); 
assign corrected[513] = (input_data[513]^invert0513); 
assign corrected[514] = (invert0514^input_data[514]); 
assign corrected[515] = (invert0515^input_data[515]); 
assign corrected[516] = (invert0516^input_data[516]); 
assign corrected[517] = (invert0517^input_data[517]); 
assign corrected[518] = (input_data[518]^invert0518); 
assign corrected[519] = (input_data[519]^invert0519); 
assign corrected[520] = (invert0520^input_data[520]); 
assign corrected[521] = (invert0521^input_data[521]); 
assign corrected[522] = (invert0522^input_data[522]); 
assign corrected[523] = (input_data[523]^invert0523); 
assign corrected[524] = (input_data[524]^invert0524); 
assign corrected[525] = (input_data[525]^invert0525); 
assign corrected[526] = (input_data[526]^invert0526); 
assign corrected[527] = (invert0527^input_data[527]); 
assign corrected[528] = (invert0528^input_data[528]); 
assign corrected[529] = (input_data[529]^invert0529); 
assign corrected[530] = (invert0530^input_data[530]); 
assign corrected[531] = (invert0531^input_data[531]); 
assign corrected[532] = (invert0532^input_data[532]); 
assign corrected[533] = (input_data[533]^invert0533); 
assign corrected[534] = (input_data[534]^invert0534); 
assign corrected[535] = (input_data[535]^invert0535); 
assign corrected[536] = (invert0536^input_data[536]); 
assign corrected[537] = (invert0537^input_data[537]); 
assign corrected[538] = (invert0538^input_data[538]); 
assign corrected[539] = (input_data[539]^invert0539); 
assign corrected[540] = (input_data[540]^invert0540); 
assign corrected[541] = (input_data[541]^invert0541); 
assign corrected[542] = (input_data[542]^invert0542); 
assign corrected[543] = (input_data[543]^invert0543); 
assign corrected[544] = (invert0544^input_data[544]); 
assign corrected[545] = (input_data[545]^invert0545); 
assign corrected[546] = (invert0546^input_data[546]); 
assign corrected[547] = (invert0547^input_data[547]); 
assign corrected[548] = (invert0548^input_data[548]); 
assign corrected[549] = (invert0549^input_data[549]); 
assign corrected[550] = (input_data[550]^invert0550); 
assign corrected[551] = (input_data[551]^invert0551); 
assign corrected[552] = (input_data[552]^invert0552); 
assign corrected[553] = (input_data[553]^invert0553); 
assign corrected[554] = (invert0554^input_data[554]); 
assign corrected[555] = (input_data[555]^invert0555); 
assign corrected[556] = (input_data[556]^invert0556); 
assign corrected[557] = (invert0557^input_data[557]); 
assign corrected[558] = (invert0558^input_data[558]); 
assign corrected[559] = (invert0559^input_data[559]); 
assign corrected[560] = (input_data[560]^invert0560); 
assign corrected[561] = (invert0561^input_data[561]); 
assign corrected[562] = (invert0562^input_data[562]); 
assign corrected[563] = (input_data[563]^invert0563); 
assign corrected[564] = (invert0564^input_data[564]); 
assign corrected[565] = (invert0565^input_data[565]); 
assign corrected[566] = (invert0566^input_data[566]); 
assign corrected[567] = (invert0567^input_data[567]); 
assign corrected[568] = (input_data[568]^invert0568); 
assign corrected[569] = (invert0569^input_data[569]); 
assign corrected[570] = (input_data[570]^invert0570); 
assign corrected[571] = (input_data[571]^invert0571); 
assign corrected[572] = (invert0572^input_data[572]); 
assign corrected[573] = (input_data[573]^invert0573); 
assign corrected[574] = (invert0574^input_data[574]); 
assign corrected[575] = (input_data[575]^invert0575); 
assign corrected[576] = (invert0576^input_data[576]); 
assign corrected[577] = (invert0577^input_data[577]); 
assign corrected[578] = (invert0578^input_data[578]); 
assign corrected[579] = (invert0579^input_data[579]); 
assign corrected[580] = (invert0580^input_data[580]); 
assign corrected[581] = (invert0581^input_data[581]); 
assign corrected[582] = (invert0582^input_data[582]); 
assign corrected[583] = (invert0583^input_data[583]); 
assign corrected[584] = (invert0584^input_data[584]); 
assign corrected[585] = (input_data[585]^invert0585); 
assign corrected[586] = (input_data[586]^invert0586); 
assign corrected[587] = (invert0587^input_data[587]); 
assign corrected[588] = (input_data[588]^invert0588); 
assign corrected[589] = (invert0589^input_data[589]); 
assign corrected[590] = (invert0590^input_data[590]); 
assign corrected[591] = (invert0591^input_data[591]); 
assign corrected[592] = (invert0592^input_data[592]); 
assign corrected[593] = (invert0593^input_data[593]); 
assign corrected[594] = (input_data[594]^invert0594); 
assign corrected[595] = (input_data[595]^invert0595); 
assign corrected[596] = (invert0596^input_data[596]); 
assign corrected[597] = (invert0597^input_data[597]); 
assign corrected[598] = (input_data[598]^invert0598); 
assign corrected[599] = (invert0599^input_data[599]); 
assign corrected[600] = (input_data[600]^invert0600); 
assign corrected[601] = (input_data[601]^invert0601); 
assign corrected[602] = (invert0602^input_data[602]); 
assign corrected[603] = (input_data[603]^invert0603); 
assign corrected[604] = (invert0604^input_data[604]); 
assign corrected[605] = (invert0605^input_data[605]); 
assign corrected[606] = (input_data[606]^invert0606); 
assign corrected[607] = (invert0607^input_data[607]); 
assign corrected[608] = (input_data[608]^invert0608); 
assign corrected[609] = (invert0609^input_data[609]); 
assign corrected[610] = (input_data[610]^invert0610); 
assign corrected[611] = (input_data[611]^invert0611); 
assign corrected[612] = (invert0612^input_data[612]); 
assign corrected[613] = (input_data[613]^invert0613); 
assign corrected[614] = (invert0614^input_data[614]); 
assign corrected[615] = (input_data[615]^invert0615); 
assign corrected[616] = (input_data[616]^invert0616); 
assign corrected[617] = (invert0617^input_data[617]); 
assign corrected[618] = (input_data[618]^invert0618); 
assign corrected[619] = (invert0619^input_data[619]); 
assign corrected[620] = (invert0620^input_data[620]); 
assign corrected[621] = (input_data[621]^invert0621); 
assign corrected[622] = (invert0622^input_data[622]); 
assign corrected[623] = (input_data[623]^invert0623); 
assign corrected[624] = (invert0624^input_data[624]); 
assign corrected[625] = (invert0625^input_data[625]); 
assign corrected[626] = (input_data[626]^invert0626); 
assign corrected[627] = (invert0627^input_data[627]); 
assign corrected[628] = (invert0628^input_data[628]); 
assign corrected[629] = (input_data[629]^invert0629); 
assign corrected[630] = (input_data[630]^invert0630); 
assign corrected[631] = (input_data[631]^invert0631); 
assign corrected[632] = (invert0632^input_data[632]); 
assign corrected[633] = (input_data[633]^invert0633); 
assign corrected[634] = (invert0634^input_data[634]); 
assign corrected[635] = (invert0635^input_data[635]); 
assign corrected[636] = (input_data[636]^invert0636); 
assign corrected[637] = (invert0637^input_data[637]); 
assign corrected[638] = (invert0638^input_data[638]); 
assign corrected[639] = (invert0639^input_data[639]); 
assign corrected[640] = (invert0640^input_data[640]); 
assign corrected[641] = (invert0641^input_data[641]); 
assign corrected[642] = (invert0642^input_data[642]); 
assign corrected[643] = (invert0643^input_data[643]); 
assign corrected[644] = (invert0644^input_data[644]); 
assign corrected[645] = (input_data[645]^invert0645); 
assign corrected[646] = (input_data[646]^invert0646); 
assign corrected[647] = (invert0647^input_data[647]); 
assign corrected[648] = (input_data[648]^invert0648); 
assign corrected[649] = (invert0649^input_data[649]); 
assign corrected[650] = (invert0650^input_data[650]); 
assign corrected[651] = (invert0651^input_data[651]); 
assign corrected[652] = (input_data[652]^invert0652); 
assign corrected[653] = (invert0653^input_data[653]); 
assign corrected[654] = (invert0654^input_data[654]); 
assign corrected[655] = (input_data[655]^invert0655); 
assign corrected[656] = (invert0656^input_data[656]); 
assign corrected[657] = (input_data[657]^invert0657); 
assign corrected[658] = (input_data[658]^invert0658); 
assign corrected[659] = (invert0659^input_data[659]); 
assign corrected[660] = (input_data[660]^invert0660); 
assign corrected[661] = (input_data[661]^invert0661); 
assign corrected[662] = (input_data[662]^invert0662); 
assign corrected[663] = (invert0663^input_data[663]); 
assign corrected[664] = (invert0664^input_data[664]); 
assign corrected[665] = (input_data[665]^invert0665); 
assign corrected[666] = (input_data[666]^invert0666); 
assign corrected[667] = (invert0667^input_data[667]); 
assign corrected[668] = (input_data[668]^invert0668); 
assign corrected[669] = (invert0669^input_data[669]); 
assign corrected[670] = (input_data[670]^invert0670); 
assign corrected[671] = (invert0671^input_data[671]); 
assign corrected[672] = (invert0672^input_data[672]); 
assign corrected[673] = (invert0673^input_data[673]); 
assign corrected[674] = (invert0674^input_data[674]); 
assign corrected[675] = (input_data[675]^invert0675); 
assign corrected[676] = (input_data[676]^invert0676); 
assign corrected[677] = (invert0677^input_data[677]); 
assign corrected[678] = (input_data[678]^invert0678); 
assign corrected[679] = (invert0679^input_data[679]); 
assign corrected[680] = (invert0680^input_data[680]); 
assign corrected[681] = (invert0681^input_data[681]); 
assign corrected[682] = (input_data[682]^invert0682); 
assign corrected[683] = (invert0683^input_data[683]); 
assign corrected[684] = (input_data[684]^invert0684); 
assign corrected[685] = (invert0685^input_data[685]); 
assign corrected[686] = (invert0686^input_data[686]); 
assign corrected[687] = (input_data[687]^invert0687); 
assign corrected[688] = (input_data[688]^invert0688); 
assign corrected[689] = (input_data[689]^invert0689); 
assign corrected[690] = (invert0690^input_data[690]); 
assign corrected[691] = (input_data[691]^invert0691); 
assign corrected[692] = (input_data[692]^invert0692); 
assign corrected[693] = (invert0693^input_data[693]); 
assign corrected[694] = (input_data[694]^invert0694); 
assign corrected[695] = (invert0695^input_data[695]); 
assign corrected[696] = (invert0696^input_data[696]); 
assign corrected[697] = (input_data[697]^invert0697); 
assign corrected[698] = (invert0698^input_data[698]); 
assign corrected[699] = (invert0699^input_data[699]); 
assign corrected[700] = (input_data[700]^invert0700); 
assign corrected[701] = (invert0701^input_data[701]); 
assign corrected[702] = (invert0702^input_data[702]); 
assign corrected[703] = (invert0703^input_data[703]); 
assign corrected[704] = (input_data[704]^invert0704); 
assign corrected[705] = (input_data[705]^invert0705); 
assign corrected[706] = (input_data[706]^invert0706); 
assign corrected[707] = (input_data[707]^invert0707); 
assign corrected[708] = (input_data[708]^invert0708); 
assign corrected[709] = (invert0709^input_data[709]); 
assign corrected[710] = (invert0710^input_data[710]); 
assign corrected[711] = (invert0711^input_data[711]); 
assign corrected[712] = (input_data[712]^invert0712); 
assign corrected[713] = (invert0713^input_data[713]); 
assign corrected[714] = (input_data[714]^invert0714); 
assign corrected[715] = (input_data[715]^invert0715); 
assign corrected[716] = (input_data[716]^invert0716); 
assign corrected[717] = (invert0717^input_data[717]); 
assign corrected[718] = (input_data[718]^invert0718); 
assign corrected[719] = (input_data[719]^invert0719); 
assign corrected[720] = (input_data[720]^invert0720); 
assign corrected[721] = (input_data[721]^invert0721); 
assign corrected[722] = (input_data[722]^invert0722); 
assign corrected[723] = (input_data[723]^invert0723); 
assign corrected[724] = (invert0724^input_data[724]); 
assign corrected[725] = (invert0725^input_data[725]); 
assign corrected[726] = (input_data[726]^invert0726); 
assign corrected[727] = (invert0727^input_data[727]); 
assign corrected[728] = (input_data[728]^invert0728); 
assign corrected[729] = (invert0729^input_data[729]); 
assign corrected[730] = (input_data[730]^invert0730); 
assign corrected[731] = (input_data[731]^invert0731); 
assign corrected[732] = (invert0732^input_data[732]); 
assign corrected[733] = (invert0733^input_data[733]); 
assign corrected[734] = (invert0734^input_data[734]); 
assign corrected[735] = (input_data[735]^invert0735); 
assign corrected[736] = (input_data[736]^invert0736); 
assign corrected[737] = (input_data[737]^invert0737); 
assign corrected[738] = (input_data[738]^invert0738); 
assign corrected[739] = (invert0739^input_data[739]); 
assign corrected[740] = (invert0740^input_data[740]); 
assign corrected[741] = (invert0741^input_data[741]); 
assign corrected[742] = (input_data[742]^invert0742); 
assign corrected[743] = (invert0743^input_data[743]); 
assign corrected[744] = (invert0744^input_data[744]); 
assign corrected[745] = (invert0745^input_data[745]); 
assign corrected[746] = (invert0746^input_data[746]); 
assign corrected[747] = (input_data[747]^invert0747); 
assign corrected[748] = (input_data[748]^invert0748); 
assign corrected[749] = (input_data[749]^invert0749); 
assign corrected[750] = (invert0750^input_data[750]); 
assign corrected[751] = (invert0751^input_data[751]); 
assign corrected[752] = (input_data[752]^invert0752); 
assign corrected[753] = (invert0753^input_data[753]); 
assign corrected[754] = (input_data[754]^invert0754); 
assign corrected[755] = (invert0755^input_data[755]); 
assign corrected[756] = (invert0756^input_data[756]); 
assign corrected[757] = (input_data[757]^invert0757); 
assign corrected[758] = (input_data[758]^invert0758); 
assign corrected[759] = (invert0759^input_data[759]); 
assign corrected[760] = (invert0760^input_data[760]); 
assign corrected[761] = (invert0761^input_data[761]); 
assign corrected[762] = (input_data[762]^invert0762); 
assign corrected[763] = (invert0763^input_data[763]); 
assign corrected[764] = (input_data[764]^invert0764); 
assign corrected[765] = (input_data[765]^invert0765); 
assign corrected[766] = (invert0766^input_data[766]); 
assign corrected[767] = (invert0767^input_data[767]); 
assign corrected[768] = (input_data[768]^invert0768); 
assign corrected[769] = (input_data[769]^invert0769); 
assign corrected[770] = (invert0770^input_data[770]); 
assign corrected[771] = (invert0771^input_data[771]); 
assign corrected[772] = (input_data[772]^invert0772); 
assign corrected[773] = (invert0773^input_data[773]); 
assign corrected[774] = (invert0774^input_data[774]); 
assign corrected[775] = (invert0775^input_data[775]); 
assign corrected[776] = (invert0776^input_data[776]); 
assign corrected[777] = (input_data[777]^invert0777); 
assign corrected[778] = (input_data[778]^invert0778); 
assign corrected[779] = (input_data[779]^invert0779); 
assign corrected[780] = (input_data[780]^invert0780); 
assign corrected[781] = (input_data[781]^invert0781); 
assign corrected[782] = (input_data[782]^invert0782); 
assign corrected[783] = (input_data[783]^invert0783); 
assign corrected[784] = (input_data[784]^invert0784); 
assign corrected[785] = (input_data[785]^invert0785); 
assign corrected[786] = (invert0786^input_data[786]); 
assign corrected[787] = (input_data[787]^invert0787); 
assign corrected[788] = (invert0788^input_data[788]); 
assign corrected[789] = (input_data[789]^invert0789); 
assign corrected[790] = (input_data[790]^invert0790); 
assign corrected[791] = (input_data[791]^invert0791); 
assign corrected[792] = (invert0792^input_data[792]); 
assign corrected[793] = (invert0793^input_data[793]); 
assign corrected[794] = (input_data[794]^invert0794); 
assign corrected[795] = (input_data[795]^invert0795); 
assign corrected[796] = (invert0796^input_data[796]); 
assign corrected[797] = (input_data[797]^invert0797); 
assign corrected[798] = (invert0798^input_data[798]); 
assign corrected[799] = (input_data[799]^invert0799); 
assign corrected[800] = (invert0800^input_data[800]); 
assign corrected[801] = (invert0801^input_data[801]); 
assign corrected[802] = (input_data[802]^invert0802); 
assign corrected[803] = (invert0803^input_data[803]); 
assign corrected[804] = (invert0804^input_data[804]); 
assign corrected[805] = (invert0805^input_data[805]); 
assign corrected[806] = (invert0806^input_data[806]); 
assign corrected[807] = (input_data[807]^invert0807); 
assign corrected[808] = (input_data[808]^invert0808); 
assign corrected[809] = (input_data[809]^invert0809); 
assign corrected[810] = (invert0810^input_data[810]); 
assign corrected[811] = (invert0811^input_data[811]); 
assign corrected[812] = (input_data[812]^invert0812); 
assign corrected[813] = (invert0813^input_data[813]); 
assign corrected[814] = (input_data[814]^invert0814); 
assign corrected[815] = (invert0815^input_data[815]); 
assign corrected[816] = (invert0816^input_data[816]); 
assign corrected[817] = (input_data[817]^invert0817); 
assign corrected[818] = (input_data[818]^invert0818); 
assign corrected[819] = (input_data[819]^invert0819); 
assign corrected[820] = (invert0820^input_data[820]); 
assign corrected[821] = (invert0821^input_data[821]); 
assign corrected[822] = (input_data[822]^invert0822); 
assign corrected[823] = (invert0823^input_data[823]); 
assign corrected[824] = (input_data[824]^invert0824); 
assign corrected[825] = (input_data[825]^invert0825); 
assign corrected[826] = (invert0826^input_data[826]); 
assign corrected[827] = (invert0827^input_data[827]); 
assign corrected[828] = (input_data[828]^invert0828); 
assign corrected[829] = (invert0829^input_data[829]); 
assign corrected[830] = (invert0830^input_data[830]); 
assign corrected[831] = (invert0831^input_data[831]); 
assign corrected[832] = (input_data[832]^invert0832); 
assign corrected[833] = (invert0833^input_data[833]); 
assign corrected[834] = (input_data[834]^invert0834); 
assign corrected[835] = (invert0835^input_data[835]); 
assign corrected[836] = (invert0836^input_data[836]); 
assign corrected[837] = (input_data[837]^invert0837); 
assign corrected[838] = (input_data[838]^invert0838); 
assign corrected[839] = (invert0839^input_data[839]); 
assign corrected[840] = (invert0840^input_data[840]); 
assign corrected[841] = (input_data[841]^invert0841); 
assign corrected[842] = (input_data[842]^invert0842); 
assign corrected[843] = (input_data[843]^invert0843); 
assign corrected[844] = (input_data[844]^invert0844); 
assign corrected[845] = (invert0845^input_data[845]); 
assign corrected[846] = (input_data[846]^invert0846); 
assign corrected[847] = (input_data[847]^invert0847); 
assign corrected[848] = (invert0848^input_data[848]); 
assign corrected[849] = (input_data[849]^invert0849); 
assign corrected[850] = (invert0850^input_data[850]); 
assign corrected[851] = (input_data[851]^invert0851); 
assign corrected[852] = (input_data[852]^invert0852); 
assign corrected[853] = (invert0853^input_data[853]); 
assign corrected[854] = (input_data[854]^invert0854); 
assign corrected[855] = (invert0855^input_data[855]); 
assign corrected[856] = (input_data[856]^invert0856); 
assign corrected[857] = (input_data[857]^invert0857); 
assign corrected[858] = (invert0858^input_data[858]); 
assign corrected[859] = (input_data[859]^invert0859); 
assign corrected[860] = (invert0860^input_data[860]); 
assign corrected[861] = (input_data[861]^invert0861); 
assign corrected[862] = (input_data[862]^invert0862); 
assign corrected[863] = (invert0863^input_data[863]); 
assign corrected[864] = (input_data[864]^invert0864); 
assign corrected[865] = (invert0865^input_data[865]); 
assign corrected[866] = (invert0866^input_data[866]); 
assign corrected[867] = (input_data[867]^invert0867); 
assign corrected[868] = (invert0868^input_data[868]); 
assign corrected[869] = (invert0869^input_data[869]); 
assign corrected[870] = (invert0870^input_data[870]); 
assign corrected[871] = (input_data[871]^invert0871); 
assign corrected[872] = (input_data[872]^invert0872); 
assign corrected[873] = (invert0873^input_data[873]); 
assign corrected[874] = (input_data[874]^invert0874); 
assign corrected[875] = (invert0875^input_data[875]); 
assign corrected[876] = (invert0876^input_data[876]); 
assign corrected[877] = (input_data[877]^invert0877); 
assign corrected[878] = (invert0878^input_data[878]); 
assign corrected[879] = (input_data[879]^invert0879); 
assign corrected[880] = (invert0880^input_data[880]); 
assign corrected[881] = (invert0881^input_data[881]); 
assign corrected[882] = (invert0882^input_data[882]); 
assign corrected[883] = (input_data[883]^invert0883); 
assign corrected[884] = (input_data[884]^invert0884); 
assign corrected[885] = (input_data[885]^invert0885); 
assign corrected[886] = (invert0886^input_data[886]); 
assign corrected[887] = (invert0887^input_data[887]); 
assign corrected[888] = (invert0888^input_data[888]); 
assign corrected[889] = (input_data[889]^invert0889); 
assign corrected[890] = (input_data[890]^invert0890); 
assign corrected[891] = (invert0891^input_data[891]); 
assign corrected[892] = (invert0892^input_data[892]); 
assign corrected[893] = (input_data[893]^invert0893); 
assign corrected[894] = (input_data[894]^invert0894); 
assign corrected[895] = (invert0895^input_data[895]); 
assign corrected[896] = (invert0896^input_data[896]); 
assign corrected[897] = (invert0897^input_data[897]); 
assign corrected[898] = (invert0898^input_data[898]); 
assign corrected[899] = (input_data[899]^invert0899); 
assign corrected[900] = (input_data[900]^invert0900); 
assign corrected[901] = (invert0901^input_data[901]); 
assign corrected[902] = (input_data[902]^invert0902); 
assign corrected[903] = (input_data[903]^invert0903); 
assign corrected[904] = (input_data[904]^invert0904); 
assign corrected[905] = (invert0905^input_data[905]); 
assign corrected[906] = (invert0906^input_data[906]); 
assign corrected[907] = (input_data[907]^invert0907); 
assign corrected[908] = (invert0908^input_data[908]); 
assign corrected[909] = (invert0909^input_data[909]); 
assign corrected[910] = (input_data[910]^invert0910); 
assign corrected[911] = (input_data[911]^invert0911); 
assign corrected[912] = (input_data[912]^invert0912); 
assign corrected[913] = (input_data[913]^invert0913); 
assign corrected[914] = (input_data[914]^invert0914); 
assign corrected[915] = (input_data[915]^invert0915); 
assign corrected[916] = (invert0916^input_data[916]); 
assign corrected[917] = (input_data[917]^invert0917); 
assign corrected[918] = (invert0918^input_data[918]); 
assign corrected[919] = (invert0919^input_data[919]); 
assign corrected[920] = (invert0920^input_data[920]); 
assign corrected[921] = (invert0921^input_data[921]); 
assign corrected[922] = (input_data[922]^invert0922); 
assign corrected[923] = (input_data[923]^invert0923); 
assign corrected[924] = (invert0924^input_data[924]); 
assign corrected[925] = (invert0925^input_data[925]); 
assign corrected[926] = (invert0926^input_data[926]); 
assign corrected[927] = (input_data[927]^invert0927); 
assign corrected[928] = (input_data[928]^invert0928); 
assign corrected[929] = (invert0929^input_data[929]); 
assign corrected[930] = (input_data[930]^invert0930); 
assign corrected[931] = (invert0931^input_data[931]); 
assign corrected[932] = (input_data[932]^invert0932); 
assign corrected[933] = (input_data[933]^invert0933); 
assign corrected[934] = (input_data[934]^invert0934); 
assign corrected[935] = (invert0935^input_data[935]); 
assign corrected[936] = (invert0936^input_data[936]); 
assign corrected[937] = (input_data[937]^invert0937); 
assign corrected[938] = (invert0938^input_data[938]); 
assign corrected[939] = (invert0939^input_data[939]); 
assign corrected[940] = (invert0940^input_data[940]); 
assign corrected[941] = (invert0941^input_data[941]); 
assign corrected[942] = (invert0942^input_data[942]); 
assign corrected[943] = (input_data[943]^invert0943); 
assign corrected[944] = (input_data[944]^invert0944); 
assign corrected[945] = (input_data[945]^invert0945); 
assign corrected[946] = (input_data[946]^invert0946); 
assign corrected[947] = (invert0947^input_data[947]); 
assign corrected[948] = (invert0948^input_data[948]); 
assign corrected[949] = (input_data[949]^invert0949); 
assign corrected[950] = (invert0950^input_data[950]); 
assign corrected[951] = (invert0951^input_data[951]); 
assign corrected[952] = (invert0952^input_data[952]); 
assign corrected[953] = (input_data[953]^invert0953); 
assign corrected[954] = (input_data[954]^invert0954); 
assign corrected[955] = (invert0955^input_data[955]); 
assign corrected[956] = (invert0956^input_data[956]); 
assign corrected[957] = (invert0957^input_data[957]); 
assign corrected[958] = (invert0958^input_data[958]); 
assign corrected[959] = (input_data[959]^invert0959); 
assign corrected[960] = (input_data[960]^invert0960); 
assign corrected[961] = (input_data[961]^invert0961); 
assign corrected[962] = (invert0962^input_data[962]); 
assign corrected[963] = (invert0963^input_data[963]); 
assign corrected[964] = (input_data[964]^invert0964); 
assign corrected[965] = (input_data[965]^invert0965); 
assign corrected[966] = (invert0966^input_data[966]); 
assign corrected[967] = (input_data[967]^invert0967); 
assign corrected[968] = (invert0968^input_data[968]); 
assign corrected[969] = (input_data[969]^invert0969); 
assign corrected[970] = (invert0970^input_data[970]); 
assign corrected[971] = (invert0971^input_data[971]); 
assign corrected[972] = (invert0972^input_data[972]); 
assign corrected[973] = (invert0973^input_data[973]); 
assign corrected[974] = (input_data[974]^invert0974); 
assign corrected[975] = (input_data[975]^invert0975); 
assign corrected[976] = (input_data[976]^invert0976); 
assign corrected[977] = (input_data[977]^invert0977); 
assign corrected[978] = (invert0978^input_data[978]); 
assign corrected[979] = (input_data[979]^invert0979); 
assign corrected[980] = (input_data[980]^invert0980); 
assign corrected[981] = (input_data[981]^invert0981); 
assign corrected[982] = (invert0982^input_data[982]); 
assign corrected[983] = (input_data[983]^invert0983); 
assign corrected[984] = (invert0984^input_data[984]); 
assign corrected[985] = (invert0985^input_data[985]); 
assign corrected[986] = (input_data[986]^invert0986); 
assign corrected[987] = (invert0987^input_data[987]); 
assign corrected[988] = (input_data[988]^invert0988); 
assign corrected[989] = (invert0989^input_data[989]); 
assign corrected[990] = (input_data[990]^invert0990); 
assign corrected[991] = (input_data[991]^invert0991); 
assign corrected[992] = (invert0992^input_data[992]); 
assign corrected[993] = (input_data[993]^invert0993); 
assign corrected[994] = (invert0994^input_data[994]); 
assign corrected[995] = (invert0995^input_data[995]); 
assign corrected[996] = (input_data[996]^invert0996); 
assign corrected[997] = (invert0997^input_data[997]); 
assign corrected[998] = (invert0998^input_data[998]); 
assign corrected[999] = (invert0999^input_data[999]); 
assign corrected[1000] = (invert1000^input_data[1000]); 
assign corrected[1001] = (input_data[1001]^invert1001); 
assign corrected[1002] = (invert1002^input_data[1002]); 
assign corrected[1003] = (invert1003^input_data[1003]); 
assign corrected[1004] = (input_data[1004]^invert1004); 
assign corrected[1005] = (input_data[1005]^invert1005); 
assign corrected[1006] = (invert1006^input_data[1006]); 
assign corrected[1007] = (input_data[1007]^invert1007); 
assign corrected[1008] = (input_data[1008]^invert1008); 
assign corrected[1009] = (invert1009^input_data[1009]); 
assign corrected[1010] = (invert1010^input_data[1010]); 
assign corrected[1011] = (input_data[1011]^invert1011); 
assign corrected[1012] = (invert1012^input_data[1012]); 
assign corrected[1013] = (invert1013^input_data[1013]); 
assign corrected[1014] = (input_data[1014]^invert1014); 
assign corrected[1015] = (input_data[1015]^invert1015); 
assign corrected[1016] = (invert1016^input_data[1016]); 
assign corrected[1017] = (input_data[1017]^invert1017); 
assign corrected[1018] = (invert1018^input_data[1018]); 
assign corrected[1019] = (input_data[1019]^invert1019); 
assign corrected[1020] = (input_data[1020]^invert1020); 
assign corrected[1021] = (invert1021^input_data[1021]); 
assign corrected[1022] = (input_data[1022]^invert1022); 
assign corrected[1023] = (invert1023^input_data[1023]); 
assign o_err_detect = |(ecc_parity[10-1:-1]);
assign o_err_multpl = o_err_detect & !ecc_parity[-1];
endmodule
