magic
tech scmos
timestamp 988943070
<< nselect >>
rect -33 27 0 90
<< pselect >>
rect 0 18 46 98
<< ndiffusion >>
rect -28 76 -8 77
rect -28 68 -8 73
rect -28 60 -8 65
rect -28 52 -8 57
rect -28 44 -8 49
rect -28 40 -8 41
<< pdiffusion >>
rect 8 86 40 87
rect 8 82 40 83
rect 28 74 40 82
rect 8 73 40 74
rect 8 69 40 70
rect 8 60 40 61
rect 8 56 40 57
rect 28 48 40 56
rect 8 47 40 48
rect 8 43 40 44
rect 8 32 40 35
rect 8 28 40 29
<< ntransistor >>
rect -28 73 -8 76
rect -28 65 -8 68
rect -28 57 -8 60
rect -28 49 -8 52
rect -28 41 -8 44
<< ptransistor >>
rect 8 83 40 86
rect 8 70 40 73
rect 8 57 40 60
rect 8 44 40 47
rect 8 29 40 32
<< polysilicon >>
rect -6 83 8 86
rect 40 83 44 86
rect -6 76 -3 83
rect -32 73 -28 76
rect -8 73 -3 76
rect 3 70 8 73
rect 40 70 44 73
rect 3 68 6 70
rect -32 65 -28 68
rect -8 65 6 68
rect -32 57 -28 60
rect -8 57 8 60
rect 40 57 44 60
rect -32 49 -28 52
rect -8 49 6 52
rect 3 47 6 49
rect 3 44 8 47
rect 40 44 44 47
rect -32 41 -28 44
rect -8 41 -4 44
rect 4 29 8 32
rect 40 29 44 32
<< ndcontact >>
rect -28 77 -8 85
rect -28 32 -8 40
<< pdcontact >>
rect 8 87 40 95
rect 8 74 28 82
rect 8 61 40 69
rect 8 48 28 56
rect 8 35 40 43
rect 8 20 40 28
<< metal1 >>
rect 8 87 40 95
rect -28 82 -8 85
rect -28 77 28 82
rect -4 74 28 77
rect -4 56 4 74
rect 32 69 40 87
rect 8 61 40 69
rect -4 48 28 56
rect -28 32 -8 40
rect -4 28 4 48
rect 32 43 40 61
rect 8 35 40 43
rect -4 20 40 28
<< labels >>
rlabel space 28 39 47 98 3 ^p
rlabel space -33 26 -28 91 7 ^n
rlabel metal1 8 61 40 69 1 Vdd!|pin|s|1
rlabel metal1 -4 20 4 82 1 x|pin|s|2
rlabel metal1 -28 77 -8 85 1 x|pin|s|2
rlabel metal1 8 74 28 82 1 x|pin|s|2
rlabel metal1 8 48 28 56 1 x|pin|s|2
rlabel metal1 -4 20 40 28 1 x|pin|s|2
rlabel polysilicon 40 44 44 47 1 a|pin|w|3|poly
rlabel polysilicon 3 44 7 47 1 a|pin|w|3|poly
rlabel polysilicon -32 49 -28 52 1 a|pin|w|3|poly
rlabel polysilicon 40 57 44 60 1 b|pin|w|4|poly
rlabel polysilicon -32 57 -28 60 1 b|pin|w|4|poly
rlabel polysilicon 40 70 44 73 1 c|pin|w|5|poly
rlabel polysilicon -32 65 -28 68 1 c|pin|w|5|poly
rlabel polysilicon 40 83 44 86 1 d|pin|w|6|poly
rlabel polysilicon -2 83 2 86 1 d|pin|w|6|poly
rlabel polysilicon -32 73 -28 76 1 d|pin|w|6|poly
rlabel polysilicon -32 41 -28 44 1 _SReset!|pin|w|7|poly
rlabel polysilicon -8 41 -4 44 1 _SReset!|pin|w|7|poly
rlabel polysilicon 4 29 8 32 1 _PReset!|pin|w|8|poly
rlabel polysilicon 40 29 44 32 1 _PReset!|pin|w|8|poly
rlabel metal1 32 43 40 95 1 Vdd!|pin|s|1
rlabel metal1 -28 32 -8 40 1 GND!|pin|s|0
rlabel metal1 8 87 40 95 1 Vdd!|pin|s|1
rlabel metal1 8 35 40 43 1 Vdd!|pin|s|1
<< end >>
