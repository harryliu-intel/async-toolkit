magic
tech scmos
timestamp 988943070
<< nselect >>
rect -87 -181 0 -110
<< pselect >>
rect 0 -181 93 -116
<< ndiffusion >>
rect -57 -122 -49 -121
rect -57 -130 -49 -125
rect -28 -130 -8 -129
rect -57 -138 -49 -133
rect -28 -138 -8 -133
rect -57 -142 -49 -141
rect -57 -151 -49 -150
rect -28 -142 -8 -141
rect -81 -159 -73 -158
rect -57 -159 -49 -154
rect -28 -151 -8 -150
rect -28 -159 -8 -154
rect -81 -163 -73 -162
rect -57 -167 -49 -162
rect -28 -163 -8 -162
rect -57 -171 -49 -170
<< pdiffusion >>
rect 8 -130 28 -129
rect 49 -130 61 -129
rect 75 -130 87 -129
rect 8 -138 28 -133
rect 8 -142 28 -141
rect 49 -138 61 -133
rect 75 -134 87 -133
rect 8 -151 28 -150
rect 49 -142 61 -141
rect 49 -151 61 -150
rect 83 -139 87 -134
rect 8 -159 28 -154
rect 49 -159 61 -154
rect 8 -163 28 -162
rect 49 -163 61 -162
rect 67 -166 79 -161
rect 67 -167 87 -166
rect 67 -171 87 -170
<< ntransistor >>
rect -57 -125 -49 -122
rect -57 -133 -49 -130
rect -28 -133 -8 -130
rect -57 -141 -49 -138
rect -28 -141 -8 -138
rect -57 -154 -49 -151
rect -28 -154 -8 -151
rect -81 -162 -73 -159
rect -57 -162 -49 -159
rect -28 -162 -8 -159
rect -57 -170 -49 -167
<< ptransistor >>
rect 8 -133 28 -130
rect 49 -133 61 -130
rect 75 -133 87 -130
rect 8 -141 28 -138
rect 49 -141 61 -138
rect 8 -154 28 -151
rect 49 -154 61 -151
rect 8 -162 28 -159
rect 49 -162 61 -159
rect 67 -170 87 -167
<< polysilicon >>
rect -61 -125 -57 -122
rect -49 -125 -45 -122
rect -61 -133 -57 -130
rect -49 -133 -28 -130
rect -8 -133 8 -130
rect 28 -133 49 -130
rect 61 -133 65 -130
rect 71 -133 75 -130
rect 87 -133 92 -130
rect -86 -146 -82 -143
rect -62 -141 -57 -138
rect -49 -141 -45 -138
rect -62 -146 -59 -141
rect -86 -159 -83 -146
rect -61 -151 -59 -146
rect -32 -141 -28 -138
rect -8 -141 8 -138
rect 28 -141 32 -138
rect -61 -154 -57 -151
rect -49 -154 -45 -151
rect -40 -159 -37 -146
rect 37 -146 40 -133
rect 45 -141 49 -138
rect 61 -141 65 -138
rect -32 -154 -28 -151
rect -8 -154 8 -151
rect 28 -154 32 -151
rect 63 -146 65 -141
rect 89 -146 92 -133
rect 63 -151 66 -146
rect 45 -154 49 -151
rect 61 -154 66 -151
rect 87 -149 92 -146
rect -86 -162 -81 -159
rect -73 -162 -69 -159
rect -61 -162 -57 -159
rect -49 -162 -28 -159
rect -8 -162 8 -159
rect 28 -162 49 -159
rect 61 -162 65 -159
rect -61 -170 -57 -167
rect -49 -170 -45 -167
rect 63 -170 67 -167
rect 87 -170 91 -167
<< ndcontact >>
rect -57 -121 -49 -113
rect -28 -129 -8 -121
rect -81 -158 -73 -150
rect -57 -150 -49 -142
rect -28 -150 -8 -142
rect -81 -171 -73 -163
rect -28 -171 -8 -163
rect -57 -179 -49 -171
<< pdcontact >>
rect 8 -129 28 -121
rect 49 -129 61 -121
rect 75 -129 87 -121
rect 8 -150 28 -142
rect 49 -150 61 -142
rect 75 -142 83 -134
rect 8 -171 28 -163
rect 49 -171 61 -163
rect 79 -166 87 -158
rect 67 -179 87 -171
<< polycontact >>
rect -82 -146 -74 -138
rect -69 -154 -61 -146
rect -40 -146 -32 -138
rect 32 -154 40 -146
rect 65 -146 73 -138
rect 79 -154 87 -146
<< metal1 >>
rect -57 -121 -8 -113
rect -28 -129 -8 -121
rect 8 -129 87 -121
rect -2 -138 83 -134
rect -82 -142 -53 -138
rect -82 -146 -74 -142
rect -69 -150 -61 -146
rect -57 -150 -49 -142
rect -40 -146 -32 -138
rect -28 -150 -8 -142
rect -81 -154 -61 -150
rect -2 -154 2 -138
rect 65 -142 83 -138
rect 8 -150 28 -142
rect 32 -154 40 -146
rect 49 -150 61 -142
rect 65 -146 73 -142
rect 79 -150 87 -146
rect 57 -154 87 -150
rect -81 -158 2 -154
rect -81 -167 -52 -163
rect -81 -171 -73 -167
rect -57 -171 -52 -167
rect -28 -171 -8 -163
rect 8 -171 74 -163
rect 79 -166 87 -154
rect -57 -179 -8 -171
rect 67 -179 87 -171
<< labels >>
rlabel metal1 32 -154 40 -146 1 b
rlabel metal1 -40 -146 -32 -138 1 a
rlabel space -88 -181 -28 -110 7 ^n
rlabel space 28 -181 94 -116 3 ^p
rlabel metal1 -81 -171 -73 -163 1 GND!|pin|s|0
rlabel metal1 -28 -171 -8 -163 1 GND!|pin|s|0
rlabel metal1 8 -171 74 -163 1 Vdd!|pin|s|1
rlabel metal1 67 -179 87 -171 1 Vdd!|pin|s|1
rlabel polysilicon -61 -170 -57 -167 1 _SReset!|pin|w|3|poly
rlabel polysilicon -49 -170 -45 -167 1 _SReset!|pin|w|3|poly
rlabel polysilicon -61 -125 -57 -122 1 _SReset!|pin|w|4|poly
rlabel polysilicon -49 -125 -45 -122 1 _SReset!|pin|w|4|poly
rlabel polysilicon 87 -170 91 -167 1 _PReset!|pin|w|5|poly
rlabel metal1 8 -129 87 -121 1 Vdd!|pin|s|2
rlabel metal1 -28 -129 -8 -121 1 GND!|pin|s|1
rlabel metal1 -57 -121 -8 -113 1 GND!|pin|s|1
rlabel metal1 -82 -142 -53 -138 1 x|pin|s|0
rlabel metal1 -57 -150 -49 -142 1 x|pin|s|0
rlabel metal1 -28 -150 -8 -142 1 x|pin|s|1
rlabel metal1 8 -150 28 -142 1 x|pin|s|2
rlabel metal1 49 -150 61 -142 1 x|pin|s|3
rlabel metal1 57 -154 87 -150 1 x|pin|s|3
rlabel metal1 79 -154 87 -146 1 x|pin|s|3
rlabel metal1 -82 -146 -74 -138 1 x|pin|s|0
rlabel metal1 -57 -179 -8 -171 1 GND!|pin|s|0
<< end >>
