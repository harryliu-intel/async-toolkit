// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

///
///  INTEL CONFIDENTIAL
///
///  Copyright 2019 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_rx_pb_pkg.vh                                           
// Creator:         ggomezde                                                   
// Time:            Wednesday Jan 30, 2019 [10:27:46 am]                       
//                                                                             
// Path:            /tmp/ggomezde/nebulon_run/2768731022_2019-01-30.10:27:12   
// Arguments:       -I                                                         
//                  /nfs/site/disks/sc_mby_00088/ggomezde/mby/work_root/models/mby_ww05_ral_TI/tools/srdl
//                  -sv_no_sai_checks -sverilog -crif -expand_handcoded_arrays 
//                  -maximize_crif -input mby_rx_pb_map.rdl -timeout 60000     
//                  -out_dir /tmp/tmp.C8ZQyTQrjK -log_file                     
//                  /nfs/site/disks/sc_mby_00088/ggomezde/mby/work_root/models/mby_ww05_ral_TI/target/GenRTL/regflow/mby/subblock/mby_rx_pb_map_crif.xml.log
//                                                                             
// MRE:             5.2018.3.p1                                                
// Machine:         sccj004303                                                 
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww52.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2019 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtlgen_pkg_template

`ifndef MBY_RX_PB_PKG_VH
`define MBY_RX_PB_PKG_VH

`include "rtlgen_include_mby_rx_pb_map.vh"
`include "rtlgen_pkg_mby_rx_pb_map.vh"

package mby_rx_pb_pkg;

import rtlgen_pkg_mby_rx_pb_map::*;

typedef cfg_req_64bit_t mby_rx_pb_cr_req_t;
typedef cfg_ack_64bit_t mby_rx_pb_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_rx_pb_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic [31:0] PORT;  // RW
} RX_PB_PORT_CFG_t;

localparam RX_PB_PORT_CFG_REG_STRIDE = 48'h8;
localparam RX_PB_PORT_CFG_REG_ENTRIES = 1;
localparam [47:0] RX_PB_PORT_CFG_CR_ADDR = 48'h0;
localparam RX_PB_PORT_CFG_SIZE = 64;
localparam RX_PB_PORT_CFG_PORT_LO = 0;
localparam RX_PB_PORT_CFG_PORT_HI = 31;
localparam RX_PB_PORT_CFG_PORT_RESET = 32'h0;
localparam RX_PB_PORT_CFG_USEMASK = 64'hFFFFFFFF;
localparam RX_PB_PORT_CFG_RO_MASK = 64'h0;
localparam RX_PB_PORT_CFG_WO_MASK = 64'h0;
localparam RX_PB_PORT_CFG_RESET = 64'h0;

typedef struct packed {
    logic [42:0] reserved0;  // RSVD
    logic  [0:0] LOSSLESS;  // RW
    logic  [9:0] XON;  // RW
    logic  [9:0] XOFF_OR_DROP;  // RW
} RX_PB_WM_t;

localparam RX_PB_WM_REG_STRIDE = 48'h8;
localparam RX_PB_WM_REG_ENTRIES = 8;
localparam RX_PB_WM_REGFILE_STRIDE = 48'h40;
localparam RX_PB_WM_REGFILE_ENTRIES = 17;
localparam [16:0][7:0][47:0] RX_PB_WM_CR_ADDR = {{48'hC38, 48'hC30, 48'hC28, 48'hC20, 48'hC18, 48'hC10, 48'hC08, 48'hC00}, {48'hBF8, 48'hBF0, 48'hBE8, 48'hBE0, 48'hBD8, 48'hBD0, 48'hBC8, 48'hBC0}, {48'hBB8, 48'hBB0, 48'hBA8, 48'hBA0, 48'hB98, 48'hB90, 48'hB88, 48'hB80}, {48'hB78, 48'hB70, 48'hB68, 48'hB60, 48'hB58, 48'hB50, 48'hB48, 48'hB40}, {48'hB38, 48'hB30, 48'hB28, 48'hB20, 48'hB18, 48'hB10, 48'hB08, 48'hB00}, {48'hAF8, 48'hAF0, 48'hAE8, 48'hAE0, 48'hAD8, 48'hAD0, 48'hAC8, 48'hAC0}, {48'hAB8, 48'hAB0, 48'hAA8, 48'hAA0, 48'hA98, 48'hA90, 48'hA88, 48'hA80}, {48'hA78, 48'hA70, 48'hA68, 48'hA60, 48'hA58, 48'hA50, 48'hA48, 48'hA40}, {48'hA38, 48'hA30, 48'hA28, 48'hA20, 48'hA18, 48'hA10, 48'hA08, 48'hA00}, {48'h9F8, 48'h9F0, 48'h9E8, 48'h9E0, 48'h9D8, 48'h9D0, 48'h9C8, 48'h9C0}, {48'h9B8, 48'h9B0, 48'h9A8, 48'h9A0, 48'h998, 48'h990, 48'h988, 48'h980}, {48'h978, 48'h970, 48'h968, 48'h960, 48'h958, 48'h950, 48'h948, 48'h940}, {48'h938, 48'h930, 48'h928, 48'h920, 48'h918, 48'h910, 48'h908, 48'h900}, {48'h8F8, 48'h8F0, 48'h8E8, 48'h8E0, 48'h8D8, 48'h8D0, 48'h8C8, 48'h8C0}, {48'h8B8, 48'h8B0, 48'h8A8, 48'h8A0, 48'h898, 48'h890, 48'h888, 48'h880}, {48'h878, 48'h870, 48'h868, 48'h860, 48'h858, 48'h850, 48'h848, 48'h840}, {48'h838, 48'h830, 48'h828, 48'h820, 48'h818, 48'h810, 48'h808, 48'h800}};
localparam RX_PB_WM_SIZE = 64;
localparam RX_PB_WM_LOSSLESS_LO = 20;
localparam RX_PB_WM_LOSSLESS_HI = 20;
localparam RX_PB_WM_LOSSLESS_RESET = 'h0;
localparam RX_PB_WM_XON_LO = 10;
localparam RX_PB_WM_XON_HI = 19;
localparam RX_PB_WM_XON_RESET = 'h200;
localparam RX_PB_WM_XOFF_OR_DROP_LO = 0;
localparam RX_PB_WM_XOFF_OR_DROP_HI = 9;
localparam RX_PB_WM_XOFF_OR_DROP_RESET = 'h200;
localparam RX_PB_WM_USEMASK = 64'h1FFFFF;
localparam RX_PB_WM_RO_MASK = 64'h0;
localparam RX_PB_WM_WO_MASK = 64'h0;
localparam RX_PB_WM_RESET = 64'h80200;

typedef struct packed {
    RX_PB_PORT_CFG_t  RX_PB_PORT_CFG;
    RX_PB_WM_t [16:0][7:0] RX_PB_WM;
} mby_rx_pb_registers_t;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// RW/V2 Structure

// ===================================================
// Parity Bit Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_rx_pb_pkg

`endif // MBY_RX_PB_PKG_VH
