///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cgrp_a_nested_map_pkg.vh                           
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_CGRP_A_NESTED_MAP_PKG_VH
`define MBY_PPE_CGRP_A_NESTED_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_cgrp_a_nested_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_cgrp_a_nested_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_cgrp_a_nested_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_cgrp_a_nested_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [43:0] reserved0;  // RSVD
    logic [19:0] PTR;  // RW
    logic [11:0] reserved1;  // RSVD
    logic  [3:0] SELECT_4;  // RW
    logic  [3:0] SELECT_3;  // RW
    logic  [3:0] SELECT_2;  // RW
    logic  [3:0] SELECT_1;  // RW
    logic  [3:0] SELECT_0;  // RW
    logic [31:0] MASK;  // RW
} EM_HASH_LOOKUP_t;

localparam EM_HASH_LOOKUP_REG_STRIDE = 48'h10;
localparam EM_HASH_LOOKUP_REG_ENTRIES = 32768;
localparam EM_HASH_LOOKUP_CR_ADDR = 48'h0;
localparam EM_HASH_LOOKUP_SIZE = 128;
localparam EM_HASH_LOOKUP_PTR_LO = 64;
localparam EM_HASH_LOOKUP_PTR_HI = 83;
localparam EM_HASH_LOOKUP_PTR_RESET = 20'h0;
localparam EM_HASH_LOOKUP_SELECT_4_LO = 48;
localparam EM_HASH_LOOKUP_SELECT_4_HI = 51;
localparam EM_HASH_LOOKUP_SELECT_4_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_3_LO = 44;
localparam EM_HASH_LOOKUP_SELECT_3_HI = 47;
localparam EM_HASH_LOOKUP_SELECT_3_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_2_LO = 40;
localparam EM_HASH_LOOKUP_SELECT_2_HI = 43;
localparam EM_HASH_LOOKUP_SELECT_2_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_1_LO = 36;
localparam EM_HASH_LOOKUP_SELECT_1_HI = 39;
localparam EM_HASH_LOOKUP_SELECT_1_RESET = 4'h0;
localparam EM_HASH_LOOKUP_SELECT_0_LO = 32;
localparam EM_HASH_LOOKUP_SELECT_0_HI = 35;
localparam EM_HASH_LOOKUP_SELECT_0_RESET = 4'h0;
localparam EM_HASH_LOOKUP_MASK_LO = 0;
localparam EM_HASH_LOOKUP_MASK_HI = 31;
localparam EM_HASH_LOOKUP_MASK_RESET = 32'h0;
localparam EM_HASH_LOOKUP_USEMASK = 128'hFFFFF000FFFFFFFFFFFFF;
localparam EM_HASH_LOOKUP_RO_MASK = 128'h0;
localparam EM_HASH_LOOKUP_WO_MASK = 128'h0;
localparam EM_HASH_LOOKUP_RESET = 128'h0;

typedef struct packed {
    logic [44:0] reserved0;  // RSVD
    logic [18:0] ACTION_BASE_PTR;  // RW
} LPM_SUBTRIE_APTR_t;

localparam LPM_SUBTRIE_APTR_REG_STRIDE = 48'h8;
localparam LPM_SUBTRIE_APTR_REG_ENTRIES = 512;
localparam LPM_SUBTRIE_APTR_REGFILE_STRIDE = 48'h1000;
localparam LPM_SUBTRIE_APTR_REGFILE_ENTRIES = 48;
localparam LPM_SUBTRIE_APTR_CR_ADDR = 48'h80000;
localparam LPM_SUBTRIE_APTR_SIZE = 64;
localparam LPM_SUBTRIE_APTR_ACTION_BASE_PTR_LO = 0;
localparam LPM_SUBTRIE_APTR_ACTION_BASE_PTR_HI = 18;
localparam LPM_SUBTRIE_APTR_ACTION_BASE_PTR_RESET = 19'h0;
localparam LPM_SUBTRIE_APTR_USEMASK = 64'h7FFFF;
localparam LPM_SUBTRIE_APTR_RO_MASK = 64'h0;
localparam LPM_SUBTRIE_APTR_WO_MASK = 64'h0;
localparam LPM_SUBTRIE_APTR_RESET = 64'h0;

typedef struct packed {
    logic [23:0] reserved0;  // RSVD
    logic  [7:0] CHILD_PTR_LEN;  // RW
    logic [15:0] CHILD_BASE_PTR;  // RW
    logic [15:0] SUBTRIE_PTR;  // RW
} LPM_SUBTRIE_CPTR_t;

localparam LPM_SUBTRIE_CPTR_REG_STRIDE = 48'h8;
localparam LPM_SUBTRIE_CPTR_REG_ENTRIES = 512;
localparam LPM_SUBTRIE_CPTR_REGFILE_STRIDE = 48'h1000;
localparam LPM_SUBTRIE_CPTR_REGFILE_ENTRIES = 48;
localparam LPM_SUBTRIE_CPTR_CR_ADDR = 48'hC0000;
localparam LPM_SUBTRIE_CPTR_SIZE = 64;
localparam LPM_SUBTRIE_CPTR_CHILD_PTR_LEN_LO = 32;
localparam LPM_SUBTRIE_CPTR_CHILD_PTR_LEN_HI = 39;
localparam LPM_SUBTRIE_CPTR_CHILD_PTR_LEN_RESET = 8'h0;
localparam LPM_SUBTRIE_CPTR_CHILD_BASE_PTR_LO = 16;
localparam LPM_SUBTRIE_CPTR_CHILD_BASE_PTR_HI = 31;
localparam LPM_SUBTRIE_CPTR_CHILD_BASE_PTR_RESET = 16'h0;
localparam LPM_SUBTRIE_CPTR_SUBTRIE_PTR_LO = 0;
localparam LPM_SUBTRIE_CPTR_SUBTRIE_PTR_HI = 15;
localparam LPM_SUBTRIE_CPTR_SUBTRIE_PTR_RESET = 16'h0;
localparam LPM_SUBTRIE_CPTR_USEMASK = 64'hFFFFFFFFFF;
localparam LPM_SUBTRIE_CPTR_RO_MASK = 64'h0;
localparam LPM_SUBTRIE_CPTR_WO_MASK = 64'h0;
localparam LPM_SUBTRIE_CPTR_RESET = 64'h0;

typedef struct packed {
    logic [63:0] BITMAP;  // RW
} LPM_SUBTRIE_BITMAPS_t;

localparam LPM_SUBTRIE_BITMAPS_REG_STRIDE = 48'h8;
localparam LPM_SUBTRIE_BITMAPS_REG_ENTRIES = 4096;
localparam LPM_SUBTRIE_BITMAPS_REGFILE_STRIDE = 48'h8000;
localparam LPM_SUBTRIE_BITMAPS_REGFILE_ENTRIES = 48;
localparam LPM_SUBTRIE_BITMAPS_CR_ADDR = 48'h200000;
localparam LPM_SUBTRIE_BITMAPS_SIZE = 64;
localparam LPM_SUBTRIE_BITMAPS_BITMAP_LO = 0;
localparam LPM_SUBTRIE_BITMAPS_BITMAP_HI = 63;
localparam LPM_SUBTRIE_BITMAPS_BITMAP_RESET = 64'h0;
localparam LPM_SUBTRIE_BITMAPS_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam LPM_SUBTRIE_BITMAPS_RO_MASK = 64'h0;
localparam LPM_SUBTRIE_BITMAPS_WO_MASK = 64'h0;
localparam LPM_SUBTRIE_BITMAPS_RESET = 64'h0;

typedef struct packed {
    logic [31:0] KEY_INVERT;  // RW
    logic [31:0] KEY;  // RW
} LPM_MATCH_TCAM_t;

localparam LPM_MATCH_TCAM_REG_STRIDE = 48'h8;
localparam LPM_MATCH_TCAM_REG_ENTRIES = 512;
localparam LPM_MATCH_TCAM_CR_ADDR = 48'h380000;
localparam LPM_MATCH_TCAM_SIZE = 64;
localparam LPM_MATCH_TCAM_KEY_INVERT_LO = 32;
localparam LPM_MATCH_TCAM_KEY_INVERT_HI = 63;
localparam LPM_MATCH_TCAM_KEY_INVERT_RESET = 32'h0;
localparam LPM_MATCH_TCAM_KEY_LO = 0;
localparam LPM_MATCH_TCAM_KEY_HI = 31;
localparam LPM_MATCH_TCAM_KEY_RESET = 32'h0;
localparam LPM_MATCH_TCAM_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam LPM_MATCH_TCAM_RO_MASK = 64'h0;
localparam LPM_MATCH_TCAM_WO_MASK = 64'h0;
localparam LPM_MATCH_TCAM_RESET = 64'h0;

typedef struct packed {
    logic [23:0] reserved0;  // RSVD
    logic  [7:0] CHILD_PTR_LEN;  // RW
    logic [15:0] CHILD_BASE_PTR;  // RW
    logic [15:0] ROOT_PTR;  // RW
} LPM_MATCH_ACTION_t;

localparam LPM_MATCH_ACTION_REG_STRIDE = 48'h8;
localparam LPM_MATCH_ACTION_REG_ENTRIES = 512;
localparam LPM_MATCH_ACTION_CR_ADDR = 48'h381000;
localparam LPM_MATCH_ACTION_SIZE = 64;
localparam LPM_MATCH_ACTION_CHILD_PTR_LEN_LO = 32;
localparam LPM_MATCH_ACTION_CHILD_PTR_LEN_HI = 39;
localparam LPM_MATCH_ACTION_CHILD_PTR_LEN_RESET = 8'h0;
localparam LPM_MATCH_ACTION_CHILD_BASE_PTR_LO = 16;
localparam LPM_MATCH_ACTION_CHILD_BASE_PTR_HI = 31;
localparam LPM_MATCH_ACTION_CHILD_BASE_PTR_RESET = 16'h0;
localparam LPM_MATCH_ACTION_ROOT_PTR_LO = 0;
localparam LPM_MATCH_ACTION_ROOT_PTR_HI = 15;
localparam LPM_MATCH_ACTION_ROOT_PTR_RESET = 16'h0;
localparam LPM_MATCH_ACTION_USEMASK = 64'hFFFFFFFFFF;
localparam LPM_MATCH_ACTION_RO_MASK = 64'h0;
localparam LPM_MATCH_ACTION_WO_MASK = 64'h0;
localparam LPM_MATCH_ACTION_RESET = 64'h0;

typedef struct packed {
    logic [63:0] MASK;  // RW
} LPM_KEY_MASK_t;

localparam LPM_KEY_MASK_REG_STRIDE = 48'h8;
localparam LPM_KEY_MASK_REG_ENTRIES = 20;
localparam LPM_KEY_MASK_REGFILE_STRIDE = 48'h100;
localparam LPM_KEY_MASK_REGFILE_ENTRIES = 64;
localparam LPM_KEY_MASK_CR_ADDR = 48'h384000;
localparam LPM_KEY_MASK_SIZE = 64;
localparam LPM_KEY_MASK_MASK_LO = 0;
localparam LPM_KEY_MASK_MASK_HI = 63;
localparam LPM_KEY_MASK_MASK_RESET = 64'h0;
localparam LPM_KEY_MASK_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam LPM_KEY_MASK_RO_MASK = 64'h0;
localparam LPM_KEY_MASK_WO_MASK = 64'h0;
localparam LPM_KEY_MASK_RESET = 64'h0;

typedef struct packed {
    logic [63:0] MD_KEY16_SEL;  // RW
} LPM_KEY_SEL0_t;

localparam LPM_KEY_SEL0_REG_STRIDE = 48'h8;
localparam LPM_KEY_SEL0_REG_ENTRIES = 64;
localparam LPM_KEY_SEL0_CR_ADDR = 48'h388000;
localparam LPM_KEY_SEL0_SIZE = 64;
localparam LPM_KEY_SEL0_MD_KEY16_SEL_LO = 0;
localparam LPM_KEY_SEL0_MD_KEY16_SEL_HI = 63;
localparam LPM_KEY_SEL0_MD_KEY16_SEL_RESET = 64'h0;
localparam LPM_KEY_SEL0_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam LPM_KEY_SEL0_RO_MASK = 64'h0;
localparam LPM_KEY_SEL0_WO_MASK = 64'h0;
localparam LPM_KEY_SEL0_RESET = 64'h0;

typedef struct packed {
    logic [31:0] ADDR_KEY8_SEL;  // RW
    logic [31:0] MD_KEY8_SEL;  // RW
} LPM_KEY_SEL1_t;

localparam LPM_KEY_SEL1_REG_STRIDE = 48'h8;
localparam LPM_KEY_SEL1_REG_ENTRIES = 64;
localparam LPM_KEY_SEL1_CR_ADDR = 48'h388200;
localparam LPM_KEY_SEL1_SIZE = 64;
localparam LPM_KEY_SEL1_ADDR_KEY8_SEL_LO = 32;
localparam LPM_KEY_SEL1_ADDR_KEY8_SEL_HI = 63;
localparam LPM_KEY_SEL1_ADDR_KEY8_SEL_RESET = 32'h0;
localparam LPM_KEY_SEL1_MD_KEY8_SEL_LO = 0;
localparam LPM_KEY_SEL1_MD_KEY8_SEL_HI = 31;
localparam LPM_KEY_SEL1_MD_KEY8_SEL_RESET = 32'h0;
localparam LPM_KEY_SEL1_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam LPM_KEY_SEL1_RO_MASK = 64'h0;
localparam LPM_KEY_SEL1_WO_MASK = 64'h0;
localparam LPM_KEY_SEL1_RESET = 64'h0;

typedef struct packed {
    logic [63:0] ADDR_KEY16_SEL;  // RW
} LPM_KEY_SEL2_t;

localparam LPM_KEY_SEL2_REG_STRIDE = 48'h8;
localparam LPM_KEY_SEL2_REG_ENTRIES = 64;
localparam LPM_KEY_SEL2_CR_ADDR = 48'h388400;
localparam LPM_KEY_SEL2_SIZE = 64;
localparam LPM_KEY_SEL2_ADDR_KEY16_SEL_LO = 0;
localparam LPM_KEY_SEL2_ADDR_KEY16_SEL_HI = 63;
localparam LPM_KEY_SEL2_ADDR_KEY16_SEL_RESET = 64'h0;
localparam LPM_KEY_SEL2_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam LPM_KEY_SEL2_RO_MASK = 64'h0;
localparam LPM_KEY_SEL2_WO_MASK = 64'h0;
localparam LPM_KEY_SEL2_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] ADDR_KEY32_SEL;  // RW
} LPM_KEY_SEL3_t;

localparam LPM_KEY_SEL3_REG_STRIDE = 48'h8;
localparam LPM_KEY_SEL3_REG_ENTRIES = 64;
localparam LPM_KEY_SEL3_CR_ADDR = 48'h388600;
localparam LPM_KEY_SEL3_SIZE = 64;
localparam LPM_KEY_SEL3_ADDR_KEY32_SEL_LO = 0;
localparam LPM_KEY_SEL3_ADDR_KEY32_SEL_HI = 15;
localparam LPM_KEY_SEL3_ADDR_KEY32_SEL_RESET = 16'h0;
localparam LPM_KEY_SEL3_USEMASK = 64'hFFFF;
localparam LPM_KEY_SEL3_RO_MASK = 64'h0;
localparam LPM_KEY_SEL3_WO_MASK = 64'h0;
localparam LPM_KEY_SEL3_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [15:0] we_EM_HASH_LOOKUP_t;

typedef logic [7:0] we_LPM_SUBTRIE_APTR_t;

typedef logic [7:0] we_LPM_SUBTRIE_CPTR_t;

typedef logic [7:0] we_LPM_SUBTRIE_BITMAPS_t;

typedef logic [7:0] we_LPM_MATCH_TCAM_t;

typedef logic [7:0] we_LPM_MATCH_ACTION_t;

typedef logic [7:0] we_LPM_KEY_MASK_t;

typedef logic [7:0] we_LPM_KEY_SEL0_t;

typedef logic [7:0] we_LPM_KEY_SEL1_t;

typedef logic [7:0] we_LPM_KEY_SEL2_t;

typedef logic [7:0] we_LPM_KEY_SEL3_t;

typedef struct packed {
    we_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    we_LPM_SUBTRIE_APTR_t LPM_SUBTRIE_APTR;
    we_LPM_SUBTRIE_CPTR_t LPM_SUBTRIE_CPTR;
    we_LPM_SUBTRIE_BITMAPS_t LPM_SUBTRIE_BITMAPS;
    we_LPM_MATCH_TCAM_t LPM_MATCH_TCAM;
    we_LPM_MATCH_ACTION_t LPM_MATCH_ACTION;
    we_LPM_KEY_MASK_t LPM_KEY_MASK;
    we_LPM_KEY_SEL0_t LPM_KEY_SEL0;
    we_LPM_KEY_SEL1_t LPM_KEY_SEL1;
    we_LPM_KEY_SEL2_t LPM_KEY_SEL2;
    we_LPM_KEY_SEL3_t LPM_KEY_SEL3;
} mby_ppe_cgrp_a_nested_map_handcoded_t;

typedef logic [15:0] re_EM_HASH_LOOKUP_t;

typedef logic [7:0] re_LPM_SUBTRIE_APTR_t;

typedef logic [7:0] re_LPM_SUBTRIE_CPTR_t;

typedef logic [7:0] re_LPM_SUBTRIE_BITMAPS_t;

typedef logic [7:0] re_LPM_MATCH_TCAM_t;

typedef logic [7:0] re_LPM_MATCH_ACTION_t;

typedef logic [7:0] re_LPM_KEY_MASK_t;

typedef logic [7:0] re_LPM_KEY_SEL0_t;

typedef logic [7:0] re_LPM_KEY_SEL1_t;

typedef logic [7:0] re_LPM_KEY_SEL2_t;

typedef logic [7:0] re_LPM_KEY_SEL3_t;

typedef struct packed {
    re_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    re_LPM_SUBTRIE_APTR_t LPM_SUBTRIE_APTR;
    re_LPM_SUBTRIE_CPTR_t LPM_SUBTRIE_CPTR;
    re_LPM_SUBTRIE_BITMAPS_t LPM_SUBTRIE_BITMAPS;
    re_LPM_MATCH_TCAM_t LPM_MATCH_TCAM;
    re_LPM_MATCH_ACTION_t LPM_MATCH_ACTION;
    re_LPM_KEY_MASK_t LPM_KEY_MASK;
    re_LPM_KEY_SEL0_t LPM_KEY_SEL0;
    re_LPM_KEY_SEL1_t LPM_KEY_SEL1;
    re_LPM_KEY_SEL2_t LPM_KEY_SEL2;
    re_LPM_KEY_SEL3_t LPM_KEY_SEL3;
} mby_ppe_cgrp_a_nested_map_hc_re_t;

typedef logic handcode_rvalid_EM_HASH_LOOKUP_t;

typedef logic handcode_rvalid_LPM_SUBTRIE_APTR_t;

typedef logic handcode_rvalid_LPM_SUBTRIE_CPTR_t;

typedef logic handcode_rvalid_LPM_SUBTRIE_BITMAPS_t;

typedef logic handcode_rvalid_LPM_MATCH_TCAM_t;

typedef logic handcode_rvalid_LPM_MATCH_ACTION_t;

typedef logic handcode_rvalid_LPM_KEY_MASK_t;

typedef logic handcode_rvalid_LPM_KEY_SEL0_t;

typedef logic handcode_rvalid_LPM_KEY_SEL1_t;

typedef logic handcode_rvalid_LPM_KEY_SEL2_t;

typedef logic handcode_rvalid_LPM_KEY_SEL3_t;

typedef struct packed {
    handcode_rvalid_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    handcode_rvalid_LPM_SUBTRIE_APTR_t LPM_SUBTRIE_APTR;
    handcode_rvalid_LPM_SUBTRIE_CPTR_t LPM_SUBTRIE_CPTR;
    handcode_rvalid_LPM_SUBTRIE_BITMAPS_t LPM_SUBTRIE_BITMAPS;
    handcode_rvalid_LPM_MATCH_TCAM_t LPM_MATCH_TCAM;
    handcode_rvalid_LPM_MATCH_ACTION_t LPM_MATCH_ACTION;
    handcode_rvalid_LPM_KEY_MASK_t LPM_KEY_MASK;
    handcode_rvalid_LPM_KEY_SEL0_t LPM_KEY_SEL0;
    handcode_rvalid_LPM_KEY_SEL1_t LPM_KEY_SEL1;
    handcode_rvalid_LPM_KEY_SEL2_t LPM_KEY_SEL2;
    handcode_rvalid_LPM_KEY_SEL3_t LPM_KEY_SEL3;
} mby_ppe_cgrp_a_nested_map_hc_rvalid_t;

typedef logic handcode_wvalid_EM_HASH_LOOKUP_t;

typedef logic handcode_wvalid_LPM_SUBTRIE_APTR_t;

typedef logic handcode_wvalid_LPM_SUBTRIE_CPTR_t;

typedef logic handcode_wvalid_LPM_SUBTRIE_BITMAPS_t;

typedef logic handcode_wvalid_LPM_MATCH_TCAM_t;

typedef logic handcode_wvalid_LPM_MATCH_ACTION_t;

typedef logic handcode_wvalid_LPM_KEY_MASK_t;

typedef logic handcode_wvalid_LPM_KEY_SEL0_t;

typedef logic handcode_wvalid_LPM_KEY_SEL1_t;

typedef logic handcode_wvalid_LPM_KEY_SEL2_t;

typedef logic handcode_wvalid_LPM_KEY_SEL3_t;

typedef struct packed {
    handcode_wvalid_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    handcode_wvalid_LPM_SUBTRIE_APTR_t LPM_SUBTRIE_APTR;
    handcode_wvalid_LPM_SUBTRIE_CPTR_t LPM_SUBTRIE_CPTR;
    handcode_wvalid_LPM_SUBTRIE_BITMAPS_t LPM_SUBTRIE_BITMAPS;
    handcode_wvalid_LPM_MATCH_TCAM_t LPM_MATCH_TCAM;
    handcode_wvalid_LPM_MATCH_ACTION_t LPM_MATCH_ACTION;
    handcode_wvalid_LPM_KEY_MASK_t LPM_KEY_MASK;
    handcode_wvalid_LPM_KEY_SEL0_t LPM_KEY_SEL0;
    handcode_wvalid_LPM_KEY_SEL1_t LPM_KEY_SEL1;
    handcode_wvalid_LPM_KEY_SEL2_t LPM_KEY_SEL2;
    handcode_wvalid_LPM_KEY_SEL3_t LPM_KEY_SEL3;
} mby_ppe_cgrp_a_nested_map_hc_wvalid_t;

typedef logic handcode_error_EM_HASH_LOOKUP_t;

typedef logic handcode_error_LPM_SUBTRIE_APTR_t;

typedef logic handcode_error_LPM_SUBTRIE_CPTR_t;

typedef logic handcode_error_LPM_SUBTRIE_BITMAPS_t;

typedef logic handcode_error_LPM_MATCH_TCAM_t;

typedef logic handcode_error_LPM_MATCH_ACTION_t;

typedef logic handcode_error_LPM_KEY_MASK_t;

typedef logic handcode_error_LPM_KEY_SEL0_t;

typedef logic handcode_error_LPM_KEY_SEL1_t;

typedef logic handcode_error_LPM_KEY_SEL2_t;

typedef logic handcode_error_LPM_KEY_SEL3_t;

typedef struct packed {
    handcode_error_EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    handcode_error_LPM_SUBTRIE_APTR_t LPM_SUBTRIE_APTR;
    handcode_error_LPM_SUBTRIE_CPTR_t LPM_SUBTRIE_CPTR;
    handcode_error_LPM_SUBTRIE_BITMAPS_t LPM_SUBTRIE_BITMAPS;
    handcode_error_LPM_MATCH_TCAM_t LPM_MATCH_TCAM;
    handcode_error_LPM_MATCH_ACTION_t LPM_MATCH_ACTION;
    handcode_error_LPM_KEY_MASK_t LPM_KEY_MASK;
    handcode_error_LPM_KEY_SEL0_t LPM_KEY_SEL0;
    handcode_error_LPM_KEY_SEL1_t LPM_KEY_SEL1;
    handcode_error_LPM_KEY_SEL2_t LPM_KEY_SEL2;
    handcode_error_LPM_KEY_SEL3_t LPM_KEY_SEL3;
} mby_ppe_cgrp_a_nested_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    LPM_SUBTRIE_APTR_t LPM_SUBTRIE_APTR;
    LPM_SUBTRIE_CPTR_t LPM_SUBTRIE_CPTR;
    LPM_SUBTRIE_BITMAPS_t LPM_SUBTRIE_BITMAPS;
    LPM_MATCH_TCAM_t LPM_MATCH_TCAM;
    LPM_MATCH_ACTION_t LPM_MATCH_ACTION;
    LPM_KEY_MASK_t LPM_KEY_MASK;
    LPM_KEY_SEL0_t LPM_KEY_SEL0;
    LPM_KEY_SEL1_t LPM_KEY_SEL1;
    LPM_KEY_SEL2_t LPM_KEY_SEL2;
    LPM_KEY_SEL3_t LPM_KEY_SEL3;
} mby_ppe_cgrp_a_nested_map_hc_reg_read_t;

typedef struct packed {
    EM_HASH_LOOKUP_t EM_HASH_LOOKUP;
    LPM_SUBTRIE_APTR_t LPM_SUBTRIE_APTR;
    LPM_SUBTRIE_CPTR_t LPM_SUBTRIE_CPTR;
    LPM_SUBTRIE_BITMAPS_t LPM_SUBTRIE_BITMAPS;
    LPM_MATCH_TCAM_t LPM_MATCH_TCAM;
    LPM_MATCH_ACTION_t LPM_MATCH_ACTION;
    LPM_KEY_MASK_t LPM_KEY_MASK;
    LPM_KEY_SEL0_t LPM_KEY_SEL0;
    LPM_KEY_SEL1_t LPM_KEY_SEL1;
    LPM_KEY_SEL2_t LPM_KEY_SEL2;
    LPM_KEY_SEL3_t LPM_KEY_SEL3;
} mby_ppe_cgrp_a_nested_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_cgrp_a_nested_map_pkg

`endif // MBY_PPE_CGRP_A_NESTED_MAP_PKG_VH
