rtlgen_pkg_v12.vh