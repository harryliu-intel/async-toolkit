package tlm_env_pkg;

`include "tlm_defines.sv"

 
`ifdef XVM
   import ovm_pkg::*;
   import xvm_pkg::*;
   `include "ovm_macros.svh"
   `include "sla_macros.svh"
`endif

import sla_pkg::*;
 import uvm_pkg::*;
 import sla_fusegen_pkg::*;
  
`include "uvm_macros.svh"
`include "slu_macros.svh"
  
`include "tlm_types.sv"
`include "tlm_params.sv"
`include "tlm_rtl_config.sv"
`include "tlm_config.sv"
`include "tlm_env_monitor.sv"
`include "tlm_base_env.sv"
`include "tlm_env.sv"
`include "tlm_ral_env.sv"
`include "tlm_sm_env.sv"
`include "tlm_im_env.sv"
`include "tlm_seqlib.sv"
`include "tlm_fuse_env.sv" // this is not reusable
  
endpackage :tlm_env_pkg
