
// vim: noai : ts=3 : sw=3 : expandtab : ft=systemverilog

//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors.  The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//   Author        : Akshay Kotian
//   Project       : Madison Bay
//------------------------------------------------------------------------------

//   Package:    mby_gpol_test_lib
//
//   This is the main Test program file which holds all tests that will be ran in GPOL env.

`ifndef __MBY_GPOL_TEST_LIB_GUARD
`define __MBY_GPOL_TEST_LIB_GUARD

program mby_gpol_test_lib;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    import shdv_base_pkg::*;
    import mby_gpol_env_pkg::*;

    `include "mby_gpol_base_test.svh"
    `include "mby_gpol_doa_test.svh"

    // UVM Start test
    initial begin
        string testname;

        if ($value$plusargs("UVM_TESTNAME=%s", testname  )) begin
            $display ("MBY_tb Started Running %s in UVM mode!\n",testname);
        end
        uvm_pkg::run_test(testname);

end

endprogram

`endif // __MBY_GPOL_TEST_LIB_GUARD
