magic
tech scmos
timestamp 988943070
<< nselect >>
rect -34 47 0 84
rect -70 -12 0 42
<< pselect >>
rect 0 47 34 84
rect 0 -12 73 42
<< ndiffusion >>
rect -28 72 -8 73
rect -28 68 -8 69
rect -28 59 -8 60
rect -28 55 -8 56
rect -58 33 -50 34
rect -28 33 -8 34
rect -58 25 -50 30
rect -28 25 -8 30
rect -58 21 -50 22
rect -58 12 -50 13
rect -58 4 -50 9
rect -28 21 -8 22
rect -28 12 -8 13
rect -28 4 -8 9
rect -58 0 -50 1
rect -28 0 -8 1
<< pdiffusion >>
rect 8 72 28 73
rect 8 68 28 69
rect 8 59 28 60
rect 8 55 28 56
rect 8 33 28 34
rect 49 33 61 34
rect 8 25 28 30
rect 8 21 28 22
rect 8 12 28 13
rect 49 25 61 30
rect 49 21 61 22
rect 49 12 61 13
rect 8 4 28 9
rect 49 4 61 9
rect 8 0 28 1
rect 49 0 61 1
<< ntransistor >>
rect -28 69 -8 72
rect -28 56 -8 59
rect -58 30 -50 33
rect -28 30 -8 33
rect -58 22 -50 25
rect -28 22 -8 25
rect -58 9 -50 12
rect -28 9 -8 12
rect -58 1 -50 4
rect -28 1 -8 4
<< ptransistor >>
rect 8 69 28 72
rect 8 56 28 59
rect 8 30 28 33
rect 49 30 61 33
rect 8 22 28 25
rect 49 22 61 25
rect 8 9 28 12
rect 49 9 61 12
rect 8 1 28 4
rect 49 1 61 4
<< polysilicon >>
rect -33 69 -28 72
rect -8 69 -4 72
rect -33 59 -30 69
rect -33 56 -28 59
rect -8 56 -4 59
rect 4 69 8 72
rect 28 69 33 72
rect 30 59 33 69
rect 4 56 8 59
rect 28 56 33 59
rect -62 30 -58 33
rect -50 30 -28 33
rect -8 30 8 33
rect 28 30 49 33
rect 61 30 65 33
rect -63 22 -58 25
rect -50 22 -45 25
rect -40 22 -28 25
rect -8 22 8 25
rect 28 22 32 25
rect -63 17 -60 22
rect -62 12 -60 17
rect -62 9 -58 12
rect -50 9 -45 12
rect -40 4 -37 22
rect 37 12 40 30
rect 45 22 49 25
rect 61 22 66 25
rect 63 17 66 22
rect 63 12 65 17
rect -32 9 -28 12
rect -8 9 8 12
rect 28 9 40 12
rect 45 9 49 12
rect 61 9 65 12
rect -62 1 -58 4
rect -50 1 -28 4
rect -8 1 8 4
rect 28 1 49 4
rect 61 1 65 4
<< ndcontact >>
rect -28 73 -8 81
rect -28 60 -8 68
rect -28 47 -8 55
rect -58 34 -50 42
rect -28 34 -8 42
rect -58 13 -50 21
rect -28 13 -8 21
rect -58 -8 -50 0
rect -28 -8 -8 0
<< pdcontact >>
rect 8 73 28 81
rect 8 60 28 68
rect 8 47 28 55
rect 8 34 28 42
rect 49 34 61 42
rect 8 13 28 21
rect 49 13 61 21
rect 8 -8 28 0
rect 49 -8 61 0
<< polycontact >>
rect -4 56 4 72
rect -70 9 -62 17
rect 65 9 73 17
<< metal1 >>
rect -28 75 -27 81
rect -9 75 -8 81
rect -28 73 -8 75
rect 8 75 9 81
rect 27 75 28 81
rect 8 73 28 75
rect -28 60 -8 63
rect -4 56 4 72
rect 8 60 28 63
rect -28 42 -8 55
rect -58 40 -8 42
rect -58 34 -27 40
rect -9 34 -8 40
rect 8 42 28 55
rect 8 40 61 42
rect 8 34 9 40
rect 27 34 61 40
rect -70 9 -62 17
rect -58 13 61 21
rect 65 9 73 17
rect -67 4 70 9
rect -58 -2 -8 0
rect -58 -8 -27 -2
rect -9 -8 -8 -2
rect 8 -2 61 0
rect 8 -8 9 -2
rect 27 -8 61 -2
<< m2contact >>
rect -27 75 -9 81
rect 9 75 27 81
rect -28 63 -8 69
rect 8 63 28 69
rect -27 34 -9 40
rect 9 34 27 40
rect -27 -8 -9 -2
rect 9 -8 27 -2
<< metal2 >>
rect -28 63 28 69
<< m3contact >>
rect -27 75 -9 81
rect 9 75 27 81
rect -27 34 -9 40
rect 9 34 27 40
rect -27 -8 -9 -2
rect 9 -8 27 -2
<< metal3 >>
rect -27 -12 -9 84
rect 9 -12 27 84
<< labels >>
rlabel metal1 -66 13 -66 13 1 x
rlabel metal1 69 13 69 13 1 x
rlabel space -71 -12 -28 46 7 ^n1
rlabel space 28 -12 74 46 3 ^p1
rlabel space 28 47 35 84 3 ^p2
rlabel space -35 47 -28 84 7 ^n2
rlabel metal3 -27 -12 -9 84 1 GND!|pin|s|0
rlabel metal3 9 -12 27 84 1 Vdd!|pin|s|1
rlabel metal1 -58 34 -8 42 1 GND!|pin|s|0
rlabel metal1 -58 -8 -8 0 1 GND!|pin|s|0
rlabel metal1 -28 -8 -8 0 1 GND!|pin|s|0
rlabel metal1 -28 34 -8 42 1 GND!|pin|s|0
rlabel metal1 -28 47 -8 55 1 GND!|pin|s|0
rlabel metal1 -28 73 -8 81 1 GND!|pin|s|0
rlabel metal1 -28 42 -8 47 1 GND!|pin|s|0
rlabel metal1 8 42 28 47 1 Vdd!|pin|s|1
rlabel metal1 8 47 28 55 1 Vdd!|pin|s|1
rlabel metal1 8 73 28 81 1 Vdd!|pin|s|1
rlabel metal1 8 34 61 42 1 Vdd!|pin|s|1
rlabel metal1 8 34 28 42 1 Vdd!|pin|s|1
rlabel metal1 8 -8 61 0 1 Vdd!|pin|s|1
rlabel metal1 8 -8 28 0 1 Vdd!|pin|s|1
rlabel polysilicon -2 1 2 4 1 a|pin|w|3|poly
rlabel polysilicon -62 1 -58 4 1 a|pin|w|3|poly
rlabel polysilicon -2 30 2 33 1 b|pin|w|4|poly
rlabel polysilicon 61 30 65 33 1 b|pin|w|4|poly
rlabel metal2 -28 63 28 69 1 x|pin|s|7
rlabel metal1 -4 56 4 72 1 _x|pin|s|6
rlabel metal1 -58 13 61 21 1 _x|pin|s|5
rlabel metal1 -67 4 70 9 1 x|pin|s|8
<< end >>
