///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cm_apply_map.sv                                    
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_cm_apply_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_FF
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_FF

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_RSTD


module rtlgen_mby_ppe_cm_apply_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_cm_apply_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_PH2_FF
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CM_APPLY_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_cm_apply_map ( //lintra s-2096
    // Clocks
    gated_clk,

    // Resets
    rst_n,


    // Register Inputs
    new_CM_APPLY_STATE,

    handcode_reg_rdata_CM_APPLY_DROP_COUNT,
    handcode_reg_rdata_CM_APPLY_LOOPBACK_SUPPRESS,
    handcode_reg_rdata_CM_APPLY_MIRROR_PROFILE_TABLE,
    handcode_reg_rdata_CM_APPLY_QCN_CFG,
    handcode_reg_rdata_CM_APPLY_RX_SMP_STATE,
    handcode_reg_rdata_CM_APPLY_SOFTDROP_CFG,
    handcode_reg_rdata_CM_APPLY_SOFTDROP_STATE,
    handcode_reg_rdata_CM_APPLY_TX_SOFTDROP_CFG,
    handcode_reg_rdata_CM_APPLY_TX_TC_QCN_WM_THRESHOLD,
    handcode_reg_rdata_CM_APPLY_TX_TC_STATE,

    handcode_rvalid_CM_APPLY_DROP_COUNT,
    handcode_rvalid_CM_APPLY_LOOPBACK_SUPPRESS,
    handcode_rvalid_CM_APPLY_MIRROR_PROFILE_TABLE,
    handcode_rvalid_CM_APPLY_QCN_CFG,
    handcode_rvalid_CM_APPLY_RX_SMP_STATE,
    handcode_rvalid_CM_APPLY_SOFTDROP_CFG,
    handcode_rvalid_CM_APPLY_SOFTDROP_STATE,
    handcode_rvalid_CM_APPLY_TX_SOFTDROP_CFG,
    handcode_rvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD,
    handcode_rvalid_CM_APPLY_TX_TC_STATE,

    handcode_wvalid_CM_APPLY_DROP_COUNT,
    handcode_wvalid_CM_APPLY_LOOPBACK_SUPPRESS,
    handcode_wvalid_CM_APPLY_MIRROR_PROFILE_TABLE,
    handcode_wvalid_CM_APPLY_QCN_CFG,
    handcode_wvalid_CM_APPLY_RX_SMP_STATE,
    handcode_wvalid_CM_APPLY_SOFTDROP_CFG,
    handcode_wvalid_CM_APPLY_SOFTDROP_STATE,
    handcode_wvalid_CM_APPLY_TX_SOFTDROP_CFG,
    handcode_wvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD,
    handcode_wvalid_CM_APPLY_TX_TC_STATE,

    handcode_error_CM_APPLY_DROP_COUNT,
    handcode_error_CM_APPLY_LOOPBACK_SUPPRESS,
    handcode_error_CM_APPLY_MIRROR_PROFILE_TABLE,
    handcode_error_CM_APPLY_QCN_CFG,
    handcode_error_CM_APPLY_RX_SMP_STATE,
    handcode_error_CM_APPLY_SOFTDROP_CFG,
    handcode_error_CM_APPLY_SOFTDROP_STATE,
    handcode_error_CM_APPLY_TX_SOFTDROP_CFG,
    handcode_error_CM_APPLY_TX_TC_QCN_WM_THRESHOLD,
    handcode_error_CM_APPLY_TX_TC_STATE,


    // Register Outputs
    CM_APPLY_CPU_TRAP_MASK,
    CM_APPLY_LOG_MIRROR_PROFILE,
    CM_APPLY_MCAST_EPOCH,
    CM_APPLY_STATE,
    CM_APPLY_TC_TO_SMP,
    CM_APPLY_TRAP_GLORT,


    // Register signals for HandCoded registers
    handcode_reg_wdata_CM_APPLY_DROP_COUNT,
    handcode_reg_wdata_CM_APPLY_LOOPBACK_SUPPRESS,
    handcode_reg_wdata_CM_APPLY_MIRROR_PROFILE_TABLE,
    handcode_reg_wdata_CM_APPLY_QCN_CFG,
    handcode_reg_wdata_CM_APPLY_RX_SMP_STATE,
    handcode_reg_wdata_CM_APPLY_SOFTDROP_CFG,
    handcode_reg_wdata_CM_APPLY_SOFTDROP_STATE,
    handcode_reg_wdata_CM_APPLY_TX_SOFTDROP_CFG,
    handcode_reg_wdata_CM_APPLY_TX_TC_QCN_WM_THRESHOLD,
    handcode_reg_wdata_CM_APPLY_TX_TC_STATE,

    we_CM_APPLY_DROP_COUNT,
    we_CM_APPLY_LOOPBACK_SUPPRESS,
    we_CM_APPLY_MIRROR_PROFILE_TABLE,
    we_CM_APPLY_QCN_CFG,
    we_CM_APPLY_RX_SMP_STATE,
    we_CM_APPLY_SOFTDROP_CFG,
    we_CM_APPLY_SOFTDROP_STATE,
    we_CM_APPLY_TX_SOFTDROP_CFG,
    we_CM_APPLY_TX_TC_QCN_WM_THRESHOLD,
    we_CM_APPLY_TX_TC_STATE,

    re_CM_APPLY_DROP_COUNT,
    re_CM_APPLY_LOOPBACK_SUPPRESS,
    re_CM_APPLY_MIRROR_PROFILE_TABLE,
    re_CM_APPLY_QCN_CFG,
    re_CM_APPLY_RX_SMP_STATE,
    re_CM_APPLY_SOFTDROP_CFG,
    re_CM_APPLY_SOFTDROP_STATE,
    re_CM_APPLY_TX_SOFTDROP_CFG,
    re_CM_APPLY_TX_TC_QCN_WM_THRESHOLD,
    re_CM_APPLY_TX_TC_STATE,




    // Config Access
    req,
    ack
    

);

import mby_ppe_cm_apply_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:0] MBY_PPE_CM_APPLY_MAP_OFFSET = {MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] CM_APPLY_SB_BAR = 3'b0;
parameter [7:0] CM_APPLY_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
`define CM_APPLY_TRAP_GLORT_CR_ADDR_def(INDEX) CM_APPLY_TRAP_GLORT_CR_ADDR``INDEX``[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_APPLY_MAP_OFFSET[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
localparam [15:0][MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_APPLY_TRAP_GLORT_DECODE_ADDR = {`CM_APPLY_TRAP_GLORT_CR_ADDR_def([15]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([14]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([13]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([12]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([11]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([10]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([9]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([8]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([7]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([6]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([5]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([4]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([3]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([2]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([1]),`CM_APPLY_TRAP_GLORT_CR_ADDR_def([0])};
localparam [MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_APPLY_TC_TO_SMP_DECODE_ADDR = CM_APPLY_TC_TO_SMP_CR_ADDR[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_APPLY_MAP_OFFSET[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_APPLY_MCAST_EPOCH_DECODE_ADDR = CM_APPLY_MCAST_EPOCH_CR_ADDR[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_APPLY_MAP_OFFSET[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_APPLY_STATE_DECODE_ADDR = CM_APPLY_STATE_CR_ADDR[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_APPLY_MAP_OFFSET[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_APPLY_CPU_TRAP_MASK_DECODE_ADDR = CM_APPLY_CPU_TRAP_MASK_CR_ADDR[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_APPLY_MAP_OFFSET[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CM_APPLY_LOG_MIRROR_PROFILE_DECODE_ADDR = CM_APPLY_LOG_MIRROR_PROFILE_CR_ADDR[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CM_APPLY_MAP_OFFSET[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];

    // Clocks
input logic  gated_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input new_CM_APPLY_STATE_t  new_CM_APPLY_STATE;

input CM_APPLY_DROP_COUNT_t  handcode_reg_rdata_CM_APPLY_DROP_COUNT;
input CM_APPLY_LOOPBACK_SUPPRESS_t  handcode_reg_rdata_CM_APPLY_LOOPBACK_SUPPRESS;
input CM_APPLY_MIRROR_PROFILE_TABLE_t  handcode_reg_rdata_CM_APPLY_MIRROR_PROFILE_TABLE;
input CM_APPLY_QCN_CFG_t  handcode_reg_rdata_CM_APPLY_QCN_CFG;
input CM_APPLY_RX_SMP_STATE_t  handcode_reg_rdata_CM_APPLY_RX_SMP_STATE;
input CM_APPLY_SOFTDROP_CFG_t  handcode_reg_rdata_CM_APPLY_SOFTDROP_CFG;
input CM_APPLY_SOFTDROP_STATE_t  handcode_reg_rdata_CM_APPLY_SOFTDROP_STATE;
input CM_APPLY_TX_SOFTDROP_CFG_t  handcode_reg_rdata_CM_APPLY_TX_SOFTDROP_CFG;
input CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t  handcode_reg_rdata_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
input CM_APPLY_TX_TC_STATE_t  handcode_reg_rdata_CM_APPLY_TX_TC_STATE;

input handcode_rvalid_CM_APPLY_DROP_COUNT_t  handcode_rvalid_CM_APPLY_DROP_COUNT;
input handcode_rvalid_CM_APPLY_LOOPBACK_SUPPRESS_t  handcode_rvalid_CM_APPLY_LOOPBACK_SUPPRESS;
input handcode_rvalid_CM_APPLY_MIRROR_PROFILE_TABLE_t  handcode_rvalid_CM_APPLY_MIRROR_PROFILE_TABLE;
input handcode_rvalid_CM_APPLY_QCN_CFG_t  handcode_rvalid_CM_APPLY_QCN_CFG;
input handcode_rvalid_CM_APPLY_RX_SMP_STATE_t  handcode_rvalid_CM_APPLY_RX_SMP_STATE;
input handcode_rvalid_CM_APPLY_SOFTDROP_CFG_t  handcode_rvalid_CM_APPLY_SOFTDROP_CFG;
input handcode_rvalid_CM_APPLY_SOFTDROP_STATE_t  handcode_rvalid_CM_APPLY_SOFTDROP_STATE;
input handcode_rvalid_CM_APPLY_TX_SOFTDROP_CFG_t  handcode_rvalid_CM_APPLY_TX_SOFTDROP_CFG;
input handcode_rvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t  handcode_rvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
input handcode_rvalid_CM_APPLY_TX_TC_STATE_t  handcode_rvalid_CM_APPLY_TX_TC_STATE;

input handcode_wvalid_CM_APPLY_DROP_COUNT_t  handcode_wvalid_CM_APPLY_DROP_COUNT;
input handcode_wvalid_CM_APPLY_LOOPBACK_SUPPRESS_t  handcode_wvalid_CM_APPLY_LOOPBACK_SUPPRESS;
input handcode_wvalid_CM_APPLY_MIRROR_PROFILE_TABLE_t  handcode_wvalid_CM_APPLY_MIRROR_PROFILE_TABLE;
input handcode_wvalid_CM_APPLY_QCN_CFG_t  handcode_wvalid_CM_APPLY_QCN_CFG;
input handcode_wvalid_CM_APPLY_RX_SMP_STATE_t  handcode_wvalid_CM_APPLY_RX_SMP_STATE;
input handcode_wvalid_CM_APPLY_SOFTDROP_CFG_t  handcode_wvalid_CM_APPLY_SOFTDROP_CFG;
input handcode_wvalid_CM_APPLY_SOFTDROP_STATE_t  handcode_wvalid_CM_APPLY_SOFTDROP_STATE;
input handcode_wvalid_CM_APPLY_TX_SOFTDROP_CFG_t  handcode_wvalid_CM_APPLY_TX_SOFTDROP_CFG;
input handcode_wvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t  handcode_wvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
input handcode_wvalid_CM_APPLY_TX_TC_STATE_t  handcode_wvalid_CM_APPLY_TX_TC_STATE;

input handcode_error_CM_APPLY_DROP_COUNT_t  handcode_error_CM_APPLY_DROP_COUNT;
input handcode_error_CM_APPLY_LOOPBACK_SUPPRESS_t  handcode_error_CM_APPLY_LOOPBACK_SUPPRESS;
input handcode_error_CM_APPLY_MIRROR_PROFILE_TABLE_t  handcode_error_CM_APPLY_MIRROR_PROFILE_TABLE;
input handcode_error_CM_APPLY_QCN_CFG_t  handcode_error_CM_APPLY_QCN_CFG;
input handcode_error_CM_APPLY_RX_SMP_STATE_t  handcode_error_CM_APPLY_RX_SMP_STATE;
input handcode_error_CM_APPLY_SOFTDROP_CFG_t  handcode_error_CM_APPLY_SOFTDROP_CFG;
input handcode_error_CM_APPLY_SOFTDROP_STATE_t  handcode_error_CM_APPLY_SOFTDROP_STATE;
input handcode_error_CM_APPLY_TX_SOFTDROP_CFG_t  handcode_error_CM_APPLY_TX_SOFTDROP_CFG;
input handcode_error_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t  handcode_error_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
input handcode_error_CM_APPLY_TX_TC_STATE_t  handcode_error_CM_APPLY_TX_TC_STATE;


    // Register Outputs
output CM_APPLY_CPU_TRAP_MASK_t  CM_APPLY_CPU_TRAP_MASK;
output CM_APPLY_LOG_MIRROR_PROFILE_t  CM_APPLY_LOG_MIRROR_PROFILE;
output CM_APPLY_MCAST_EPOCH_t  CM_APPLY_MCAST_EPOCH;
output CM_APPLY_STATE_t  CM_APPLY_STATE;
output CM_APPLY_TC_TO_SMP_t  CM_APPLY_TC_TO_SMP;
output CM_APPLY_TRAP_GLORT_t [15:0] CM_APPLY_TRAP_GLORT;


    // Register signals for HandCoded registers
output CM_APPLY_DROP_COUNT_t  handcode_reg_wdata_CM_APPLY_DROP_COUNT;
output CM_APPLY_LOOPBACK_SUPPRESS_t  handcode_reg_wdata_CM_APPLY_LOOPBACK_SUPPRESS;
output CM_APPLY_MIRROR_PROFILE_TABLE_t  handcode_reg_wdata_CM_APPLY_MIRROR_PROFILE_TABLE;
output CM_APPLY_QCN_CFG_t  handcode_reg_wdata_CM_APPLY_QCN_CFG;
output CM_APPLY_RX_SMP_STATE_t  handcode_reg_wdata_CM_APPLY_RX_SMP_STATE;
output CM_APPLY_SOFTDROP_CFG_t  handcode_reg_wdata_CM_APPLY_SOFTDROP_CFG;
output CM_APPLY_SOFTDROP_STATE_t  handcode_reg_wdata_CM_APPLY_SOFTDROP_STATE;
output CM_APPLY_TX_SOFTDROP_CFG_t  handcode_reg_wdata_CM_APPLY_TX_SOFTDROP_CFG;
output CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t  handcode_reg_wdata_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
output CM_APPLY_TX_TC_STATE_t  handcode_reg_wdata_CM_APPLY_TX_TC_STATE;

output we_CM_APPLY_DROP_COUNT_t  we_CM_APPLY_DROP_COUNT;
output we_CM_APPLY_LOOPBACK_SUPPRESS_t  we_CM_APPLY_LOOPBACK_SUPPRESS;
output we_CM_APPLY_MIRROR_PROFILE_TABLE_t  we_CM_APPLY_MIRROR_PROFILE_TABLE;
output we_CM_APPLY_QCN_CFG_t  we_CM_APPLY_QCN_CFG;
output we_CM_APPLY_RX_SMP_STATE_t  we_CM_APPLY_RX_SMP_STATE;
output we_CM_APPLY_SOFTDROP_CFG_t  we_CM_APPLY_SOFTDROP_CFG;
output we_CM_APPLY_SOFTDROP_STATE_t  we_CM_APPLY_SOFTDROP_STATE;
output we_CM_APPLY_TX_SOFTDROP_CFG_t  we_CM_APPLY_TX_SOFTDROP_CFG;
output we_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t  we_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
output we_CM_APPLY_TX_TC_STATE_t  we_CM_APPLY_TX_TC_STATE;

output re_CM_APPLY_DROP_COUNT_t  re_CM_APPLY_DROP_COUNT;
output re_CM_APPLY_LOOPBACK_SUPPRESS_t  re_CM_APPLY_LOOPBACK_SUPPRESS;
output re_CM_APPLY_MIRROR_PROFILE_TABLE_t  re_CM_APPLY_MIRROR_PROFILE_TABLE;
output re_CM_APPLY_QCN_CFG_t  re_CM_APPLY_QCN_CFG;
output re_CM_APPLY_RX_SMP_STATE_t  re_CM_APPLY_RX_SMP_STATE;
output re_CM_APPLY_SOFTDROP_CFG_t  re_CM_APPLY_SOFTDROP_CFG;
output re_CM_APPLY_SOFTDROP_STATE_t  re_CM_APPLY_SOFTDROP_STATE;
output re_CM_APPLY_TX_SOFTDROP_CFG_t  re_CM_APPLY_TX_SOFTDROP_CFG;
output re_CM_APPLY_TX_TC_QCN_WM_THRESHOLD_t  re_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
output re_CM_APPLY_TX_TC_STATE_t  re_CM_APPLY_TX_TC_STATE;




    // Config Access
input mby_ppe_cm_apply_map_cr_req_t  req;
output mby_ppe_cm_apply_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_cm_apply_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_CM_APPLY_MAP_MEM;
assign case_req_addr_MBY_PPE_CM_APPLY_MAP_MEM = req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_cm_apply;
always_comb begin : sb_fid_cond_cm_apply_BLOCK
    unique casez (req_fid) 
		CM_APPLY_SB_FID: sb_fid_cond_cm_apply = 1;
		default: sb_fid_cond_cm_apply = 0;
    endcase 
end


logic sb_bar_cond_cm_apply;
always_comb begin : sb_bar_cond_cm_apply_BLOCK
    unique casez (req_bar) 
		CM_APPLY_SB_BAR: sb_bar_cond_cm_apply = 1;
		default: sb_bar_cond_cm_apply = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// CM_APPLY_TX_SOFTDROP_CFG using HANDCODED_REG template.
logic addr_decode_CM_APPLY_TX_SOFTDROP_CFG;
logic write_req_CM_APPLY_TX_SOFTDROP_CFG;
logic read_req_CM_APPLY_TX_SOFTDROP_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h0??,1'b?}: 
         addr_decode_CM_APPLY_TX_SOFTDROP_CFG = req.valid;
      default: 
         addr_decode_CM_APPLY_TX_SOFTDROP_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_TX_SOFTDROP_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_TX_SOFTDROP_CFG ;
always_comb read_req_CM_APPLY_TX_SOFTDROP_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_TX_SOFTDROP_CFG ;

always_comb we_CM_APPLY_TX_SOFTDROP_CFG = {8{write_req_CM_APPLY_TX_SOFTDROP_CFG}} & be;
always_comb re_CM_APPLY_TX_SOFTDROP_CFG = {8{read_req_CM_APPLY_TX_SOFTDROP_CFG}} & be;
always_comb handcode_reg_wdata_CM_APPLY_TX_SOFTDROP_CFG = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_TX_TC_STATE using HANDCODED_REG template.
logic addr_decode_CM_APPLY_TX_TC_STATE;
logic write_req_CM_APPLY_TX_TC_STATE;
logic read_req_CM_APPLY_TX_TC_STATE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h1??,1'b?}: 
         addr_decode_CM_APPLY_TX_TC_STATE = req.valid;
      default: 
         addr_decode_CM_APPLY_TX_TC_STATE = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_TX_TC_STATE = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_TX_TC_STATE ;
always_comb read_req_CM_APPLY_TX_TC_STATE  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_TX_TC_STATE ;

always_comb we_CM_APPLY_TX_TC_STATE = {8{write_req_CM_APPLY_TX_TC_STATE}} & be;
always_comb re_CM_APPLY_TX_TC_STATE = {8{read_req_CM_APPLY_TX_TC_STATE}} & be;
always_comb handcode_reg_wdata_CM_APPLY_TX_TC_STATE = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_TX_TC_QCN_WM_THRESHOLD using HANDCODED_REG template.
logic addr_decode_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
logic write_req_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
logic read_req_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h2??,1'b?}: 
         addr_decode_CM_APPLY_TX_TC_QCN_WM_THRESHOLD = req.valid;
      default: 
         addr_decode_CM_APPLY_TX_TC_QCN_WM_THRESHOLD = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_TX_TC_QCN_WM_THRESHOLD = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_TX_TC_QCN_WM_THRESHOLD ;
always_comb read_req_CM_APPLY_TX_TC_QCN_WM_THRESHOLD  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_TX_TC_QCN_WM_THRESHOLD ;

always_comb we_CM_APPLY_TX_TC_QCN_WM_THRESHOLD = {8{write_req_CM_APPLY_TX_TC_QCN_WM_THRESHOLD}} & be;
always_comb re_CM_APPLY_TX_TC_QCN_WM_THRESHOLD = {8{read_req_CM_APPLY_TX_TC_QCN_WM_THRESHOLD}} & be;
always_comb handcode_reg_wdata_CM_APPLY_TX_TC_QCN_WM_THRESHOLD = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_RX_SMP_STATE using HANDCODED_REG template.
logic addr_decode_CM_APPLY_RX_SMP_STATE;
logic write_req_CM_APPLY_RX_SMP_STATE;
logic read_req_CM_APPLY_RX_SMP_STATE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h3,4'b000?,4'h?,1'b?}: 
         addr_decode_CM_APPLY_RX_SMP_STATE = req.valid;
      default: 
         addr_decode_CM_APPLY_RX_SMP_STATE = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_RX_SMP_STATE = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_RX_SMP_STATE ;
always_comb read_req_CM_APPLY_RX_SMP_STATE  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_RX_SMP_STATE ;

always_comb we_CM_APPLY_RX_SMP_STATE = {8{write_req_CM_APPLY_RX_SMP_STATE}} & be;
always_comb re_CM_APPLY_RX_SMP_STATE = {8{read_req_CM_APPLY_RX_SMP_STATE}} & be;
always_comb handcode_reg_wdata_CM_APPLY_RX_SMP_STATE = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_MIRROR_PROFILE_TABLE using HANDCODED_REG template.
logic addr_decode_CM_APPLY_MIRROR_PROFILE_TABLE;
logic write_req_CM_APPLY_MIRROR_PROFILE_TABLE;
logic read_req_CM_APPLY_MIRROR_PROFILE_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h3,4'b001?,4'h?,1'b?}: 
         addr_decode_CM_APPLY_MIRROR_PROFILE_TABLE = req.valid;
      default: 
         addr_decode_CM_APPLY_MIRROR_PROFILE_TABLE = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_MIRROR_PROFILE_TABLE = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_MIRROR_PROFILE_TABLE ;
always_comb read_req_CM_APPLY_MIRROR_PROFILE_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_MIRROR_PROFILE_TABLE ;

always_comb we_CM_APPLY_MIRROR_PROFILE_TABLE = {8{write_req_CM_APPLY_MIRROR_PROFILE_TABLE}} & be;
always_comb re_CM_APPLY_MIRROR_PROFILE_TABLE = {8{read_req_CM_APPLY_MIRROR_PROFILE_TABLE}} & be;
always_comb handcode_reg_wdata_CM_APPLY_MIRROR_PROFILE_TABLE = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_DROP_COUNT using HANDCODED_REG template.
logic addr_decode_CM_APPLY_DROP_COUNT;
logic write_req_CM_APPLY_DROP_COUNT;
logic read_req_CM_APPLY_DROP_COUNT;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h34?,1'b?}: 
         addr_decode_CM_APPLY_DROP_COUNT = req.valid;
      default: 
         addr_decode_CM_APPLY_DROP_COUNT = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_DROP_COUNT = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_DROP_COUNT ;
always_comb read_req_CM_APPLY_DROP_COUNT  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_DROP_COUNT ;

always_comb we_CM_APPLY_DROP_COUNT = {8{write_req_CM_APPLY_DROP_COUNT}} & be;
always_comb re_CM_APPLY_DROP_COUNT = {8{read_req_CM_APPLY_DROP_COUNT}} & be;
always_comb handcode_reg_wdata_CM_APPLY_DROP_COUNT = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_LOOPBACK_SUPPRESS using HANDCODED_REG template.
logic addr_decode_CM_APPLY_LOOPBACK_SUPPRESS;
logic write_req_CM_APPLY_LOOPBACK_SUPPRESS;
logic read_req_CM_APPLY_LOOPBACK_SUPPRESS;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h35?,1'b?}: 
         addr_decode_CM_APPLY_LOOPBACK_SUPPRESS = req.valid;
      default: 
         addr_decode_CM_APPLY_LOOPBACK_SUPPRESS = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_LOOPBACK_SUPPRESS = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_LOOPBACK_SUPPRESS ;
always_comb read_req_CM_APPLY_LOOPBACK_SUPPRESS  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_LOOPBACK_SUPPRESS ;

always_comb we_CM_APPLY_LOOPBACK_SUPPRESS = {8{write_req_CM_APPLY_LOOPBACK_SUPPRESS}} & be;
always_comb re_CM_APPLY_LOOPBACK_SUPPRESS = {8{read_req_CM_APPLY_LOOPBACK_SUPPRESS}} & be;
always_comb handcode_reg_wdata_CM_APPLY_LOOPBACK_SUPPRESS = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_SOFTDROP_CFG using HANDCODED_REG template.
logic addr_decode_CM_APPLY_SOFTDROP_CFG;
logic write_req_CM_APPLY_SOFTDROP_CFG;
logic read_req_CM_APPLY_SOFTDROP_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h36,4'b00??,1'b?}: 
         addr_decode_CM_APPLY_SOFTDROP_CFG = req.valid;
      default: 
         addr_decode_CM_APPLY_SOFTDROP_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_SOFTDROP_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_SOFTDROP_CFG ;
always_comb read_req_CM_APPLY_SOFTDROP_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_SOFTDROP_CFG ;

always_comb we_CM_APPLY_SOFTDROP_CFG = {8{write_req_CM_APPLY_SOFTDROP_CFG}} & be;
always_comb re_CM_APPLY_SOFTDROP_CFG = {8{read_req_CM_APPLY_SOFTDROP_CFG}} & be;
always_comb handcode_reg_wdata_CM_APPLY_SOFTDROP_CFG = write_data;


// ----------------------------------------------------------------------
// CM_APPLY_SOFTDROP_STATE using HANDCODED_REG template.
logic addr_decode_CM_APPLY_SOFTDROP_STATE;
logic write_req_CM_APPLY_SOFTDROP_STATE;
logic read_req_CM_APPLY_SOFTDROP_STATE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h36,4'b01??,1'b?}: 
         addr_decode_CM_APPLY_SOFTDROP_STATE = req.valid;
      default: 
         addr_decode_CM_APPLY_SOFTDROP_STATE = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_SOFTDROP_STATE = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_SOFTDROP_STATE ;
always_comb read_req_CM_APPLY_SOFTDROP_STATE  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_SOFTDROP_STATE ;

always_comb we_CM_APPLY_SOFTDROP_STATE = {8{write_req_CM_APPLY_SOFTDROP_STATE}} & be;
always_comb re_CM_APPLY_SOFTDROP_STATE = {8{read_req_CM_APPLY_SOFTDROP_STATE}} & be;
always_comb handcode_reg_wdata_CM_APPLY_SOFTDROP_STATE = write_data;


//---------------------------------------------------------------------
// CM_APPLY_TRAP_GLORT Address Decode
logic [15:0] addr_decode_CM_APPLY_TRAP_GLORT;
logic [15:0] write_req_CM_APPLY_TRAP_GLORT;
always_comb begin
   addr_decode_CM_APPLY_TRAP_GLORT[0] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[0]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[1] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[1]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[2] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[2]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[3] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[3]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[4] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[4]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[5] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[5]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[6] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[6]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[7] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[7]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[8] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[8]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[9] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[9]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[10] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[10]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[11] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[11]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[12] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[12]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[13] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[13]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[14] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[14]) && req.valid ;
   addr_decode_CM_APPLY_TRAP_GLORT[15] = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TRAP_GLORT_DECODE_ADDR[15]) && req.valid ;
   write_req_CM_APPLY_TRAP_GLORT[0] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[0] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[1] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[1] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[2] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[2] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[3] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[3] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[4] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[4] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[5] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[5] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[6] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[6] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[7] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[7] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[8] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[8] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[9] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[9] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[10] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[10] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[11] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[11] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[12] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[12] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[13] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[13] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[14] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[14] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
   write_req_CM_APPLY_TRAP_GLORT[15] = IsMEMWr && addr_decode_CM_APPLY_TRAP_GLORT[15] && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
end

// ----------------------------------------------------------------------
// CM_APPLY_TRAP_GLORT.TRAP_GLORT x8 RW, using RW template.
logic [15:0][1:0] up_CM_APPLY_TRAP_GLORT_TRAP_GLORT;
always_comb begin
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[0] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[0] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[1] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[1] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[2] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[2] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[3] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[3] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[4] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[4] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[5] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[5] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[6] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[6] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[7] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[7] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[8] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[8] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[9] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[9] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[10] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[10] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[11] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[11] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[12] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[12] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[13] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[13] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[14] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[14] }} &
    be[1:0]);
 up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[15] =
    ({2{write_req_CM_APPLY_TRAP_GLORT[15] }} &
    be[1:0]);
end

logic [15:0][15:0] nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT;
always_comb begin
 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[0] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[1] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[2] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[3] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[4] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[5] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[6] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[7] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[8] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[9] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[10] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[11] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[12] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[13] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[14] = write_data[15:0];

 nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[15] = write_data[15:0];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[0][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[0][7:0], CM_APPLY_TRAP_GLORT[0].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[0][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[0][15:8], CM_APPLY_TRAP_GLORT[0].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[1][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[1][7:0], CM_APPLY_TRAP_GLORT[1].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[1][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[1][15:8], CM_APPLY_TRAP_GLORT[1].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[2][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[2][7:0], CM_APPLY_TRAP_GLORT[2].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[2][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[2][15:8], CM_APPLY_TRAP_GLORT[2].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[3][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[3][7:0], CM_APPLY_TRAP_GLORT[3].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[3][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[3][15:8], CM_APPLY_TRAP_GLORT[3].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[4][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[4][7:0], CM_APPLY_TRAP_GLORT[4].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[4][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[4][15:8], CM_APPLY_TRAP_GLORT[4].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[5][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[5][7:0], CM_APPLY_TRAP_GLORT[5].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[5][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[5][15:8], CM_APPLY_TRAP_GLORT[5].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[6][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[6][7:0], CM_APPLY_TRAP_GLORT[6].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[6][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[6][15:8], CM_APPLY_TRAP_GLORT[6].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[7][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[7][7:0], CM_APPLY_TRAP_GLORT[7].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[7][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[7][15:8], CM_APPLY_TRAP_GLORT[7].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[8][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[8][7:0], CM_APPLY_TRAP_GLORT[8].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[8][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[8][15:8], CM_APPLY_TRAP_GLORT[8].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[9][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[9][7:0], CM_APPLY_TRAP_GLORT[9].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[9][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[9][15:8], CM_APPLY_TRAP_GLORT[9].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[10][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[10][7:0], CM_APPLY_TRAP_GLORT[10].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[10][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[10][15:8], CM_APPLY_TRAP_GLORT[10].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[11][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[11][7:0], CM_APPLY_TRAP_GLORT[11].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[11][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[11][15:8], CM_APPLY_TRAP_GLORT[11].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[12][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[12][7:0], CM_APPLY_TRAP_GLORT[12].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[12][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[12][15:8], CM_APPLY_TRAP_GLORT[12].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[13][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[13][7:0], CM_APPLY_TRAP_GLORT[13].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[13][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[13][15:8], CM_APPLY_TRAP_GLORT[13].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[14][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[14][7:0], CM_APPLY_TRAP_GLORT[14].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[14][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[14][15:8], CM_APPLY_TRAP_GLORT[14].TRAP_GLORT[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[15][0], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[15][7:0], CM_APPLY_TRAP_GLORT[15].TRAP_GLORT[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_TRAP_GLORT_TRAP_GLORT[15][1], nxt_CM_APPLY_TRAP_GLORT_TRAP_GLORT[15][15:8], CM_APPLY_TRAP_GLORT[15].TRAP_GLORT[15:8])

//---------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP Address Decode
logic  addr_decode_CM_APPLY_TC_TO_SMP;
logic  write_req_CM_APPLY_TC_TO_SMP;
always_comb begin
   addr_decode_CM_APPLY_TC_TO_SMP = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_TC_TO_SMP_DECODE_ADDR) && req.valid ;
   write_req_CM_APPLY_TC_TO_SMP = IsMEMWr && addr_decode_CM_APPLY_TC_TO_SMP && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
end

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_0 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_0;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_0 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_0;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_0 = write_data[0:0];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_0[0], nxt_CM_APPLY_TC_TO_SMP_SMP_0[0:0], CM_APPLY_TC_TO_SMP.SMP_0[0:0])

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_1 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_1;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_1 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_1;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_1 = write_data[1:1];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_1[0], nxt_CM_APPLY_TC_TO_SMP_SMP_1[0:0], CM_APPLY_TC_TO_SMP.SMP_1[0:0])

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_2 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_2;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_2 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_2;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_2 = write_data[2:2];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_2[0], nxt_CM_APPLY_TC_TO_SMP_SMP_2[0:0], CM_APPLY_TC_TO_SMP.SMP_2[0:0])

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_3 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_3;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_3 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_3;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_3 = write_data[3:3];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_3[0], nxt_CM_APPLY_TC_TO_SMP_SMP_3[0:0], CM_APPLY_TC_TO_SMP.SMP_3[0:0])

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_4 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_4;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_4 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_4;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_4 = write_data[4:4];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_4[0], nxt_CM_APPLY_TC_TO_SMP_SMP_4[0:0], CM_APPLY_TC_TO_SMP.SMP_4[0:0])

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_5 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_5;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_5 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_5;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_5 = write_data[5:5];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_5[0], nxt_CM_APPLY_TC_TO_SMP_SMP_5[0:0], CM_APPLY_TC_TO_SMP.SMP_5[0:0])

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_6 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_6;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_6 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_6;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_6 = write_data[6:6];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_6[0], nxt_CM_APPLY_TC_TO_SMP_SMP_6[0:0], CM_APPLY_TC_TO_SMP.SMP_6[0:0])

// ----------------------------------------------------------------------
// CM_APPLY_TC_TO_SMP.SMP_7 x1 RW, using RW template.
logic [0:0] up_CM_APPLY_TC_TO_SMP_SMP_7;
always_comb begin
 up_CM_APPLY_TC_TO_SMP_SMP_7 =
    ({1{write_req_CM_APPLY_TC_TO_SMP }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_TC_TO_SMP_SMP_7;
always_comb begin
 nxt_CM_APPLY_TC_TO_SMP_SMP_7 = write_data[7:7];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_TC_TO_SMP_SMP_7[0], nxt_CM_APPLY_TC_TO_SMP_SMP_7[0:0], CM_APPLY_TC_TO_SMP.SMP_7[0:0])

//---------------------------------------------------------------------
// CM_APPLY_MCAST_EPOCH Address Decode
logic  addr_decode_CM_APPLY_MCAST_EPOCH;
logic  write_req_CM_APPLY_MCAST_EPOCH;
always_comb begin
   addr_decode_CM_APPLY_MCAST_EPOCH = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_MCAST_EPOCH_DECODE_ADDR) && req.valid ;
   write_req_CM_APPLY_MCAST_EPOCH = IsMEMWr && addr_decode_CM_APPLY_MCAST_EPOCH && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
end

// ----------------------------------------------------------------------
// CM_APPLY_MCAST_EPOCH.CURRENT x1 RW, using RW template.
logic [0:0] up_CM_APPLY_MCAST_EPOCH_CURRENT;
always_comb begin
 up_CM_APPLY_MCAST_EPOCH_CURRENT =
    ({1{write_req_CM_APPLY_MCAST_EPOCH }} &
    be[0:0]);
end

logic [0:0] nxt_CM_APPLY_MCAST_EPOCH_CURRENT;
always_comb begin
 nxt_CM_APPLY_MCAST_EPOCH_CURRENT = write_data[0:0];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_CM_APPLY_MCAST_EPOCH_CURRENT[0], nxt_CM_APPLY_MCAST_EPOCH_CURRENT[0:0], CM_APPLY_MCAST_EPOCH.CURRENT[0:0])

//---------------------------------------------------------------------
// CM_APPLY_STATE Address Decode
// ----------------------------------------------------------------------
// CM_APPLY_STATE.GLOBAL_EX x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.GLOBAL_EX = new_CM_APPLY_STATE.GLOBAL_EX;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_0 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_0 = new_CM_APPLY_STATE.RXS_0;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_1 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_1 = new_CM_APPLY_STATE.RXS_1;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_2 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_2 = new_CM_APPLY_STATE.RXS_2;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_3 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_3 = new_CM_APPLY_STATE.RXS_3;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_4 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_4 = new_CM_APPLY_STATE.RXS_4;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_5 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_5 = new_CM_APPLY_STATE.RXS_5;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_6 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_6 = new_CM_APPLY_STATE.RXS_6;



// ----------------------------------------------------------------------
// CM_APPLY_STATE.RXS_7 x1 RO/V, using RO/V template.
assign CM_APPLY_STATE.RXS_7 = new_CM_APPLY_STATE.RXS_7;




//---------------------------------------------------------------------
// CM_APPLY_CPU_TRAP_MASK Address Decode
logic  addr_decode_CM_APPLY_CPU_TRAP_MASK;
logic  write_req_CM_APPLY_CPU_TRAP_MASK;
always_comb begin
   addr_decode_CM_APPLY_CPU_TRAP_MASK = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_CPU_TRAP_MASK_DECODE_ADDR) && req.valid ;
   write_req_CM_APPLY_CPU_TRAP_MASK = IsMEMWr && addr_decode_CM_APPLY_CPU_TRAP_MASK && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
end

// ----------------------------------------------------------------------
// CM_APPLY_CPU_TRAP_MASK.DEST_MASK x8 RW, using RW template.
logic [2:0] up_CM_APPLY_CPU_TRAP_MASK_DEST_MASK;
always_comb begin
 up_CM_APPLY_CPU_TRAP_MASK_DEST_MASK =
    ({3{write_req_CM_APPLY_CPU_TRAP_MASK }} &
    be[2:0]);
end

logic [23:0] nxt_CM_APPLY_CPU_TRAP_MASK_DEST_MASK;
always_comb begin
 nxt_CM_APPLY_CPU_TRAP_MASK_DEST_MASK = write_data[23:0];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h1, up_CM_APPLY_CPU_TRAP_MASK_DEST_MASK[0], nxt_CM_APPLY_CPU_TRAP_MASK_DEST_MASK[7:0], CM_APPLY_CPU_TRAP_MASK.DEST_MASK[7:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_CPU_TRAP_MASK_DEST_MASK[1], nxt_CM_APPLY_CPU_TRAP_MASK_DEST_MASK[15:8], CM_APPLY_CPU_TRAP_MASK.DEST_MASK[15:8])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_CM_APPLY_CPU_TRAP_MASK_DEST_MASK[2], nxt_CM_APPLY_CPU_TRAP_MASK_DEST_MASK[23:16], CM_APPLY_CPU_TRAP_MASK.DEST_MASK[23:16])

//---------------------------------------------------------------------
// CM_APPLY_LOG_MIRROR_PROFILE Address Decode
logic  addr_decode_CM_APPLY_LOG_MIRROR_PROFILE;
logic  write_req_CM_APPLY_LOG_MIRROR_PROFILE;
always_comb begin
   addr_decode_CM_APPLY_LOG_MIRROR_PROFILE = (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CM_APPLY_LOG_MIRROR_PROFILE_DECODE_ADDR) && req.valid ;
   write_req_CM_APPLY_LOG_MIRROR_PROFILE = IsMEMWr && addr_decode_CM_APPLY_LOG_MIRROR_PROFILE && sb_fid_cond_cm_apply && sb_bar_cond_cm_apply;
end

// ----------------------------------------------------------------------
// CM_APPLY_LOG_MIRROR_PROFILE.FFU x6 RW, using RW template.
logic [0:0] up_CM_APPLY_LOG_MIRROR_PROFILE_FFU;
always_comb begin
 up_CM_APPLY_LOG_MIRROR_PROFILE_FFU =
    ({1{write_req_CM_APPLY_LOG_MIRROR_PROFILE }} &
    be[0:0]);
end

logic [5:0] nxt_CM_APPLY_LOG_MIRROR_PROFILE_FFU;
always_comb begin
 nxt_CM_APPLY_LOG_MIRROR_PROFILE_FFU = write_data[5:0];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 6'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_FFU[0], nxt_CM_APPLY_LOG_MIRROR_PROFILE_FFU[5:0], CM_APPLY_LOG_MIRROR_PROFILE.FFU[5:0])

// ----------------------------------------------------------------------
// CM_APPLY_LOG_MIRROR_PROFILE.RESERVED_MAC x4 RW, using RW template.
logic [1:0] up_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC;
always_comb begin
 up_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC =
    ({2{write_req_CM_APPLY_LOG_MIRROR_PROFILE }} &
    be[1:0]);
end

logic [5:0] nxt_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC;
always_comb begin
 nxt_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC = write_data[11:6];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC[0], nxt_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC[1:0], CM_APPLY_LOG_MIRROR_PROFILE.RESERVED_MAC[1:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 4'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC[1], nxt_CM_APPLY_LOG_MIRROR_PROFILE_RESERVED_MAC[5:2], CM_APPLY_LOG_MIRROR_PROFILE.RESERVED_MAC[5:2])

// ----------------------------------------------------------------------
// CM_APPLY_LOG_MIRROR_PROFILE.ARP_REDIRECT x2 RW, using RW template.
logic [1:0] up_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT;
always_comb begin
 up_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT =
    ({2{write_req_CM_APPLY_LOG_MIRROR_PROFILE }} &
    be[2:1]);
end

logic [5:0] nxt_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT;
always_comb begin
 nxt_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT = write_data[17:12];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 4'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT[0], nxt_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT[3:0], CM_APPLY_LOG_MIRROR_PROFILE.ARP_REDIRECT[3:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT[1], nxt_CM_APPLY_LOG_MIRROR_PROFILE_ARP_REDIRECT[5:4], CM_APPLY_LOG_MIRROR_PROFILE.ARP_REDIRECT[5:4])

// ----------------------------------------------------------------------
// CM_APPLY_LOG_MIRROR_PROFILE.ICMP x6 RW, using RW template.
logic [0:0] up_CM_APPLY_LOG_MIRROR_PROFILE_ICMP;
always_comb begin
 up_CM_APPLY_LOG_MIRROR_PROFILE_ICMP =
    ({1{write_req_CM_APPLY_LOG_MIRROR_PROFILE }} &
    be[2:2]);
end

logic [5:0] nxt_CM_APPLY_LOG_MIRROR_PROFILE_ICMP;
always_comb begin
 nxt_CM_APPLY_LOG_MIRROR_PROFILE_ICMP = write_data[23:18];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 6'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_ICMP[0], nxt_CM_APPLY_LOG_MIRROR_PROFILE_ICMP[5:0], CM_APPLY_LOG_MIRROR_PROFILE.ICMP[5:0])

// ----------------------------------------------------------------------
// CM_APPLY_LOG_MIRROR_PROFILE.TTL x6 RW, using RW template.
logic [0:0] up_CM_APPLY_LOG_MIRROR_PROFILE_TTL;
always_comb begin
 up_CM_APPLY_LOG_MIRROR_PROFILE_TTL =
    ({1{write_req_CM_APPLY_LOG_MIRROR_PROFILE }} &
    be[3:3]);
end

logic [5:0] nxt_CM_APPLY_LOG_MIRROR_PROFILE_TTL;
always_comb begin
 nxt_CM_APPLY_LOG_MIRROR_PROFILE_TTL = write_data[29:24];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 6'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_TTL[0], nxt_CM_APPLY_LOG_MIRROR_PROFILE_TTL[5:0], CM_APPLY_LOG_MIRROR_PROFILE.TTL[5:0])

// ----------------------------------------------------------------------
// CM_APPLY_LOG_MIRROR_PROFILE.TRIGGER x4 RW, using RW template.
logic [1:0] up_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER;
always_comb begin
 up_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER =
    ({2{write_req_CM_APPLY_LOG_MIRROR_PROFILE }} &
    be[4:3]);
end

logic [5:0] nxt_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER;
always_comb begin
 nxt_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER = write_data[35:30];

end


`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 2'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER[0], nxt_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER[1:0], CM_APPLY_LOG_MIRROR_PROFILE.TRIGGER[1:0])
`RTLGEN_MBY_PPE_CM_APPLY_MAP_EN_FF(gated_clk, rst_n, 4'h0, up_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER[1], nxt_CM_APPLY_LOG_MIRROR_PROFILE_TRIGGER[5:2], CM_APPLY_LOG_MIRROR_PROFILE.TRIGGER[5:2])

// ----------------------------------------------------------------------
// CM_APPLY_QCN_CFG using HANDCODED_REG template.
logic addr_decode_CM_APPLY_QCN_CFG;
logic write_req_CM_APPLY_QCN_CFG;
logic read_req_CM_APPLY_QCN_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CM_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h372,1'b1}: 
         addr_decode_CM_APPLY_QCN_CFG = req.valid;
      default: 
         addr_decode_CM_APPLY_QCN_CFG = 1'b0; 
   endcase
end

always_comb write_req_CM_APPLY_QCN_CFG = f_IsMEMWr(req_opcode) && addr_decode_CM_APPLY_QCN_CFG ;
always_comb read_req_CM_APPLY_QCN_CFG  = f_IsMEMRd(req_opcode) && addr_decode_CM_APPLY_QCN_CFG ;

always_comb we_CM_APPLY_QCN_CFG = {8{write_req_CM_APPLY_QCN_CFG}} & be;
always_comb re_CM_APPLY_QCN_CFG = {8{read_req_CM_APPLY_QCN_CFG}} & be;
always_comb handcode_reg_wdata_CM_APPLY_QCN_CFG = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_CM_APPLY_MAP_MEM) 
           {44'h0??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_TX_SOFTDROP_CFG;
                    ack.read_miss = handcode_error_CM_APPLY_TX_SOFTDROP_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h1??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_TX_TC_STATE;
                    ack.read_miss = handcode_error_CM_APPLY_TX_TC_STATE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h2??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
                    ack.read_miss = handcode_error_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h3,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_RX_SMP_STATE;
                    ack.read_miss = handcode_error_CM_APPLY_RX_SMP_STATE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h3,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_MIRROR_PROFILE_TABLE;
                    ack.read_miss = handcode_error_CM_APPLY_MIRROR_PROFILE_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h34?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_DROP_COUNT;
                    ack.read_miss = handcode_error_CM_APPLY_DROP_COUNT;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h35?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_LOOPBACK_SUPPRESS;
                    ack.read_miss = handcode_error_CM_APPLY_LOOPBACK_SUPPRESS;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h36,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_SOFTDROP_CFG;
                    ack.read_miss = handcode_error_CM_APPLY_SOFTDROP_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h36,4'b01??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_SOFTDROP_STATE;
                    ack.read_miss = handcode_error_CM_APPLY_SOFTDROP_STATE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_TC_TO_SMP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_MCAST_EPOCH_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_STATE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_CPU_TRAP_MASK_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           CM_APPLY_LOG_MIRROR_PROFILE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h372,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CM_APPLY_QCN_CFG;
                    ack.read_miss = handcode_error_CM_APPLY_QCN_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_CM_APPLY_MAP_MEM) 
           {44'h0??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_TX_SOFTDROP_CFG;
                    ack.write_miss = handcode_error_CM_APPLY_TX_SOFTDROP_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h1??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_TX_TC_STATE;
                    ack.write_miss = handcode_error_CM_APPLY_TX_TC_STATE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h2??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
                    ack.write_miss = handcode_error_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h3,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_RX_SMP_STATE;
                    ack.write_miss = handcode_error_CM_APPLY_RX_SMP_STATE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h3,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_MIRROR_PROFILE_TABLE;
                    ack.write_miss = handcode_error_CM_APPLY_MIRROR_PROFILE_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h34?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_DROP_COUNT;
                    ack.write_miss = handcode_error_CM_APPLY_DROP_COUNT;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h35?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_LOOPBACK_SUPPRESS;
                    ack.write_miss = handcode_error_CM_APPLY_LOOPBACK_SUPPRESS;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h36,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_SOFTDROP_CFG;
                    ack.write_miss = handcode_error_CM_APPLY_SOFTDROP_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h36,4'b01??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_SOFTDROP_STATE;
                    ack.write_miss = handcode_error_CM_APPLY_SOFTDROP_STATE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_TC_TO_SMP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_MCAST_EPOCH_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_STATE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_CPU_TRAP_MASK_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           CM_APPLY_LOG_MIRROR_PROFILE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h372,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CM_APPLY_QCN_CFG;
                    ack.write_miss = handcode_error_CM_APPLY_QCN_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_CM_APPLY_MAP_MEM) 
           {44'h0??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_TX_SOFTDROP_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'h1??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_TX_TC_STATE;
                 default: read_data = '0;
              endcase
           end
           {44'h2??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_TX_TC_QCN_WM_THRESHOLD;
                 default: read_data = '0;
              endcase
           end
           {36'h3,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_RX_SMP_STATE;
                 default: read_data = '0;
              endcase
           end
           {36'h3,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_MIRROR_PROFILE_TABLE;
                 default: read_data = '0;
              endcase
           end
           {44'h34?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_DROP_COUNT;
                 default: read_data = '0;
              endcase
           end
           {44'h35?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_LOOPBACK_SUPPRESS;
                 default: read_data = '0;
              endcase
           end
           {40'h36,4'b00??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_SOFTDROP_CFG;
                 default: read_data = '0;
              endcase
           end
           {40'h36,4'b01??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_SOFTDROP_STATE;
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[0]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[1]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[2]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[3]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[4]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[5]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[6]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[7]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[8]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[9]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[10]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[11]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[12]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[13]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[14]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TRAP_GLORT_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TRAP_GLORT[15]};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_TC_TO_SMP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_TC_TO_SMP};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_MCAST_EPOCH_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_MCAST_EPOCH};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_STATE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_STATE};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_CPU_TRAP_MASK_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_CPU_TRAP_MASK};
                 default: read_data = '0;
              endcase
           end
           CM_APPLY_LOG_MIRROR_PROFILE_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = {CM_APPLY_LOG_MIRROR_PROFILE};
                 default: read_data = '0;
              endcase
           end
           {44'h372,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {CM_APPLY_SB_FID,CM_APPLY_SB_BAR}: read_data = handcode_reg_rdata_CM_APPLY_QCN_CFG;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    CM_APPLY_TRAP_GLORT[0].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[1].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[2].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[3].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[4].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[5].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[6].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[7].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[8].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[9].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[10].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[11].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[12].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[13].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[14].reserved0 = '0;
    CM_APPLY_TRAP_GLORT[15].reserved0 = '0;
    CM_APPLY_TC_TO_SMP.reserved0 = '0;
    CM_APPLY_MCAST_EPOCH.reserved0 = '0;
    CM_APPLY_STATE.reserved0 = '0;
    CM_APPLY_CPU_TRAP_MASK.reserved0 = '0;
    CM_APPLY_LOG_MIRROR_PROFILE.reserved0 = '0;
end

// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
