magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -217 -713 -211 -712
rect -217 -719 -211 -715
rect -217 -725 -211 -721
rect -217 -731 -211 -727
rect -217 -734 -211 -733
rect -217 -738 -215 -734
rect -217 -739 -211 -738
rect -217 -745 -211 -741
rect -217 -751 -211 -747
rect -217 -757 -211 -753
rect -217 -760 -211 -759
<< pdiffusion >>
rect -199 -707 -189 -706
rect -199 -710 -189 -709
rect -191 -714 -189 -710
rect -199 -715 -189 -714
rect -199 -718 -189 -717
rect -199 -722 -193 -718
rect -199 -723 -189 -722
rect -199 -726 -189 -725
rect -191 -730 -189 -726
rect -199 -731 -189 -730
rect -199 -734 -189 -733
rect -199 -738 -193 -734
rect -199 -739 -189 -738
rect -199 -742 -189 -741
rect -191 -746 -189 -742
rect -199 -747 -189 -746
rect -199 -750 -189 -749
rect -199 -754 -193 -750
rect -199 -755 -189 -754
rect -199 -758 -189 -757
rect -191 -762 -189 -758
rect -199 -763 -189 -762
rect -199 -766 -189 -765
<< ntransistor >>
rect -217 -715 -211 -713
rect -217 -721 -211 -719
rect -217 -727 -211 -725
rect -217 -733 -211 -731
rect -217 -741 -211 -739
rect -217 -747 -211 -745
rect -217 -753 -211 -751
rect -217 -759 -211 -757
<< ptransistor >>
rect -199 -709 -189 -707
rect -199 -717 -189 -715
rect -199 -725 -189 -723
rect -199 -733 -189 -731
rect -199 -741 -189 -739
rect -199 -749 -189 -747
rect -199 -757 -189 -755
rect -199 -765 -189 -763
<< polysilicon >>
rect -203 -709 -199 -707
rect -189 -709 -186 -707
rect -203 -713 -201 -709
rect -220 -715 -217 -713
rect -211 -715 -201 -713
rect -203 -717 -199 -715
rect -189 -717 -186 -715
rect -220 -721 -217 -719
rect -211 -721 -208 -719
rect -203 -725 -199 -723
rect -189 -725 -186 -723
rect -220 -727 -217 -725
rect -211 -727 -201 -725
rect -203 -731 -201 -727
rect -220 -733 -217 -731
rect -211 -733 -208 -731
rect -203 -733 -199 -731
rect -189 -733 -186 -731
rect -220 -741 -217 -739
rect -211 -741 -208 -739
rect -203 -741 -199 -739
rect -189 -741 -186 -739
rect -203 -745 -201 -741
rect -220 -747 -217 -745
rect -211 -747 -201 -745
rect -203 -749 -199 -747
rect -189 -749 -186 -747
rect -220 -753 -217 -751
rect -211 -753 -208 -751
rect -203 -757 -199 -755
rect -189 -757 -186 -755
rect -220 -759 -217 -757
rect -211 -759 -201 -757
rect -203 -763 -201 -759
rect -203 -765 -199 -763
rect -189 -765 -186 -763
<< ndcontact >>
rect -217 -712 -211 -708
rect -215 -738 -211 -734
rect -217 -764 -211 -760
<< pdcontact >>
rect -199 -706 -189 -702
rect -199 -714 -191 -710
rect -193 -722 -189 -718
rect -199 -730 -191 -726
rect -193 -738 -189 -734
rect -199 -746 -191 -742
rect -193 -754 -189 -750
rect -199 -762 -191 -758
rect -199 -770 -189 -766
<< metal1 >>
rect -199 -706 -189 -702
rect -217 -712 -211 -708
rect -199 -714 -191 -710
rect -199 -726 -196 -714
rect -193 -722 -189 -718
rect -199 -730 -191 -726
rect -199 -734 -196 -730
rect -215 -738 -196 -734
rect -193 -738 -189 -734
rect -199 -742 -196 -738
rect -199 -746 -191 -742
rect -199 -758 -196 -746
rect -193 -754 -189 -750
rect -217 -764 -211 -760
rect -199 -762 -191 -758
rect -199 -770 -189 -766
<< labels >>
rlabel space -220 -765 -214 -707 7 ^n
rlabel polysilicon -218 -758 -218 -758 3 a
rlabel polysilicon -218 -714 -218 -714 3 d
rlabel polysilicon -218 -752 -218 -752 3 b
rlabel polysilicon -218 -746 -218 -746 3 c
rlabel polysilicon -218 -732 -218 -732 3 a
rlabel polysilicon -218 -740 -218 -740 3 d
rlabel polysilicon -218 -726 -218 -726 3 b
rlabel polysilicon -218 -720 -218 -720 3 c
rlabel polysilicon -188 -716 -188 -716 7 d
rlabel polysilicon -188 -708 -188 -708 7 d
rlabel polysilicon -188 -732 -188 -732 7 b
rlabel polysilicon -188 -724 -188 -724 7 b
rlabel polysilicon -188 -740 -188 -740 7 c
rlabel polysilicon -188 -748 -188 -748 7 c
rlabel polysilicon -188 -764 -188 -764 7 a
rlabel polysilicon -188 -756 -188 -756 7 a
rlabel space -192 -771 -185 -701 3 ^p
rlabel ndcontact -213 -710 -213 -710 5 GND!
rlabel ndcontact -213 -736 -213 -736 1 x
rlabel ndcontact -213 -762 -213 -762 1 GND!
rlabel pdcontact -197 -760 -197 -760 1 x
rlabel pdcontact -197 -744 -197 -744 1 x
rlabel pdcontact -197 -728 -197 -728 1 x
rlabel pdcontact -197 -712 -197 -712 1 x
rlabel pdcontact -191 -720 -191 -720 1 Vdd!
rlabel pdcontact -191 -736 -191 -736 1 Vdd!
rlabel pdcontact -191 -752 -191 -752 1 Vdd!
rlabel pdcontact -191 -768 -191 -768 1 Vdd!
rlabel pdcontact -191 -704 -191 -704 1 Vdd!
<< end >>
