magic
tech scmos
timestamp 970030226
<< ndiffusion >>
rect -21 151 -16 159
rect -21 150 -8 151
rect -24 141 -8 142
rect -24 133 -8 138
rect -67 117 -51 118
rect -24 125 -8 130
rect -24 117 -8 122
rect -67 109 -51 114
rect -24 109 -8 114
rect -67 105 -51 106
rect -67 97 -63 105
rect -55 97 -51 105
rect -24 105 -8 106
rect -67 96 -51 97
rect -24 97 -23 105
rect -24 96 -8 97
rect -67 88 -51 93
rect -24 88 -8 93
rect -67 84 -51 85
rect -24 80 -8 85
rect -24 72 -8 77
rect -67 64 -51 65
rect -24 64 -8 69
rect -67 56 -51 61
rect -24 60 -8 61
rect -67 52 -51 53
rect -67 44 -65 52
rect -67 43 -51 44
rect -67 39 -51 40
<< pdiffusion >>
rect 22 163 38 164
rect 22 157 38 160
rect 44 149 48 154
rect 22 148 48 149
rect 53 149 57 154
rect 53 148 65 149
rect 22 144 48 145
rect 44 136 48 144
rect 22 135 48 136
rect 53 144 65 145
rect 61 136 65 144
rect 53 135 65 136
rect 22 131 48 132
rect 22 123 30 131
rect 22 122 48 123
rect 53 131 65 132
rect 53 123 57 131
rect 53 122 65 123
rect 22 118 48 119
rect 44 110 48 118
rect 22 109 48 110
rect 53 118 65 119
rect 61 110 65 118
rect 53 109 65 110
rect 22 105 48 106
rect 41 97 48 105
rect 22 96 48 97
rect 53 105 65 106
rect 53 97 57 105
rect 53 96 65 97
rect 22 92 48 93
rect 41 84 48 92
rect 22 83 48 84
rect 53 92 65 93
rect 61 84 65 92
rect 53 83 65 84
rect 22 79 48 80
rect 22 71 30 79
rect 22 70 48 71
rect 53 79 65 80
rect 53 71 57 79
rect 53 70 65 71
rect 22 66 48 67
rect 44 58 48 66
rect 22 57 48 58
rect 53 66 65 67
rect 61 58 65 66
rect 53 57 65 58
rect 22 53 48 54
rect 22 51 32 53
rect 15 46 32 51
rect 15 43 27 46
rect 53 53 65 54
rect 53 45 57 53
rect 53 43 65 45
rect 15 39 27 40
rect 53 39 65 40
<< ntransistor >>
rect -24 138 -8 141
rect -24 130 -8 133
rect -24 122 -8 125
rect -67 114 -51 117
rect -24 114 -8 117
rect -67 106 -51 109
rect -24 106 -8 109
rect -67 93 -51 96
rect -24 93 -8 96
rect -67 85 -51 88
rect -24 85 -8 88
rect -24 77 -8 80
rect -24 69 -8 72
rect -67 61 -51 64
rect -24 61 -8 64
rect -67 53 -51 56
rect -67 40 -51 43
<< ptransistor >>
rect 22 160 38 163
rect 22 145 48 148
rect 53 145 65 148
rect 22 132 48 135
rect 53 132 65 135
rect 22 119 48 122
rect 53 119 65 122
rect 22 106 48 109
rect 53 106 65 109
rect 22 93 48 96
rect 53 93 65 96
rect 22 80 48 83
rect 53 80 65 83
rect 22 67 48 70
rect 53 67 65 70
rect 22 54 48 57
rect 53 54 65 57
rect 15 40 27 43
rect 53 40 65 43
<< polysilicon >>
rect 40 173 42 176
rect 40 163 43 173
rect 18 160 22 163
rect 38 160 43 163
rect -79 138 -38 141
rect 1 145 22 148
rect 48 145 53 148
rect 65 145 73 148
rect -30 138 -24 141
rect -8 138 -4 141
rect -79 64 -76 138
rect 1 133 4 145
rect -49 130 -24 133
rect -8 130 4 133
rect 9 132 22 135
rect 48 132 53 135
rect 65 132 69 135
rect -49 117 -46 130
rect 9 125 12 132
rect -33 122 -24 125
rect -8 122 12 125
rect 17 119 22 122
rect 48 119 53 122
rect 65 119 81 122
rect 17 117 20 119
rect -71 114 -67 117
rect -51 114 -46 117
rect -28 114 -24 117
rect -8 114 20 117
rect -71 106 -67 109
rect -51 106 -35 109
rect -27 106 -24 109
rect -8 106 22 109
rect 48 106 53 109
rect 65 106 69 109
rect -71 93 -67 96
rect -51 93 -48 96
rect -40 93 -24 96
rect -8 93 22 96
rect 48 93 53 96
rect 65 93 69 96
rect -71 85 -67 88
rect -51 85 -46 88
rect -28 85 -24 88
rect -8 85 20 88
rect -49 72 -46 85
rect 17 83 20 85
rect 17 80 22 83
rect 48 80 53 83
rect 65 80 73 83
rect -33 77 -24 80
rect -8 77 12 80
rect -49 69 -24 72
rect -8 69 4 72
rect -79 61 -67 64
rect -51 61 -24 64
rect -8 61 -4 64
rect -69 53 -67 56
rect -51 53 -45 56
rect 1 57 4 69
rect 9 70 12 77
rect 9 67 22 70
rect 48 67 53 70
rect 65 67 69 70
rect 1 54 22 57
rect 48 54 53 57
rect 65 54 81 57
rect -71 40 -67 43
rect -51 40 -4 43
rect 4 40 15 43
rect 27 40 31 43
rect 41 40 53 43
rect 65 40 69 43
rect 41 39 44 40
<< ndcontact >>
rect -24 142 -8 150
rect -67 118 -51 126
rect -63 97 -55 105
rect -23 97 -8 105
rect -67 65 -51 84
rect -65 44 -51 52
rect -24 52 -8 60
rect -67 31 -51 39
<< pdcontact >>
rect 22 164 38 172
rect 22 149 44 157
rect 57 149 65 157
rect 22 136 44 144
rect 53 136 61 144
rect 30 123 48 131
rect 57 123 65 131
rect 22 110 44 118
rect 53 110 61 118
rect 22 97 41 105
rect 57 97 65 105
rect 22 84 41 92
rect 53 84 61 92
rect 30 71 48 79
rect 57 71 65 79
rect 22 58 44 66
rect 53 58 61 66
rect 32 45 48 53
rect 57 45 65 53
rect 15 31 27 39
rect 53 31 65 39
<< psubstratepcontact >>
rect -16 151 -8 159
rect -41 45 -33 53
<< nsubstratencontact >>
rect 74 39 82 47
<< polycontact >>
rect 42 173 50 181
rect -38 138 -30 146
rect 73 140 81 148
rect -41 117 -33 125
rect 81 114 89 122
rect -35 101 -27 109
rect -48 93 -40 101
rect -41 77 -33 85
rect 73 80 81 88
rect -77 48 -69 56
rect 81 54 89 62
rect -4 40 4 48
rect 36 31 44 39
<< metal1 >>
rect -38 138 -30 175
rect -21 150 -8 175
rect -24 142 -8 150
rect 12 157 17 175
rect 42 173 50 175
rect 22 168 38 172
rect 22 164 53 168
rect 12 149 44 157
rect -71 118 -51 126
rect -41 121 -33 125
rect -71 84 -67 118
rect -44 115 -41 121
rect -63 97 -55 105
rect -44 101 -40 115
rect -48 93 -40 101
rect 12 105 18 149
rect 48 144 53 164
rect 57 153 65 157
rect 57 149 69 153
rect 22 136 44 144
rect 48 136 61 144
rect 22 118 26 136
rect 48 131 53 136
rect 65 131 69 149
rect 30 123 53 131
rect 57 123 69 131
rect 48 118 53 123
rect 22 110 44 118
rect 48 110 61 118
rect -35 101 -27 103
rect -35 85 -31 101
rect -23 97 -8 105
rect 12 97 41 105
rect 48 97 53 110
rect 65 105 69 123
rect 57 97 69 105
rect -71 80 -51 84
rect -67 65 -51 80
rect -41 81 -31 85
rect -41 77 -33 81
rect -77 48 -69 56
rect -41 52 -33 53
rect -24 52 -8 60
rect -73 39 -69 48
rect -65 49 -8 52
rect -65 44 -21 49
rect -3 48 3 91
rect 22 84 41 92
rect 53 91 61 92
rect 48 84 61 91
rect 22 66 26 84
rect 48 79 53 84
rect 65 79 69 97
rect 73 140 81 148
rect 73 88 77 140
rect 81 114 89 122
rect 73 85 81 88
rect 30 71 53 79
rect 57 71 69 79
rect 85 73 89 114
rect 48 66 53 71
rect 22 58 44 66
rect 48 62 61 66
rect 53 58 61 62
rect 65 53 69 71
rect 81 54 89 67
rect 32 49 53 53
rect -4 40 4 48
rect 57 49 69 53
rect 57 45 65 49
rect 48 39 53 43
rect 74 39 82 47
rect -73 35 -51 39
rect 15 35 44 39
rect -67 34 44 35
rect -67 31 27 34
rect 36 31 44 34
rect 48 35 78 39
rect 48 31 65 35
<< m2contact >>
rect -38 175 -30 181
rect -21 175 -3 181
rect 3 175 17 181
rect 42 175 50 181
rect -41 115 -33 121
rect -63 91 -55 97
rect -35 103 -27 109
rect -23 91 3 97
rect -21 43 -8 49
rect 45 91 53 97
rect 73 79 81 85
rect 81 67 89 73
rect 32 43 53 49
<< metal2 >>
rect -38 175 -27 181
rect 27 175 50 181
rect -41 115 0 121
rect -35 103 0 109
rect -63 91 53 97
rect 0 79 81 85
rect 0 67 89 73
rect 21 43 53 49
<< m3contact >>
rect -21 175 -3 181
rect 3 175 21 181
rect -21 43 -3 49
rect 3 43 21 49
<< metal3 >>
rect -21 28 -3 184
rect 3 28 21 184
<< labels >>
rlabel metal1 26 153 26 153 5 Vdd!
rlabel metal1 26 101 26 101 1 Vdd!
rlabel metal1 -12 146 -12 146 5 GND!
rlabel metal1 -12 56 -12 56 1 GND!
rlabel metal1 44 127 44 127 1 x
rlabel pdcontact 44 75 44 75 5 x
rlabel metal1 61 35 61 35 1 Vdd!
rlabel polysilicon 66 55 66 55 1 _a0
rlabel polysilicon 66 68 66 68 1 _b0
rlabel polysilicon 66 81 66 81 1 _b1
rlabel polysilicon 66 94 66 94 1 _a1
rlabel polysilicon 66 107 66 107 1 _b0
rlabel polysilicon 66 120 66 120 1 _a0
rlabel polysilicon 66 133 66 133 1 _a1
rlabel polysilicon 66 146 66 146 1 _b1
rlabel metal1 39 49 39 49 1 Vdd!
rlabel metal1 27 168 27 168 5 x
rlabel polysilicon 39 161 39 161 1 _PReset!
rlabel polysilicon -25 139 -25 139 1 _SReset!
rlabel polysilicon -68 62 -68 62 1 _SReset!
rlabel metal1 -59 101 -59 101 1 x
rlabel metal1 -15 101 -15 101 1 x
rlabel metal1 78 43 78 43 7 Vdd!
rlabel metal1 -37 50 -37 50 1 GND!
rlabel metal2 0 94 0 94 1 x
rlabel metal2 0 67 0 73 3 _a0
rlabel metal2 0 79 0 85 3 _b1
rlabel metal2 0 103 0 109 7 _b0
rlabel metal2 0 115 0 121 7 _a1
rlabel metal2 46 178 46 178 1 _PReset!
rlabel metal1 -58 48 -58 48 1 GND!
rlabel metal2 -34 178 -34 178 1 _SReset!
rlabel space -80 30 -24 182 7 ^n
rlabel metal2 -27 175 -27 181 3 ^n
rlabel space 35 30 83 50 3 ^p
rlabel space 35 51 91 151 3 ^p
rlabel space 44 152 70 169 3 ^p
rlabel metal2 -37 118 -37 118 1 _a1
rlabel metal2 -31 106 -31 106 1 _b0
rlabel metal2 -59 94 -59 94 1 x
rlabel metal2 49 94 49 94 1 x
rlabel metal2 77 82 77 82 1 _b1
rlabel metal2 85 70 85 70 1 _a0
<< end >>
