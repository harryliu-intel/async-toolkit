// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

module clkgen(output logic clk);

parameter FREQ_MHZ = 100.0;

initial begin
    clk = 0;
    forever #(1.0us/FREQ_MHZ/2.0) clk = !clk;
end

endmodule
