magic
tech scmos
timestamp 982690832
<< nselect >>
rect -47 22 -1 71
<< pselect >>
rect -1 22 77 76
<< ndiffusion >>
rect -43 50 -35 51
rect -21 52 -13 53
rect -43 46 -35 47
rect -21 44 -13 49
rect -21 36 -13 41
rect -21 32 -13 33
<< pdiffusion >>
rect 63 65 67 70
rect 55 64 67 65
rect 55 58 67 61
rect 55 49 71 50
rect 8 41 12 44
rect 8 32 12 37
rect 25 36 33 37
rect 55 45 71 46
rect 69 37 71 45
rect 55 36 71 37
rect 25 32 33 33
rect 55 32 71 33
<< ntransistor >>
rect -43 47 -35 50
rect -21 49 -13 52
rect -21 41 -13 44
rect -21 33 -13 36
<< ptransistor >>
rect 55 61 67 64
rect 55 46 71 49
rect 8 37 12 41
rect 25 33 33 36
rect 55 33 71 36
<< polysilicon >>
rect -33 50 -30 66
rect 51 61 55 64
rect 67 61 71 64
rect -47 47 -43 50
rect -35 47 -30 50
rect -25 49 -21 52
rect -13 49 -9 52
rect 50 46 55 49
rect 71 46 76 49
rect -25 41 -21 44
rect -13 41 -4 44
rect 4 37 8 41
rect 12 37 16 41
rect -25 33 -21 36
rect -13 33 -9 36
rect 37 36 40 37
rect 21 33 25 36
rect 33 33 40 36
rect 50 36 53 46
rect 73 36 76 46
rect 50 33 55 36
rect 71 33 76 36
<< ndcontact >>
rect -43 51 -35 59
rect -21 53 -13 61
rect -43 38 -35 46
rect -21 24 -13 32
<< pdcontact >>
rect 55 65 63 73
rect 8 44 16 52
rect 55 50 71 58
rect 25 37 33 45
rect 55 37 69 45
rect 8 24 16 32
rect 25 24 33 32
rect 55 24 71 32
<< polycontact >>
rect -41 63 -33 71
rect -4 36 4 44
rect 37 37 45 45
<< metal1 >>
rect -41 65 63 73
rect -41 63 -33 65
rect -43 55 -35 59
rect -43 51 -27 55
rect -21 53 -13 65
rect 8 55 16 65
rect 55 56 71 58
rect -43 32 -35 46
rect -31 44 -27 51
rect 8 49 42 55
rect 63 50 71 56
rect 8 44 16 49
rect 37 45 42 49
rect -31 40 4 44
rect 25 40 33 45
rect -4 37 33 40
rect 37 37 69 45
rect -4 36 29 37
rect -43 30 -13 32
rect 8 30 71 32
rect -43 24 -27 30
rect 8 24 9 30
rect 27 24 71 30
<< m2contact >>
rect 55 50 63 56
rect -27 24 -9 30
rect 9 24 27 30
<< metal2 >>
rect 27 50 63 56
<< m3contact >>
rect 9 50 27 56
rect -27 24 -9 30
rect 9 24 27 30
<< metal3 >>
rect -27 22 -9 76
rect 9 22 27 76
<< labels >>
rlabel space 71 22 78 58 3 ^p
rlabel metal3 -27 22 -9 76 1 GND!|pin|s|0
rlabel metal3 9 22 27 76 1 Vdd!|pin|s|1
rlabel metal1 -43 24 -13 32 1 GND!|pin|s|0
rlabel metal1 -43 24 -35 46 1 GND!|pin|s|0
rlabel metal1 8 24 71 32 1 Vdd!|pin|s|1
rlabel metal1 55 50 71 58 1 Vdd!|pin|s|1
rlabel metal1 -41 65 63 73 1 x|pin|s|2
rlabel metal1 8 44 16 73 1 x|pin|s|2
rlabel metal1 37 37 69 45 1 x|pin|s|2
rlabel polysilicon 50 33 53 49 1 a|pin|w|3|poly
rlabel polysilicon 73 33 76 49 1 a|pin|w|3|poly
rlabel polysilicon -13 49 -9 52 1 a|pin|w|4|poly
rlabel polysilicon -25 49 -21 52 1 a|pin|w|4|poly
rlabel polysilicon -25 33 -21 36 1 _SReset!|pin|w|5|poly
rlabel polysilicon -13 33 -9 36 1 _SReset!|pin|w|5|poly
rlabel polysilicon 51 61 55 64 1 _PReset!|pin|w|6|poly
rlabel polysilicon 67 61 71 64 1 _PReset!|pin|w|6|poly
<< end >>
