package mby_env_pkg;

`include "mby_defines.sv"

 
`ifdef XVM
   import ovm_pkg::*;
   import xvm_pkg::*;
   `include "ovm_macros.svh"
   `include "sla_macros.svh"
`endif

import sla_pkg::*;
import uvm_pkg::*;

import shdv_base_pkg::*;
import mby_wm_dpi_pkg::*;    
    
// START IOSF_NOT_PRESENT
// import svlib_pkg::*;
// import IosfPkg::*;    
// END IOSF_NOT_PRESENT

// START CHASSIS_NOT_PRESENT
// import PowerGatingCommonPkg::*;
// import CCAgentPkg::*;
// import chassis_reset_pkg::*;
// import ccu_vc_pkg::*;
// END CHASSIS_NOT_PRESENT

// START FUSE_NOT_PRESENT
// import sla_fusegen_pkg::*;
// END FUSE_NOT_PRESENT
  
`include "uvm_macros.svh"
`include "slu_macros.svh"
  
`include "mby_types.sv"
`include "mby_params.sv"
`include "mby_ti_config.sv"
`include "mby_config.sv"

// START IOSF_NOT_PRESENT
//`include "mby_pri_scbd.sv"
//`include "mby_ral_iosf_sb_access.sv"
//`include "mby_ral_iosf_pri_access.sv"
// END IOSF_NOT_PRESENT

`include "mby_ral_env.sv"
`include "mby_env_monitor.sv"
`include "mby_base_env.sv"
`include "mby_env.sv"
`include "mby_seqlib.sv"
`include "mby_sm_env.sv"
`include "mby_im_env.sv"

// START FUSE_NOT_PRESENT
//`include "mby_fuse_env.sv" // this is not reusable
// END FUSE_NOT_PRESENT
  
endpackage :mby_env_pkg
