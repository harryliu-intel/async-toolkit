///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_policers_map_pkg.vh                                
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_POLICERS_MAP_PKG_VH
`define MBY_PPE_POLICERS_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_policers_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_policers_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_policers_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_policers_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic  [0:0] GO_COMPL;  // RW/V
    logic  [0:0] STATUS;  // RW/V
    logic  [0:0] OP_TYPE;  // RW
    logic [12:0] reserved0;  // RSVD
    logic  [7:0] REG_ID;  // RW
    logic  [7:0] REG_SUB_ID;  // RW
    logic [31:0] REG_INDX;  // RW
} POL_DIRECT_MAP_CTRL_t;

localparam POL_DIRECT_MAP_CTRL_REG_STRIDE = 48'h8;
localparam POL_DIRECT_MAP_CTRL_REG_ENTRIES = 1;
localparam POL_DIRECT_MAP_CTRL_CR_ADDR = 48'h0;
localparam POL_DIRECT_MAP_CTRL_SIZE = 64;
localparam POL_DIRECT_MAP_CTRL_GO_COMPL_LO = 63;
localparam POL_DIRECT_MAP_CTRL_GO_COMPL_HI = 63;
localparam POL_DIRECT_MAP_CTRL_GO_COMPL_RESET = 1'h0;
localparam POL_DIRECT_MAP_CTRL_STATUS_LO = 62;
localparam POL_DIRECT_MAP_CTRL_STATUS_HI = 62;
localparam POL_DIRECT_MAP_CTRL_STATUS_RESET = 1'h0;
localparam POL_DIRECT_MAP_CTRL_OP_TYPE_LO = 61;
localparam POL_DIRECT_MAP_CTRL_OP_TYPE_HI = 61;
localparam POL_DIRECT_MAP_CTRL_OP_TYPE_RESET = 1'h0;
localparam POL_DIRECT_MAP_CTRL_REG_ID_LO = 40;
localparam POL_DIRECT_MAP_CTRL_REG_ID_HI = 47;
localparam POL_DIRECT_MAP_CTRL_REG_ID_RESET = 8'h0;
localparam POL_DIRECT_MAP_CTRL_REG_SUB_ID_LO = 32;
localparam POL_DIRECT_MAP_CTRL_REG_SUB_ID_HI = 39;
localparam POL_DIRECT_MAP_CTRL_REG_SUB_ID_RESET = 8'h0;
localparam POL_DIRECT_MAP_CTRL_REG_INDX_LO = 0;
localparam POL_DIRECT_MAP_CTRL_REG_INDX_HI = 31;
localparam POL_DIRECT_MAP_CTRL_REG_INDX_RESET = 32'h0;
localparam POL_DIRECT_MAP_CTRL_USEMASK = 64'hE000FFFFFFFFFFFF;
localparam POL_DIRECT_MAP_CTRL_RO_MASK = 64'h0;
localparam POL_DIRECT_MAP_CTRL_WO_MASK = 64'h0;
localparam POL_DIRECT_MAP_CTRL_RESET = 64'h0;

typedef struct packed {
    logic [19:0] reserved0;  // RSVD
    logic [43:0] DATA_CNTB;  // RW/V
} POL_DIRECT_MAP_CTR0_t;

localparam POL_DIRECT_MAP_CTR0_REG_STRIDE = 48'h8;
localparam POL_DIRECT_MAP_CTR0_REG_ENTRIES = 1;
localparam POL_DIRECT_MAP_CTR0_CR_ADDR = 48'h8;
localparam POL_DIRECT_MAP_CTR0_SIZE = 64;
localparam POL_DIRECT_MAP_CTR0_DATA_CNTB_LO = 0;
localparam POL_DIRECT_MAP_CTR0_DATA_CNTB_HI = 43;
localparam POL_DIRECT_MAP_CTR0_DATA_CNTB_RESET = 44'h0;
localparam POL_DIRECT_MAP_CTR0_USEMASK = 64'hFFFFFFFFFFF;
localparam POL_DIRECT_MAP_CTR0_RO_MASK = 64'h0;
localparam POL_DIRECT_MAP_CTR0_WO_MASK = 64'h0;
localparam POL_DIRECT_MAP_CTR0_RESET = 64'h0;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic [35:0] DATA_CNTP;  // RW/V
} POL_DIRECT_MAP_CTR1_t;

localparam POL_DIRECT_MAP_CTR1_REG_STRIDE = 48'h8;
localparam POL_DIRECT_MAP_CTR1_REG_ENTRIES = 1;
localparam POL_DIRECT_MAP_CTR1_CR_ADDR = 48'h10;
localparam POL_DIRECT_MAP_CTR1_SIZE = 64;
localparam POL_DIRECT_MAP_CTR1_DATA_CNTP_LO = 0;
localparam POL_DIRECT_MAP_CTR1_DATA_CNTP_HI = 35;
localparam POL_DIRECT_MAP_CTR1_DATA_CNTP_RESET = 36'h0;
localparam POL_DIRECT_MAP_CTR1_USEMASK = 64'hFFFFFFFFF;
localparam POL_DIRECT_MAP_CTR1_RO_MASK = 64'h0;
localparam POL_DIRECT_MAP_CTR1_WO_MASK = 64'h0;
localparam POL_DIRECT_MAP_CTR1_RESET = 64'h0;

typedef struct packed {
    logic [23:0] ETOK_HI;  // RW/V
    logic  [2:0] reserved0;  // RSVD
    logic [12:0] ETOK_LO;  // RW/V
    logic [23:0] TIME_STORED;  // RO/V
} POL_DIRECT_MAP_POL0_t;

localparam POL_DIRECT_MAP_POL0_REG_STRIDE = 48'h8;
localparam POL_DIRECT_MAP_POL0_REG_ENTRIES = 1;
localparam POL_DIRECT_MAP_POL0_CR_ADDR = 48'h18;
localparam POL_DIRECT_MAP_POL0_SIZE = 64;
localparam POL_DIRECT_MAP_POL0_ETOK_HI_LO = 40;
localparam POL_DIRECT_MAP_POL0_ETOK_HI_HI = 63;
localparam POL_DIRECT_MAP_POL0_ETOK_HI_RESET = 24'h0;
localparam POL_DIRECT_MAP_POL0_ETOK_LO_LO = 24;
localparam POL_DIRECT_MAP_POL0_ETOK_LO_HI = 36;
localparam POL_DIRECT_MAP_POL0_ETOK_LO_RESET = 13'h0;
localparam POL_DIRECT_MAP_POL0_TIME_STORED_LO = 0;
localparam POL_DIRECT_MAP_POL0_TIME_STORED_HI = 23;
localparam POL_DIRECT_MAP_POL0_TIME_STORED_RESET = 24'h0;
localparam POL_DIRECT_MAP_POL0_USEMASK = 64'hFFFFFF1FFFFFFFFF;
localparam POL_DIRECT_MAP_POL0_RO_MASK = 64'hFFFFFF;
localparam POL_DIRECT_MAP_POL0_WO_MASK = 64'h0;
localparam POL_DIRECT_MAP_POL0_RESET = 64'h0;

typedef struct packed {
    logic [23:0] CTOK_HI;  // RW/V
    logic  [2:0] reserved0;  // RSVD
    logic [12:0] CTOK_LO;  // RW/V
    logic [19:0] reserved1;  // RSVD
    logic  [3:0] CFG;  // RW
} POL_DIRECT_MAP_POL1_t;

localparam POL_DIRECT_MAP_POL1_REG_STRIDE = 48'h8;
localparam POL_DIRECT_MAP_POL1_REG_ENTRIES = 1;
localparam POL_DIRECT_MAP_POL1_CR_ADDR = 48'h20;
localparam POL_DIRECT_MAP_POL1_SIZE = 64;
localparam POL_DIRECT_MAP_POL1_CTOK_HI_LO = 40;
localparam POL_DIRECT_MAP_POL1_CTOK_HI_HI = 63;
localparam POL_DIRECT_MAP_POL1_CTOK_HI_RESET = 24'h0;
localparam POL_DIRECT_MAP_POL1_CTOK_LO_LO = 24;
localparam POL_DIRECT_MAP_POL1_CTOK_LO_HI = 36;
localparam POL_DIRECT_MAP_POL1_CTOK_LO_RESET = 13'h0;
localparam POL_DIRECT_MAP_POL1_CFG_LO = 0;
localparam POL_DIRECT_MAP_POL1_CFG_HI = 3;
localparam POL_DIRECT_MAP_POL1_CFG_RESET = 4'h0;
localparam POL_DIRECT_MAP_POL1_USEMASK = 64'hFFFFFF1FFF00000F;
localparam POL_DIRECT_MAP_POL1_RO_MASK = 64'h0;
localparam POL_DIRECT_MAP_POL1_WO_MASK = 64'h0;
localparam POL_DIRECT_MAP_POL1_RESET = 64'h0;

typedef struct packed {
    logic [33:0] reserved0;  // RSVD
    logic  [2:0] EIR_UNIT;  // RW
    logic [10:0] EIR;  // RW
    logic  [0:0] reserved1;  // RSVD
    logic  [1:0] EBS_UNIT;  // RW
    logic [12:0] EBS;  // RW
} POL_DIRECT_MAP_POL2_t;

localparam POL_DIRECT_MAP_POL2_REG_STRIDE = 48'h8;
localparam POL_DIRECT_MAP_POL2_REG_ENTRIES = 1;
localparam POL_DIRECT_MAP_POL2_CR_ADDR = 48'h28;
localparam POL_DIRECT_MAP_POL2_SIZE = 64;
localparam POL_DIRECT_MAP_POL2_EIR_UNIT_LO = 27;
localparam POL_DIRECT_MAP_POL2_EIR_UNIT_HI = 29;
localparam POL_DIRECT_MAP_POL2_EIR_UNIT_RESET = 3'h0;
localparam POL_DIRECT_MAP_POL2_EIR_LO = 16;
localparam POL_DIRECT_MAP_POL2_EIR_HI = 26;
localparam POL_DIRECT_MAP_POL2_EIR_RESET = 11'h0;
localparam POL_DIRECT_MAP_POL2_EBS_UNIT_LO = 13;
localparam POL_DIRECT_MAP_POL2_EBS_UNIT_HI = 14;
localparam POL_DIRECT_MAP_POL2_EBS_UNIT_RESET = 2'h0;
localparam POL_DIRECT_MAP_POL2_EBS_LO = 0;
localparam POL_DIRECT_MAP_POL2_EBS_HI = 12;
localparam POL_DIRECT_MAP_POL2_EBS_RESET = 13'h0;
localparam POL_DIRECT_MAP_POL2_USEMASK = 64'h3FFF7FFF;
localparam POL_DIRECT_MAP_POL2_RO_MASK = 64'h0;
localparam POL_DIRECT_MAP_POL2_WO_MASK = 64'h0;
localparam POL_DIRECT_MAP_POL2_RESET = 64'h0;

typedef struct packed {
    logic [33:0] reserved0;  // RSVD
    logic  [2:0] CIR_UNIT;  // RW
    logic [10:0] CIR;  // RW
    logic  [0:0] reserved1;  // RSVD
    logic  [1:0] CBS_UNIT;  // RW
    logic [12:0] CBS;  // RW
} POL_DIRECT_MAP_POL3_t;

localparam POL_DIRECT_MAP_POL3_REG_STRIDE = 48'h8;
localparam POL_DIRECT_MAP_POL3_REG_ENTRIES = 1;
localparam POL_DIRECT_MAP_POL3_CR_ADDR = 48'h30;
localparam POL_DIRECT_MAP_POL3_SIZE = 64;
localparam POL_DIRECT_MAP_POL3_CIR_UNIT_LO = 27;
localparam POL_DIRECT_MAP_POL3_CIR_UNIT_HI = 29;
localparam POL_DIRECT_MAP_POL3_CIR_UNIT_RESET = 3'h0;
localparam POL_DIRECT_MAP_POL3_CIR_LO = 16;
localparam POL_DIRECT_MAP_POL3_CIR_HI = 26;
localparam POL_DIRECT_MAP_POL3_CIR_RESET = 11'h0;
localparam POL_DIRECT_MAP_POL3_CBS_UNIT_LO = 13;
localparam POL_DIRECT_MAP_POL3_CBS_UNIT_HI = 14;
localparam POL_DIRECT_MAP_POL3_CBS_UNIT_RESET = 2'h0;
localparam POL_DIRECT_MAP_POL3_CBS_LO = 0;
localparam POL_DIRECT_MAP_POL3_CBS_HI = 12;
localparam POL_DIRECT_MAP_POL3_CBS_RESET = 13'h0;
localparam POL_DIRECT_MAP_POL3_USEMASK = 64'h3FFF7FFF;
localparam POL_DIRECT_MAP_POL3_RO_MASK = 64'h0;
localparam POL_DIRECT_MAP_POL3_WO_MASK = 64'h0;
localparam POL_DIRECT_MAP_POL3_RESET = 64'h0;

typedef struct packed {
    logic [40:0] reserved0;  // RSVD
    logic  [0:0] UNPOLICE_DROP_CM;  // RW
    logic  [0:0] UNPOLICE_DROP_PRECM;  // RW
    logic  [0:0] CREDIT_FRAME_ERR;  // RW
    logic  [0:0] CREDIT_L3_LEN_ERR;  // RW
    logic  [1:0] reserved1;  // RSVD
    logic  [0:0] CB;  // RW
    logic  [0:0] CF;  // RW
    logic  [0:0] COLOR_SELECT;  // RW
    logic  [0:0] PRECEDENCE;  // RW
    logic  [0:0] DEBIT_MODE;  // RW
    logic  [0:0] L3_LEN_MODE;  // RW
    logic [10:0] reserved2;  // RSVD
} POL_CFG_t;

localparam POL_CFG_REG_STRIDE = 48'h8;
localparam POL_CFG_REG_ENTRIES = 16;
localparam POL_CFG_REGFILE_STRIDE = 48'h80;
localparam POL_CFG_REGFILE_ENTRIES = 2;
localparam POL_CFG_CR_ADDR = 48'h40;
localparam POL_CFG_SIZE = 64;
localparam POL_CFG_UNPOLICE_DROP_CM_LO = 22;
localparam POL_CFG_UNPOLICE_DROP_CM_HI = 22;
localparam POL_CFG_UNPOLICE_DROP_CM_RESET = 1'h0;
localparam POL_CFG_UNPOLICE_DROP_PRECM_LO = 21;
localparam POL_CFG_UNPOLICE_DROP_PRECM_HI = 21;
localparam POL_CFG_UNPOLICE_DROP_PRECM_RESET = 1'h1;
localparam POL_CFG_CREDIT_FRAME_ERR_LO = 20;
localparam POL_CFG_CREDIT_FRAME_ERR_HI = 20;
localparam POL_CFG_CREDIT_FRAME_ERR_RESET = 1'h1;
localparam POL_CFG_CREDIT_L3_LEN_ERR_LO = 19;
localparam POL_CFG_CREDIT_L3_LEN_ERR_HI = 19;
localparam POL_CFG_CREDIT_L3_LEN_ERR_RESET = 1'h0;
localparam POL_CFG_CB_LO = 16;
localparam POL_CFG_CB_HI = 16;
localparam POL_CFG_CB_RESET = 1'h0;
localparam POL_CFG_CF_LO = 15;
localparam POL_CFG_CF_HI = 15;
localparam POL_CFG_CF_RESET = 1'h0;
localparam POL_CFG_COLOR_SELECT_LO = 14;
localparam POL_CFG_COLOR_SELECT_HI = 14;
localparam POL_CFG_COLOR_SELECT_RESET = 1'h0;
localparam POL_CFG_PRECEDENCE_LO = 13;
localparam POL_CFG_PRECEDENCE_HI = 13;
localparam POL_CFG_PRECEDENCE_RESET = 1'h0;
localparam POL_CFG_DEBIT_MODE_LO = 12;
localparam POL_CFG_DEBIT_MODE_HI = 12;
localparam POL_CFG_DEBIT_MODE_RESET = 1'h0;
localparam POL_CFG_L3_LEN_MODE_LO = 11;
localparam POL_CFG_L3_LEN_MODE_HI = 11;
localparam POL_CFG_L3_LEN_MODE_RESET = 1'h0;
localparam POL_CFG_USEMASK = 64'h79F800;
localparam POL_CFG_RO_MASK = 64'h0;
localparam POL_CFG_WO_MASK = 64'h0;
localparam POL_CFG_RESET = 64'h300000;

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic  [0:0] IR;  // RW
    logic  [0:0] IG;  // RW
    logic  [0:0] DROP_ER;  // RW
    logic  [5:0] TO_YELLOW;  // RW
    logic  [5:0] TO_RED;  // RW
} POL_DSCP_t;

localparam POL_DSCP_REG_STRIDE = 48'h8;
localparam POL_DSCP_REG_ENTRIES = 64;
localparam POL_DSCP_REGFILE_STRIDE = 48'h200;
localparam POL_DSCP_REGFILE_ENTRIES = 16;
localparam POL_DSCP_CR_ADDR = 48'h2040;
localparam POL_DSCP_SIZE = 64;
localparam POL_DSCP_IR_LO = 14;
localparam POL_DSCP_IR_HI = 14;
localparam POL_DSCP_IR_RESET = 1'h0;
localparam POL_DSCP_IG_LO = 13;
localparam POL_DSCP_IG_HI = 13;
localparam POL_DSCP_IG_RESET = 1'h0;
localparam POL_DSCP_DROP_ER_LO = 12;
localparam POL_DSCP_DROP_ER_HI = 12;
localparam POL_DSCP_DROP_ER_RESET = 1'h0;
localparam POL_DSCP_TO_YELLOW_LO = 6;
localparam POL_DSCP_TO_YELLOW_HI = 11;
localparam POL_DSCP_TO_YELLOW_RESET = 6'h0;
localparam POL_DSCP_TO_RED_LO = 0;
localparam POL_DSCP_TO_RED_HI = 5;
localparam POL_DSCP_TO_RED_RESET = 6'h0;
localparam POL_DSCP_USEMASK = 64'h7FFF;
localparam POL_DSCP_RO_MASK = 64'h0;
localparam POL_DSCP_WO_MASK = 64'h0;
localparam POL_DSCP_RESET = 64'h0;

typedef struct packed {
    logic [52:0] reserved0;  // RSVD
    logic  [0:0] IR;  // RW
    logic  [0:0] IG;  // RW
    logic  [0:0] DROP_ER;  // RW
    logic  [3:0] TO_YELLOW;  // RW
    logic  [3:0] TO_RED;  // RW
} POL_VPRI_t;

localparam POL_VPRI_REG_STRIDE = 48'h8;
localparam POL_VPRI_REG_ENTRIES = 16;
localparam POL_VPRI_REGFILE_STRIDE = 48'h80;
localparam POL_VPRI_REGFILE_ENTRIES = 16;
localparam POL_VPRI_CR_ADDR = 48'h4040;
localparam POL_VPRI_SIZE = 64;
localparam POL_VPRI_IR_LO = 10;
localparam POL_VPRI_IR_HI = 10;
localparam POL_VPRI_IR_RESET = 1'h0;
localparam POL_VPRI_IG_LO = 9;
localparam POL_VPRI_IG_HI = 9;
localparam POL_VPRI_IG_RESET = 1'h0;
localparam POL_VPRI_DROP_ER_LO = 8;
localparam POL_VPRI_DROP_ER_HI = 8;
localparam POL_VPRI_DROP_ER_RESET = 1'h0;
localparam POL_VPRI_TO_YELLOW_LO = 4;
localparam POL_VPRI_TO_YELLOW_HI = 7;
localparam POL_VPRI_TO_YELLOW_RESET = 4'h0;
localparam POL_VPRI_TO_RED_LO = 0;
localparam POL_VPRI_TO_RED_HI = 3;
localparam POL_VPRI_TO_RED_RESET = 4'h0;
localparam POL_VPRI_USEMASK = 64'h7FF;
localparam POL_VPRI_RO_MASK = 64'h0;
localparam POL_VPRI_WO_MASK = 64'h0;
localparam POL_VPRI_RESET = 64'h0;

typedef struct packed {
    logic [43:0] reserved0;  // RSVD
    logic [19:0] POL_TIME_UNIT;  // RW
} POL_TIME_UNIT_t;

localparam POL_TIME_UNIT_REG_STRIDE = 48'h8;
localparam POL_TIME_UNIT_REG_ENTRIES = 1;
localparam POL_TIME_UNIT_CR_ADDR = 48'h4840;
localparam POL_TIME_UNIT_SIZE = 64;
localparam POL_TIME_UNIT_POL_TIME_UNIT_LO = 0;
localparam POL_TIME_UNIT_POL_TIME_UNIT_HI = 19;
localparam POL_TIME_UNIT_POL_TIME_UNIT_RESET = 20'h0;
localparam POL_TIME_UNIT_USEMASK = 64'hFFFFF;
localparam POL_TIME_UNIT_RO_MASK = 64'h0;
localparam POL_TIME_UNIT_WO_MASK = 64'h0;
localparam POL_TIME_UNIT_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] POL_TIME;  // RW/V
} POL_TIME_t;

localparam POL_TIME_REG_STRIDE = 48'h8;
localparam POL_TIME_REG_ENTRIES = 1;
localparam POL_TIME_CR_ADDR = 48'h4848;
localparam POL_TIME_SIZE = 64;
localparam POL_TIME_POL_TIME_LO = 0;
localparam POL_TIME_POL_TIME_HI = 47;
localparam POL_TIME_POL_TIME_RESET = 48'h0;
localparam POL_TIME_USEMASK = 64'hFFFFFFFFFFFF;
localparam POL_TIME_RO_MASK = 64'h0;
localparam POL_TIME_WO_MASK = 64'h0;
localparam POL_TIME_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [15:0] ELAPSE_CYCLE;  // RW
    logic  [7:0] ELAPSE_SLOT;  // RW
    logic [11:0] POL0_HI;  // RW
    logic [11:0] POL1_HI;  // RW
} POL_SWEEP_t;

localparam POL_SWEEP_REG_STRIDE = 48'h8;
localparam POL_SWEEP_REG_ENTRIES = 1;
localparam POL_SWEEP_CR_ADDR = 48'h4850;
localparam POL_SWEEP_SIZE = 64;
localparam POL_SWEEP_ELAPSE_CYCLE_LO = 32;
localparam POL_SWEEP_ELAPSE_CYCLE_HI = 47;
localparam POL_SWEEP_ELAPSE_CYCLE_RESET = 16'h0;
localparam POL_SWEEP_ELAPSE_SLOT_LO = 24;
localparam POL_SWEEP_ELAPSE_SLOT_HI = 31;
localparam POL_SWEEP_ELAPSE_SLOT_RESET = 8'h0;
localparam POL_SWEEP_POL0_HI_LO = 12;
localparam POL_SWEEP_POL0_HI_HI = 23;
localparam POL_SWEEP_POL0_HI_RESET = 12'h0;
localparam POL_SWEEP_POL1_HI_LO = 0;
localparam POL_SWEEP_POL1_HI_HI = 11;
localparam POL_SWEEP_POL1_HI_RESET = 12'h0;
localparam POL_SWEEP_USEMASK = 64'hFFFFFFFFFFFF;
localparam POL_SWEEP_RO_MASK = 64'h0;
localparam POL_SWEEP_WO_MASK = 64'h0;
localparam POL_SWEEP_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] POL_SWEEP_LAST;  // RW/V
} POL_SWEEP_LAST_t;

localparam POL_SWEEP_LAST_REG_STRIDE = 48'h8;
localparam POL_SWEEP_LAST_REG_ENTRIES = 1;
localparam POL_SWEEP_LAST_CR_ADDR = 48'h4858;
localparam POL_SWEEP_LAST_SIZE = 64;
localparam POL_SWEEP_LAST_POL_SWEEP_LAST_LO = 0;
localparam POL_SWEEP_LAST_POL_SWEEP_LAST_HI = 47;
localparam POL_SWEEP_LAST_POL_SWEEP_LAST_RESET = 48'h0;
localparam POL_SWEEP_LAST_USEMASK = 64'hFFFFFFFFFFFF;
localparam POL_SWEEP_LAST_RO_MASK = 64'h0;
localparam POL_SWEEP_LAST_WO_MASK = 64'h0;
localparam POL_SWEEP_LAST_RESET = 64'h0;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] POL_SWEEP_PERIOD_MAX;  // RW/V
} POL_SWEEP_PERIOD_MAX_t;

localparam POL_SWEEP_PERIOD_MAX_REG_STRIDE = 48'h8;
localparam POL_SWEEP_PERIOD_MAX_REG_ENTRIES = 1;
localparam POL_SWEEP_PERIOD_MAX_CR_ADDR = 48'h4860;
localparam POL_SWEEP_PERIOD_MAX_SIZE = 64;
localparam POL_SWEEP_PERIOD_MAX_POL_SWEEP_PERIOD_MAX_LO = 0;
localparam POL_SWEEP_PERIOD_MAX_POL_SWEEP_PERIOD_MAX_HI = 47;
localparam POL_SWEEP_PERIOD_MAX_POL_SWEEP_PERIOD_MAX_RESET = 48'h0;
localparam POL_SWEEP_PERIOD_MAX_USEMASK = 64'hFFFFFFFFFFFF;
localparam POL_SWEEP_PERIOD_MAX_RO_MASK = 64'h0;
localparam POL_SWEEP_PERIOD_MAX_WO_MASK = 64'h0;
localparam POL_SWEEP_PERIOD_MAX_RESET = 64'h0;

// ===================================================
// load

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_POL_DIRECT_MAP_CTRL_t;

typedef logic [7:0] we_POL_DIRECT_MAP_CTR0_t;

typedef logic [7:0] we_POL_DIRECT_MAP_CTR1_t;

typedef logic [7:0] we_POL_DIRECT_MAP_POL0_t;

typedef logic [7:0] we_POL_DIRECT_MAP_POL1_t;

typedef logic [7:0] we_POL_DIRECT_MAP_POL2_t;

typedef logic [7:0] we_POL_DIRECT_MAP_POL3_t;

typedef logic [7:0] we_POL_CFG_t;

typedef logic [7:0] we_POL_DSCP_t;

typedef logic [7:0] we_POL_VPRI_t;

typedef logic [7:0] we_POL_TIME_UNIT_t;

typedef logic [7:0] we_POL_TIME_t;

typedef logic [7:0] we_POL_SWEEP_t;

typedef logic [7:0] we_POL_SWEEP_LAST_t;

typedef logic [7:0] we_POL_SWEEP_PERIOD_MAX_t;

typedef struct packed {
    we_POL_DIRECT_MAP_CTRL_t POL_DIRECT_MAP_CTRL;
    we_POL_DIRECT_MAP_CTR0_t POL_DIRECT_MAP_CTR0;
    we_POL_DIRECT_MAP_CTR1_t POL_DIRECT_MAP_CTR1;
    we_POL_DIRECT_MAP_POL0_t POL_DIRECT_MAP_POL0;
    we_POL_DIRECT_MAP_POL1_t POL_DIRECT_MAP_POL1;
    we_POL_DIRECT_MAP_POL2_t POL_DIRECT_MAP_POL2;
    we_POL_DIRECT_MAP_POL3_t POL_DIRECT_MAP_POL3;
    we_POL_CFG_t POL_CFG;
    we_POL_DSCP_t POL_DSCP;
    we_POL_VPRI_t POL_VPRI;
    we_POL_TIME_UNIT_t POL_TIME_UNIT;
    we_POL_TIME_t POL_TIME;
    we_POL_SWEEP_t POL_SWEEP;
    we_POL_SWEEP_LAST_t POL_SWEEP_LAST;
    we_POL_SWEEP_PERIOD_MAX_t POL_SWEEP_PERIOD_MAX;
} mby_ppe_policers_map_handcoded_t;

typedef logic [7:0] re_POL_DIRECT_MAP_CTRL_t;

typedef logic [7:0] re_POL_DIRECT_MAP_CTR0_t;

typedef logic [7:0] re_POL_DIRECT_MAP_CTR1_t;

typedef logic [7:0] re_POL_DIRECT_MAP_POL0_t;

typedef logic [7:0] re_POL_DIRECT_MAP_POL1_t;

typedef logic [7:0] re_POL_DIRECT_MAP_POL2_t;

typedef logic [7:0] re_POL_DIRECT_MAP_POL3_t;

typedef logic [7:0] re_POL_CFG_t;

typedef logic [7:0] re_POL_DSCP_t;

typedef logic [7:0] re_POL_VPRI_t;

typedef logic [7:0] re_POL_TIME_UNIT_t;

typedef logic [7:0] re_POL_TIME_t;

typedef logic [7:0] re_POL_SWEEP_t;

typedef logic [7:0] re_POL_SWEEP_LAST_t;

typedef logic [7:0] re_POL_SWEEP_PERIOD_MAX_t;

typedef struct packed {
    re_POL_DIRECT_MAP_CTRL_t POL_DIRECT_MAP_CTRL;
    re_POL_DIRECT_MAP_CTR0_t POL_DIRECT_MAP_CTR0;
    re_POL_DIRECT_MAP_CTR1_t POL_DIRECT_MAP_CTR1;
    re_POL_DIRECT_MAP_POL0_t POL_DIRECT_MAP_POL0;
    re_POL_DIRECT_MAP_POL1_t POL_DIRECT_MAP_POL1;
    re_POL_DIRECT_MAP_POL2_t POL_DIRECT_MAP_POL2;
    re_POL_DIRECT_MAP_POL3_t POL_DIRECT_MAP_POL3;
    re_POL_CFG_t POL_CFG;
    re_POL_DSCP_t POL_DSCP;
    re_POL_VPRI_t POL_VPRI;
    re_POL_TIME_UNIT_t POL_TIME_UNIT;
    re_POL_TIME_t POL_TIME;
    re_POL_SWEEP_t POL_SWEEP;
    re_POL_SWEEP_LAST_t POL_SWEEP_LAST;
    re_POL_SWEEP_PERIOD_MAX_t POL_SWEEP_PERIOD_MAX;
} mby_ppe_policers_map_hc_re_t;

typedef logic handcode_rvalid_POL_DIRECT_MAP_CTRL_t;

typedef logic handcode_rvalid_POL_DIRECT_MAP_CTR0_t;

typedef logic handcode_rvalid_POL_DIRECT_MAP_CTR1_t;

typedef logic handcode_rvalid_POL_DIRECT_MAP_POL0_t;

typedef logic handcode_rvalid_POL_DIRECT_MAP_POL1_t;

typedef logic handcode_rvalid_POL_DIRECT_MAP_POL2_t;

typedef logic handcode_rvalid_POL_DIRECT_MAP_POL3_t;

typedef logic handcode_rvalid_POL_CFG_t;

typedef logic handcode_rvalid_POL_DSCP_t;

typedef logic handcode_rvalid_POL_VPRI_t;

typedef logic handcode_rvalid_POL_TIME_UNIT_t;

typedef logic handcode_rvalid_POL_TIME_t;

typedef logic handcode_rvalid_POL_SWEEP_t;

typedef logic handcode_rvalid_POL_SWEEP_LAST_t;

typedef logic handcode_rvalid_POL_SWEEP_PERIOD_MAX_t;

typedef struct packed {
    handcode_rvalid_POL_DIRECT_MAP_CTRL_t POL_DIRECT_MAP_CTRL;
    handcode_rvalid_POL_DIRECT_MAP_CTR0_t POL_DIRECT_MAP_CTR0;
    handcode_rvalid_POL_DIRECT_MAP_CTR1_t POL_DIRECT_MAP_CTR1;
    handcode_rvalid_POL_DIRECT_MAP_POL0_t POL_DIRECT_MAP_POL0;
    handcode_rvalid_POL_DIRECT_MAP_POL1_t POL_DIRECT_MAP_POL1;
    handcode_rvalid_POL_DIRECT_MAP_POL2_t POL_DIRECT_MAP_POL2;
    handcode_rvalid_POL_DIRECT_MAP_POL3_t POL_DIRECT_MAP_POL3;
    handcode_rvalid_POL_CFG_t POL_CFG;
    handcode_rvalid_POL_DSCP_t POL_DSCP;
    handcode_rvalid_POL_VPRI_t POL_VPRI;
    handcode_rvalid_POL_TIME_UNIT_t POL_TIME_UNIT;
    handcode_rvalid_POL_TIME_t POL_TIME;
    handcode_rvalid_POL_SWEEP_t POL_SWEEP;
    handcode_rvalid_POL_SWEEP_LAST_t POL_SWEEP_LAST;
    handcode_rvalid_POL_SWEEP_PERIOD_MAX_t POL_SWEEP_PERIOD_MAX;
} mby_ppe_policers_map_hc_rvalid_t;

typedef logic handcode_wvalid_POL_DIRECT_MAP_CTRL_t;

typedef logic handcode_wvalid_POL_DIRECT_MAP_CTR0_t;

typedef logic handcode_wvalid_POL_DIRECT_MAP_CTR1_t;

typedef logic handcode_wvalid_POL_DIRECT_MAP_POL0_t;

typedef logic handcode_wvalid_POL_DIRECT_MAP_POL1_t;

typedef logic handcode_wvalid_POL_DIRECT_MAP_POL2_t;

typedef logic handcode_wvalid_POL_DIRECT_MAP_POL3_t;

typedef logic handcode_wvalid_POL_CFG_t;

typedef logic handcode_wvalid_POL_DSCP_t;

typedef logic handcode_wvalid_POL_VPRI_t;

typedef logic handcode_wvalid_POL_TIME_UNIT_t;

typedef logic handcode_wvalid_POL_TIME_t;

typedef logic handcode_wvalid_POL_SWEEP_t;

typedef logic handcode_wvalid_POL_SWEEP_LAST_t;

typedef logic handcode_wvalid_POL_SWEEP_PERIOD_MAX_t;

typedef struct packed {
    handcode_wvalid_POL_DIRECT_MAP_CTRL_t POL_DIRECT_MAP_CTRL;
    handcode_wvalid_POL_DIRECT_MAP_CTR0_t POL_DIRECT_MAP_CTR0;
    handcode_wvalid_POL_DIRECT_MAP_CTR1_t POL_DIRECT_MAP_CTR1;
    handcode_wvalid_POL_DIRECT_MAP_POL0_t POL_DIRECT_MAP_POL0;
    handcode_wvalid_POL_DIRECT_MAP_POL1_t POL_DIRECT_MAP_POL1;
    handcode_wvalid_POL_DIRECT_MAP_POL2_t POL_DIRECT_MAP_POL2;
    handcode_wvalid_POL_DIRECT_MAP_POL3_t POL_DIRECT_MAP_POL3;
    handcode_wvalid_POL_CFG_t POL_CFG;
    handcode_wvalid_POL_DSCP_t POL_DSCP;
    handcode_wvalid_POL_VPRI_t POL_VPRI;
    handcode_wvalid_POL_TIME_UNIT_t POL_TIME_UNIT;
    handcode_wvalid_POL_TIME_t POL_TIME;
    handcode_wvalid_POL_SWEEP_t POL_SWEEP;
    handcode_wvalid_POL_SWEEP_LAST_t POL_SWEEP_LAST;
    handcode_wvalid_POL_SWEEP_PERIOD_MAX_t POL_SWEEP_PERIOD_MAX;
} mby_ppe_policers_map_hc_wvalid_t;

typedef logic handcode_error_POL_DIRECT_MAP_CTRL_t;

typedef logic handcode_error_POL_DIRECT_MAP_CTR0_t;

typedef logic handcode_error_POL_DIRECT_MAP_CTR1_t;

typedef logic handcode_error_POL_DIRECT_MAP_POL0_t;

typedef logic handcode_error_POL_DIRECT_MAP_POL1_t;

typedef logic handcode_error_POL_DIRECT_MAP_POL2_t;

typedef logic handcode_error_POL_DIRECT_MAP_POL3_t;

typedef logic handcode_error_POL_CFG_t;

typedef logic handcode_error_POL_DSCP_t;

typedef logic handcode_error_POL_VPRI_t;

typedef logic handcode_error_POL_TIME_UNIT_t;

typedef logic handcode_error_POL_TIME_t;

typedef logic handcode_error_POL_SWEEP_t;

typedef logic handcode_error_POL_SWEEP_LAST_t;

typedef logic handcode_error_POL_SWEEP_PERIOD_MAX_t;

typedef struct packed {
    handcode_error_POL_DIRECT_MAP_CTRL_t POL_DIRECT_MAP_CTRL;
    handcode_error_POL_DIRECT_MAP_CTR0_t POL_DIRECT_MAP_CTR0;
    handcode_error_POL_DIRECT_MAP_CTR1_t POL_DIRECT_MAP_CTR1;
    handcode_error_POL_DIRECT_MAP_POL0_t POL_DIRECT_MAP_POL0;
    handcode_error_POL_DIRECT_MAP_POL1_t POL_DIRECT_MAP_POL1;
    handcode_error_POL_DIRECT_MAP_POL2_t POL_DIRECT_MAP_POL2;
    handcode_error_POL_DIRECT_MAP_POL3_t POL_DIRECT_MAP_POL3;
    handcode_error_POL_CFG_t POL_CFG;
    handcode_error_POL_DSCP_t POL_DSCP;
    handcode_error_POL_VPRI_t POL_VPRI;
    handcode_error_POL_TIME_UNIT_t POL_TIME_UNIT;
    handcode_error_POL_TIME_t POL_TIME;
    handcode_error_POL_SWEEP_t POL_SWEEP;
    handcode_error_POL_SWEEP_LAST_t POL_SWEEP_LAST;
    handcode_error_POL_SWEEP_PERIOD_MAX_t POL_SWEEP_PERIOD_MAX;
} mby_ppe_policers_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    POL_DIRECT_MAP_CTRL_t POL_DIRECT_MAP_CTRL;
    POL_DIRECT_MAP_CTR0_t POL_DIRECT_MAP_CTR0;
    POL_DIRECT_MAP_CTR1_t POL_DIRECT_MAP_CTR1;
    POL_DIRECT_MAP_POL0_t POL_DIRECT_MAP_POL0;
    POL_DIRECT_MAP_POL1_t POL_DIRECT_MAP_POL1;
    POL_DIRECT_MAP_POL2_t POL_DIRECT_MAP_POL2;
    POL_DIRECT_MAP_POL3_t POL_DIRECT_MAP_POL3;
    POL_CFG_t POL_CFG;
    POL_DSCP_t POL_DSCP;
    POL_VPRI_t POL_VPRI;
    POL_TIME_UNIT_t POL_TIME_UNIT;
    POL_TIME_t POL_TIME;
    POL_SWEEP_t POL_SWEEP;
    POL_SWEEP_LAST_t POL_SWEEP_LAST;
    POL_SWEEP_PERIOD_MAX_t POL_SWEEP_PERIOD_MAX;
} mby_ppe_policers_map_hc_reg_read_t;

typedef struct packed {
    POL_DIRECT_MAP_CTRL_t POL_DIRECT_MAP_CTRL;
    POL_DIRECT_MAP_CTR0_t POL_DIRECT_MAP_CTR0;
    POL_DIRECT_MAP_CTR1_t POL_DIRECT_MAP_CTR1;
    POL_DIRECT_MAP_POL0_t POL_DIRECT_MAP_POL0;
    POL_DIRECT_MAP_POL1_t POL_DIRECT_MAP_POL1;
    POL_DIRECT_MAP_POL2_t POL_DIRECT_MAP_POL2;
    POL_DIRECT_MAP_POL3_t POL_DIRECT_MAP_POL3;
    POL_CFG_t POL_CFG;
    POL_DSCP_t POL_DSCP;
    POL_VPRI_t POL_VPRI;
    POL_TIME_UNIT_t POL_TIME_UNIT;
    POL_TIME_t POL_TIME;
    POL_SWEEP_t POL_SWEEP;
    POL_SWEEP_LAST_t POL_SWEEP_LAST;
    POL_SWEEP_PERIOD_MAX_t POL_SWEEP_PERIOD_MAX;
} mby_ppe_policers_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_policers_map_pkg

`endif // MBY_PPE_POLICERS_MAP_PKG_VH
