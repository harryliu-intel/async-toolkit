magic
tech scmos
timestamp 969760391
<< ndiffusion >>
rect -57 67 -49 68
rect -57 63 -49 64
rect -57 54 -49 55
rect -57 50 -49 51
rect -57 28 -49 29
rect -57 20 -49 25
rect -57 16 -49 17
rect -57 7 -49 8
rect -57 3 -49 4
rect -57 -6 -49 -5
rect -57 -10 -49 -9
<< pdiffusion >>
rect -33 62 -25 63
rect -33 54 -25 59
rect -33 50 -25 51
rect -33 33 -25 34
rect -33 29 -25 30
rect -33 20 -25 21
rect -33 16 -25 17
rect -33 7 -25 8
rect -33 -1 -25 4
rect -33 -5 -25 -4
<< ntransistor >>
rect -57 64 -49 67
rect -57 51 -49 54
rect -57 25 -49 28
rect -57 17 -49 20
rect -57 4 -49 7
rect -57 -9 -49 -6
<< ptransistor >>
rect -33 59 -25 62
rect -33 51 -25 54
rect -33 30 -25 33
rect -33 17 -25 20
rect -33 4 -25 7
rect -33 -4 -25 -1
<< polysilicon >>
rect -61 64 -57 67
rect -49 64 -44 67
rect -47 62 -44 64
rect -47 59 -33 62
rect -25 59 -21 62
rect -61 51 -57 54
rect -49 51 -33 54
rect -25 51 -21 54
rect -40 33 -37 38
rect -40 30 -33 33
rect -25 30 -21 33
rect -40 28 -37 30
rect -61 25 -57 28
rect -49 25 -37 28
rect -61 17 -57 20
rect -49 17 -45 20
rect -37 17 -33 20
rect -25 17 -21 20
rect -61 4 -57 7
rect -49 4 -33 7
rect -25 4 -21 7
rect -47 -4 -33 -1
rect -25 -4 -21 -1
rect -47 -6 -44 -4
rect -61 -9 -57 -6
rect -49 -9 -44 -6
<< ndcontact >>
rect -57 68 -49 76
rect -57 55 -49 63
rect -57 42 -49 50
rect -57 29 -49 37
rect -57 8 -49 16
rect -57 -5 -49 3
rect -57 -18 -49 -10
<< pdcontact >>
rect -33 63 -25 71
rect -33 34 -25 50
rect -33 21 -25 29
rect -33 8 -25 16
rect -33 -13 -25 -5
<< polycontact >>
rect -45 38 -37 46
rect -45 12 -37 20
<< metal1 >>
rect -57 68 -49 76
rect -33 63 -25 71
rect -57 59 -29 63
rect -57 55 -49 59
rect -57 42 -49 50
rect -43 46 -39 59
rect -45 38 -37 46
rect -57 29 -49 37
rect -33 34 -25 50
rect -53 25 -25 29
rect -33 21 -25 25
rect -57 8 -49 16
rect -45 12 -37 20
rect -57 -1 -49 3
rect -43 -1 -39 12
rect -33 8 -25 16
rect -57 -5 -29 -1
rect -57 -18 -49 -10
rect -33 -13 -25 -5
<< labels >>
rlabel metal1 -53 46 -53 46 1 GND!
rlabel metal1 -53 72 -53 72 5 GND!
rlabel polysilicon -58 52 -58 52 3 a2
rlabel polysilicon -24 52 -24 52 7 a2
rlabel polysilicon -24 60 -24 60 7 a3
rlabel polysilicon -58 65 -58 65 3 a3
rlabel metal1 -53 59 -53 59 1 _a_23
rlabel metal1 -53 33 -53 33 1 av
rlabel metal1 -29 25 -29 25 1 av
rlabel metal1 -53 -1 -53 -1 1 _a_01
rlabel polysilicon -24 -3 -24 -3 7 a0
rlabel polysilicon -24 5 -24 5 7 a1
rlabel polysilicon -58 5 -58 5 3 a1
rlabel polysilicon -58 -8 -58 -8 3 a0
rlabel metal1 -29 12 -29 12 5 Vdd!
rlabel metal1 -53 -14 -53 -14 1 GND!
rlabel metal1 -53 12 -53 12 5 GND!
rlabel metal1 -29 42 -29 42 1 Vdd!
rlabel space -62 -18 -57 11 7 ^n01
rlabel space -25 -13 -20 9 3 ^p01
rlabel space -62 15 -57 30 7 ^n03
rlabel space -25 15 -20 35 3 ^p03
rlabel space -25 49 -20 64 3 ^p23
rlabel space -62 42 -57 76 7 ^n23
<< end >>
