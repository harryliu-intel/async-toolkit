///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Jon Bagge <jon.bagge.com> 
// -- Project Name : MBY 
// -- Description  : rx_ppe netlist. 
// ------------------------------------------------------------------- 

module rx_ppe (
rx_ppe_ppe_stm_if.ppe rx_ppe_ppe_stm_if, 
rx_ppe_igr_if.ppe rx_ppe_igr_if, 
//Input List
input                   cclk,                                     
input                   reset,                                    

//Interface List
ahb_rx_ppe_if.ppe                 ahb_rx_ppe_if,  
glb_rx_ppe_if.ppe                 glb_rx_ppe_if,  
igr_rx_ppe_if.ppe                 igr_rx_ppe_if   
);



// module parser_top    from parser_top using parser_top.map 
parser_top    parser_top(
/* input  logic                */ .reset         (reset),             
/* Interface ahb_rx_ppe_if.ppe */ .ahb_rx_ppe_if (ahb_rx_ppe_if),     
/* Interface glb_rx_ppe_if.ppe */ .glb_rx_ppe_if (glb_rx_ppe_if),     
/* Interface igr_rx_ppe_if.ppe */ .igr_rx_ppe_if (igr_rx_ppe_if),     
/* input  logic                */ .cclk          (cclk));              
// End of module parser_top from parser_top

endmodule // rx_ppe
