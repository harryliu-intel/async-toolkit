//-----------------------------------------------------------------------------
// Title         : Egress types
// Project       : Madison Bay
//-----------------------------------------------------------------------------
// File          : egress_types.svh
// Author        : jose.j.godinez.carrillo  <jjgodine@ichips.intel.com>
// Created       : 21.08.2018
// Last modified : 21.08.2018
//-----------------------------------------------------------------------------
// Description :
// Type definitions for egress cte
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by Intel Corporation This model is the confidential and
// proprietary property of Intel Corporation and the possession or use of this
// file requires a written license from Intel Corporation.
//------------------------------------------------------------------------------
// Modification history :
// 21.08.2018 : created
//-----------------------------------------------------------------------------
`ifndef EGRESS_TYPES_SV
`define EGRESS_TYPES_SV


`endif // EGRESS_TYPES_SV

