// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

//                                                                             
// File:       mby_regs_regs.svh                                               
// Creator:    romanb                                                          
// Time:       Monday Sep 16, 2013 [12:53:28 am]                               
//                                                                             
// Path:       /tmp/romanb/nebulon_run/31199                                   
// Arguments:  /p/com/eda/denali/blueprint/3.7.4/Linux/blueprint -html -I      
//             /p/com/eda/intel/nebulon/2.06p1/include -I source/rdl/ -ovm     
//             mby_ip.rdl                                                      
//                                                                             
// Sources:    /tmp/romanb/nebulon_run/31199/mby_cfg.rdl                       
//             /tmp/romanb/nebulon_run/31199/lib_udp.rdl                       
//             /tmp/romanb/nebulon_run/31199/mby_ip.rdl                        
//             /tmp/romanb/nebulon_run/31199/mby_mem.rdl                       
//             /p/com/eda/intel/nebulon/2.06p1/generators/html.pm              
//             /p/com/eda/intel/nebulon/2.06p1/generators/ovm.pm               
//             /p/com/eda/intel/nebulon/2.06p1/generators/generator_common.pm  
//                                                                             
// Blueprint:   3.7.4 (Tue Jun 23 00:17:01 PDT 2009)                           
// Machine:    icsl0407                                                        
// OS:         Linux 2.6.16.60-0.58.1.3835.0.PTF.638363-smp                    
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2013 Denali Software Inc.  All rights reserved                
// THIS FILE IS AUTOMATICALLY GENERATED BY DENALI BLUEPRINT, DO NOT EDIT       
//                                                                             


//RAL code compatible with Saola versions: v20130603 and newer 

`ifndef RAL_MBY_REGS_FILE
`define RAL_MBY_REGS_FILE

class mby_regs_DEVVENDID_reg extends sla_ral_reg;

  // --------------------------
  sla_ral_field VENDORID;
  sla_ral_field DEVICEID;

  // --------------------------
  `ovm_object_utils(mby_regs_DEVVENDID_reg)

  // --------------------------
  function new(
                string         name = "",
                `ifdef SLA_RAL_COVERAGE
                slu_ral_coverage_t cov_t = COVERAGE_OFF,
                `endif
                int            bus_num=0,
                int            dev_num=0,
                int            func_num=0,
                int            offset=0,
                int            size=0,
                slu_ral_data_t reset_val=0,
                boolean_t      mon_enabled = SLA_FALSE
             );
      super.new();
      set_space_addr("CFG",undef);
      set_space_addr("MEM",undef);
      set_space_addr("IO",undef);
      set_space_addr("MSG",undef);
      set_space_addr("CREG",undef); 
      set_space_addr("LT_MEM",undef);     

      build();

      `ifdef SLA_RAL_COVERAGE
      `CONFIG_RAL_COVERAGE(regname, COVERAGE_ON, FD_RW_SAMPLE)
      if(_coverage_type != COVERAGE_OFF) begin
        if(_sample_type inside {FD_RO_SAMPLE, RO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_WRITE)
        else if(_sample_type inside {FD_WO_SAMPLE, WO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_READ)
        else
        `CREATE_OP_SAMPLE_COV(RAL_NONE)
        `CREATE_DESIRED_COV
        `CREATE_ACTUAL_COV
      end
      `endif

  endfunction

  `ifdef SLA_RAL_COVERAGE
  `CREATE_RAL_OP_COVERGROUP
  covergroup desired_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(VENDORID, VENDORID.desired)
     `RAL_FIELD_CP_16(VENDORID, VENDORID.desired, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
     `RAL_FIELD_CP(DEVICEID, DEVICEID.desired)
     `RAL_FIELD_CP_16(DEVICEID, DEVICEID.desired, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
  endgroup

  covergroup actual_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(VENDORID, VENDORID.actual)
     `RAL_FIELD_CP_16(VENDORID, VENDORID.actual, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
     `RAL_FIELD_CP(DEVICEID, DEVICEID.actual)
     `RAL_FIELD_CP_16(DEVICEID, DEVICEID.actual, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
  endgroup
  `endif

  // --------------------------
  // add constraint based on database legal values
  // --------------------------
  function void build();
    VENDORID = new("VENDORID", "RW", 16, 0, {""});
    VENDORID.set_rand_mode(0);
    void'(add_field( VENDORID ));

    DEVICEID = new("DEVICEID", "RW", 16, 16, {""});
    DEVICEID.set_rand_mode(0);
    void'(add_field( DEVICEID ));

  endfunction

endclass : mby_regs_DEVVENDID_reg

// ================================================

class mby_regs_BASE_ADDR_0_reg extends sla_ral_reg;

  // --------------------------
  sla_ral_field MEMORY_IO_SPACE;
  sla_ral_field MEMORY_TYPE;
  sla_ral_field PREFETCHABLE_MEMORY;
  sla_ral_field MEMORY_SIZE;
  sla_ral_field BASE_ADDR;

  // --------------------------
  `ovm_object_utils(mby_regs_BASE_ADDR_0_reg)

  // --------------------------
  function new(
                string         name = "",
                `ifdef SLA_RAL_COVERAGE
                slu_ral_coverage_t cov_t = COVERAGE_OFF,
                `endif
                int            bus_num=0,
                int            dev_num=0,
                int            func_num=0,
                int            offset=0,
                int            size=0,
                slu_ral_data_t reset_val=0,
                boolean_t      mon_enabled = SLA_FALSE
             );
      super.new();
      set_space_addr("CFG",undef);
      set_space_addr("MEM",undef);
      set_space_addr("IO",undef);
      set_space_addr("MSG",undef);
      set_space_addr("CREG",undef); 
      set_space_addr("LT_MEM",undef);     

      build();

      `ifdef SLA_RAL_COVERAGE
      `CONFIG_RAL_COVERAGE(regname, COVERAGE_ON, FD_RW_SAMPLE)
      if(_coverage_type != COVERAGE_OFF) begin
        if(_sample_type inside {FD_RO_SAMPLE, RO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_WRITE)
        else if(_sample_type inside {FD_WO_SAMPLE, WO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_READ)
        else
        `CREATE_OP_SAMPLE_COV(RAL_NONE)
        `CREATE_DESIRED_COV
        `CREATE_ACTUAL_COV
      end
      `endif

  endfunction

  `ifdef SLA_RAL_COVERAGE
  `CREATE_RAL_OP_COVERGROUP
  covergroup desired_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(MEMORY_IO_SPACE, MEMORY_IO_SPACE.desired)
     `RAL_FIELD_CP_1(MEMORY_IO_SPACE, MEMORY_IO_SPACE.desired, 0)
     `RAL_FIELD_CP(MEMORY_TYPE, MEMORY_TYPE.desired)
     `RAL_FIELD_CP_2(MEMORY_TYPE, MEMORY_TYPE.desired, 0,1)
     `RAL_FIELD_CP(PREFETCHABLE_MEMORY, PREFETCHABLE_MEMORY.desired)
     `RAL_FIELD_CP_1(PREFETCHABLE_MEMORY, PREFETCHABLE_MEMORY.desired, 0)
     `RAL_FIELD_CP(MEMORY_SIZE, MEMORY_SIZE.desired)
     `RAL_FIELD_CP_13(MEMORY_SIZE, MEMORY_SIZE.desired, 0,1,2,3,4,5,6,7,8,9,10,11,12)
     `RAL_FIELD_CP(BASE_ADDR, BASE_ADDR.desired)
     `RAL_FIELD_CP_15(BASE_ADDR, BASE_ADDR.desired, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14)
  endgroup

  covergroup actual_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(MEMORY_IO_SPACE, MEMORY_IO_SPACE.actual)
     `RAL_FIELD_CP_1(MEMORY_IO_SPACE, MEMORY_IO_SPACE.actual, 0)
     `RAL_FIELD_CP(MEMORY_TYPE, MEMORY_TYPE.actual)
     `RAL_FIELD_CP_2(MEMORY_TYPE, MEMORY_TYPE.actual, 0,1)
     `RAL_FIELD_CP(PREFETCHABLE_MEMORY, PREFETCHABLE_MEMORY.actual)
     `RAL_FIELD_CP_1(PREFETCHABLE_MEMORY, PREFETCHABLE_MEMORY.actual, 0)
     `RAL_FIELD_CP(MEMORY_SIZE, MEMORY_SIZE.actual)
     `RAL_FIELD_CP_13(MEMORY_SIZE, MEMORY_SIZE.actual, 0,1,2,3,4,5,6,7,8,9,10,11,12)
     `RAL_FIELD_CP(BASE_ADDR, BASE_ADDR.actual)
     `RAL_FIELD_CP_15(BASE_ADDR, BASE_ADDR.actual, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14)
  endgroup
  `endif

  // --------------------------
  // add constraint based on database legal values
  // --------------------------
  function void build();
    MEMORY_IO_SPACE = new("MEMORY_IO_SPACE", "RO", 1, 0, {""});
    MEMORY_IO_SPACE.set_rand_mode(0);
    void'(add_field( MEMORY_IO_SPACE ));

    MEMORY_TYPE = new("MEMORY_TYPE", "RO", 2, 1, {""});
    MEMORY_TYPE.set_rand_mode(0);
    void'(add_field( MEMORY_TYPE ));

    PREFETCHABLE_MEMORY = new("PREFETCHABLE_MEMORY", "RO", 1, 3, {""});
    PREFETCHABLE_MEMORY.set_rand_mode(0);
    void'(add_field( PREFETCHABLE_MEMORY ));

    MEMORY_SIZE = new("MEMORY_SIZE", "RO", 13, 4, {""});
    MEMORY_SIZE.set_rand_mode(0);
    void'(add_field( MEMORY_SIZE ));

    BASE_ADDR = new("BASE_ADDR", "RW", 15, 17, {""});
    BASE_ADDR.set_rand_mode(0);
    void'(add_field( BASE_ADDR ));

  endfunction

endclass : mby_regs_BASE_ADDR_0_reg

// ================================================

class mby_regs_MEM_reg extends sla_ral_reg;

  // --------------------------
  sla_ral_field MEM2;
  sla_ral_field MEM1;

  // --------------------------
  `ovm_object_utils(mby_regs_MEM_reg)

  // --------------------------
  function new(
                string         name = "",
                `ifdef SLA_RAL_COVERAGE
                slu_ral_coverage_t cov_t = COVERAGE_OFF,
                `endif
                int            bus_num=0,
                int            dev_num=0,
                int            func_num=0,
                int            offset=0,
                int            size=0,
                slu_ral_data_t reset_val=0,
                boolean_t      mon_enabled = SLA_FALSE
             );
      super.new();
      set_space_addr("CFG",undef);
      set_space_addr("MEM",undef);
      set_space_addr("IO",undef);
      set_space_addr("MSG",undef);
      set_space_addr("CREG",undef); 
      set_space_addr("LT_MEM",undef);     

      build();

      `ifdef SLA_RAL_COVERAGE
      `CONFIG_RAL_COVERAGE(regname, COVERAGE_ON, FD_RW_SAMPLE)
      if(_coverage_type != COVERAGE_OFF) begin
        if(_sample_type inside {FD_RO_SAMPLE, RO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_WRITE)
        else if(_sample_type inside {FD_WO_SAMPLE, WO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_READ)
        else
        `CREATE_OP_SAMPLE_COV(RAL_NONE)
        `CREATE_DESIRED_COV
        `CREATE_ACTUAL_COV
      end
      `endif

  endfunction

  `ifdef SLA_RAL_COVERAGE
  `CREATE_RAL_OP_COVERGROUP
  covergroup desired_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(MEM2, MEM2.desired)
     `RAL_FIELD_CP_16(MEM2, MEM2.desired, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
     `RAL_FIELD_CP(MEM1, MEM1.desired)
     `RAL_FIELD_CP_16(MEM1, MEM1.desired, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
  endgroup

  covergroup actual_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(MEM2, MEM2.actual)
     `RAL_FIELD_CP_16(MEM2, MEM2.actual, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
     `RAL_FIELD_CP(MEM1, MEM1.actual)
     `RAL_FIELD_CP_16(MEM1, MEM1.actual, 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15)
  endgroup
  `endif

  // --------------------------
  // add constraint based on database legal values
  // --------------------------
  function void build();
    MEM2 = new("MEM2", "RO", 16, 0, {""});
    MEM2.set_rand_mode(0);
    void'(add_field( MEM2 ));

    MEM1 = new("MEM1", "RW", 16, 16, {""});
    MEM1.set_rand_mode(0);
    void'(add_field( MEM1 ));

  endfunction

endclass : mby_regs_MEM_reg

// ================================================

class ingress_regs_file extends sla_ral_file;

  rand mby_regs_DEVVENDID_reg DEVVENDID;
  rand mby_regs_BASE_ADDR_0_reg BASE_ADDR_0;
  rand mby_regs_MEM_reg MEM;

  `ovm_component_utils(ingress_regs_file)

  function new(string n, ovm_component p);
    super.new(n,p);
  endfunction

  // --------------------------
  function void build();
    `ifdef SLA_RAL_COVERAGE
    regfilename = this.get_name();
    `endif


    `ifdef SLA_RAL_COVERAGE
    sla_ral_reg::regname = "DEVVENDID";
    `endif
    DEVVENDID = mby_regs_DEVVENDID_reg::type_id::create("DEVVENDID", this);
    DEVVENDID.set_cfg(16'h00, 16'h0A, 16'h00, 4'h0, 32, 32'b00000000000000000000000000000000);
    DEVVENDID.set_space_addr("CFG", 4'h0);
    DEVVENDID.set_space_addr("MSG", 4'h0);
    DEVVENDID.set_space_addr("msg_bus_port", 'haa);
    DEVVENDID.set_space("CFG");
    if ( $test$plusargs("DEVVENDID:dont_test") ) DEVVENDID.set_test_reg(1'b0);
    if (!add_reg( DEVVENDID )) begin
      `slu_error(get_name(), ("Could not add register DEVVENDID"));
    end

    `ifdef SLA_RAL_COVERAGE
    sla_ral_reg::regname = "BASE_ADDR_0";
    `endif
    BASE_ADDR_0 = mby_regs_BASE_ADDR_0_reg::type_id::create("BASE_ADDR_0", this);
    BASE_ADDR_0.set_cfg(16'h00, 16'h0A, 16'h00, 8'h10, 32, 32'b00000000000000000000000000000000);
    BASE_ADDR_0.set_space_addr("CFG", 8'h10);
    BASE_ADDR_0.set_space_addr("MSG", 8'h10);
    BASE_ADDR_0.set_space_addr("msg_bus_port", 'haa);
    BASE_ADDR_0.set_space("CFG");
    if ( $test$plusargs("BASE_ADDR_0:dont_test") ) BASE_ADDR_0.set_test_reg(1'b0);
    if (!add_reg( BASE_ADDR_0 )) begin
      `slu_error(get_name(), ("Could not add register BASE_ADDR_0"));
    end

    `ifdef SLA_RAL_COVERAGE
    sla_ral_reg::regname = "MEM";
    `endif
    MEM = mby_regs_MEM_reg::type_id::create("MEM", this);
    MEM.set_cfg(16'h0, 16'h0, 16'h0, 4'h0, 32, 32'b00000000000000000000000000000000);
    MEM.set_space_addr("MSG", 4'h0);
    MEM.set_space_addr("msg_bus_port", 'haa);
    MEM.set_space_addr("MEM", 4'h0);
    MEM.set_space("MEM");
    if ( $test$plusargs("MEM:dont_test") ) MEM.set_test_reg(1'b0);
    if (!add_reg( MEM )) begin
      `slu_error(get_name(), ("Could not add register MEM"));
    end

    MEM.set_base_addr_reg(BASE_ADDR_0);
  endfunction

endclass : ingress_regs_file

// ================================================


`endif
