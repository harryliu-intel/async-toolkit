///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_trig_apply_map.sv                                  
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_trig_apply_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_RSTD


module rtlgen_mby_ppe_trig_apply_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_trig_apply_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_PH2_FF
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_TRIG_APPLY_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_trig_apply_map ( //lintra s-2096
    // Clocks


    // Resets



    // Register Inputs
    handcode_reg_rdata_TRIGGER_ACTION_CFG_1,
    handcode_reg_rdata_TRIGGER_ACTION_CFG_2,
    handcode_reg_rdata_TRIGGER_ACTION_GLORT,
    handcode_reg_rdata_TRIGGER_ACTION_MIRROR,
    handcode_reg_rdata_TRIGGER_CONDITION_AMASK_1,
    handcode_reg_rdata_TRIGGER_CONDITION_AMASK_2,
    handcode_reg_rdata_TRIGGER_CONDITION_CFG,
    handcode_reg_rdata_TRIGGER_CONDITION_CGRP,
    handcode_reg_rdata_TRIGGER_CONDITION_GLORT,
    handcode_reg_rdata_TRIGGER_CONDITION_PARAM,
    handcode_reg_rdata_TRIGGER_CONDITION_RX,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM0,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM1,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM2,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM3,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM4,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR0,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR1,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR2,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR3,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR4,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTRL,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX0,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX1,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX2,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX3,
    handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX4,
    handcode_reg_rdata_TRIGGER_STATS,

    handcode_rvalid_TRIGGER_ACTION_CFG_1,
    handcode_rvalid_TRIGGER_ACTION_CFG_2,
    handcode_rvalid_TRIGGER_ACTION_GLORT,
    handcode_rvalid_TRIGGER_ACTION_MIRROR,
    handcode_rvalid_TRIGGER_CONDITION_AMASK_1,
    handcode_rvalid_TRIGGER_CONDITION_AMASK_2,
    handcode_rvalid_TRIGGER_CONDITION_CFG,
    handcode_rvalid_TRIGGER_CONDITION_CGRP,
    handcode_rvalid_TRIGGER_CONDITION_GLORT,
    handcode_rvalid_TRIGGER_CONDITION_PARAM,
    handcode_rvalid_TRIGGER_CONDITION_RX,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM0,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM1,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM2,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM3,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADM4,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR0,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR1,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR2,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR3,
    handcode_rvalid_TRIGGER_DIRECT_MAP_ADR4,
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTRL,
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX0,
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX1,
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX2,
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX3,
    handcode_rvalid_TRIGGER_DIRECT_MAP_CTX4,
    handcode_rvalid_TRIGGER_STATS,

    handcode_wvalid_TRIGGER_ACTION_CFG_1,
    handcode_wvalid_TRIGGER_ACTION_CFG_2,
    handcode_wvalid_TRIGGER_ACTION_GLORT,
    handcode_wvalid_TRIGGER_ACTION_MIRROR,
    handcode_wvalid_TRIGGER_CONDITION_AMASK_1,
    handcode_wvalid_TRIGGER_CONDITION_AMASK_2,
    handcode_wvalid_TRIGGER_CONDITION_CFG,
    handcode_wvalid_TRIGGER_CONDITION_CGRP,
    handcode_wvalid_TRIGGER_CONDITION_GLORT,
    handcode_wvalid_TRIGGER_CONDITION_PARAM,
    handcode_wvalid_TRIGGER_CONDITION_RX,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM0,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM1,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM2,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM3,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADM4,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR0,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR1,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR2,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR3,
    handcode_wvalid_TRIGGER_DIRECT_MAP_ADR4,
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTRL,
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX0,
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX1,
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX2,
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX3,
    handcode_wvalid_TRIGGER_DIRECT_MAP_CTX4,
    handcode_wvalid_TRIGGER_STATS,

    handcode_error_TRIGGER_ACTION_CFG_1,
    handcode_error_TRIGGER_ACTION_CFG_2,
    handcode_error_TRIGGER_ACTION_GLORT,
    handcode_error_TRIGGER_ACTION_MIRROR,
    handcode_error_TRIGGER_CONDITION_AMASK_1,
    handcode_error_TRIGGER_CONDITION_AMASK_2,
    handcode_error_TRIGGER_CONDITION_CFG,
    handcode_error_TRIGGER_CONDITION_CGRP,
    handcode_error_TRIGGER_CONDITION_GLORT,
    handcode_error_TRIGGER_CONDITION_PARAM,
    handcode_error_TRIGGER_CONDITION_RX,
    handcode_error_TRIGGER_DIRECT_MAP_ADM0,
    handcode_error_TRIGGER_DIRECT_MAP_ADM1,
    handcode_error_TRIGGER_DIRECT_MAP_ADM2,
    handcode_error_TRIGGER_DIRECT_MAP_ADM3,
    handcode_error_TRIGGER_DIRECT_MAP_ADM4,
    handcode_error_TRIGGER_DIRECT_MAP_ADR0,
    handcode_error_TRIGGER_DIRECT_MAP_ADR1,
    handcode_error_TRIGGER_DIRECT_MAP_ADR2,
    handcode_error_TRIGGER_DIRECT_MAP_ADR3,
    handcode_error_TRIGGER_DIRECT_MAP_ADR4,
    handcode_error_TRIGGER_DIRECT_MAP_CTRL,
    handcode_error_TRIGGER_DIRECT_MAP_CTX0,
    handcode_error_TRIGGER_DIRECT_MAP_CTX1,
    handcode_error_TRIGGER_DIRECT_MAP_CTX2,
    handcode_error_TRIGGER_DIRECT_MAP_CTX3,
    handcode_error_TRIGGER_DIRECT_MAP_CTX4,
    handcode_error_TRIGGER_STATS,


    // Register Outputs

    // Register signals for HandCoded registers
    handcode_reg_wdata_TRIGGER_ACTION_CFG_1,
    handcode_reg_wdata_TRIGGER_ACTION_CFG_2,
    handcode_reg_wdata_TRIGGER_ACTION_GLORT,
    handcode_reg_wdata_TRIGGER_ACTION_MIRROR,
    handcode_reg_wdata_TRIGGER_CONDITION_AMASK_1,
    handcode_reg_wdata_TRIGGER_CONDITION_AMASK_2,
    handcode_reg_wdata_TRIGGER_CONDITION_CFG,
    handcode_reg_wdata_TRIGGER_CONDITION_CGRP,
    handcode_reg_wdata_TRIGGER_CONDITION_GLORT,
    handcode_reg_wdata_TRIGGER_CONDITION_PARAM,
    handcode_reg_wdata_TRIGGER_CONDITION_RX,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM0,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM1,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM2,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM3,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM4,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR0,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR1,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR2,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR3,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR4,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTRL,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX0,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX1,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX2,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX3,
    handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX4,
    handcode_reg_wdata_TRIGGER_STATS,

    we_TRIGGER_ACTION_CFG_1,
    we_TRIGGER_ACTION_CFG_2,
    we_TRIGGER_ACTION_GLORT,
    we_TRIGGER_ACTION_MIRROR,
    we_TRIGGER_CONDITION_AMASK_1,
    we_TRIGGER_CONDITION_AMASK_2,
    we_TRIGGER_CONDITION_CFG,
    we_TRIGGER_CONDITION_CGRP,
    we_TRIGGER_CONDITION_GLORT,
    we_TRIGGER_CONDITION_PARAM,
    we_TRIGGER_CONDITION_RX,
    we_TRIGGER_DIRECT_MAP_ADM0,
    we_TRIGGER_DIRECT_MAP_ADM1,
    we_TRIGGER_DIRECT_MAP_ADM2,
    we_TRIGGER_DIRECT_MAP_ADM3,
    we_TRIGGER_DIRECT_MAP_ADM4,
    we_TRIGGER_DIRECT_MAP_ADR0,
    we_TRIGGER_DIRECT_MAP_ADR1,
    we_TRIGGER_DIRECT_MAP_ADR2,
    we_TRIGGER_DIRECT_MAP_ADR3,
    we_TRIGGER_DIRECT_MAP_ADR4,
    we_TRIGGER_DIRECT_MAP_CTRL,
    we_TRIGGER_DIRECT_MAP_CTX0,
    we_TRIGGER_DIRECT_MAP_CTX1,
    we_TRIGGER_DIRECT_MAP_CTX2,
    we_TRIGGER_DIRECT_MAP_CTX3,
    we_TRIGGER_DIRECT_MAP_CTX4,
    we_TRIGGER_STATS,

    re_TRIGGER_ACTION_CFG_1,
    re_TRIGGER_ACTION_CFG_2,
    re_TRIGGER_ACTION_GLORT,
    re_TRIGGER_ACTION_MIRROR,
    re_TRIGGER_CONDITION_AMASK_1,
    re_TRIGGER_CONDITION_AMASK_2,
    re_TRIGGER_CONDITION_CFG,
    re_TRIGGER_CONDITION_CGRP,
    re_TRIGGER_CONDITION_GLORT,
    re_TRIGGER_CONDITION_PARAM,
    re_TRIGGER_CONDITION_RX,
    re_TRIGGER_DIRECT_MAP_ADM0,
    re_TRIGGER_DIRECT_MAP_ADM1,
    re_TRIGGER_DIRECT_MAP_ADM2,
    re_TRIGGER_DIRECT_MAP_ADM3,
    re_TRIGGER_DIRECT_MAP_ADM4,
    re_TRIGGER_DIRECT_MAP_ADR0,
    re_TRIGGER_DIRECT_MAP_ADR1,
    re_TRIGGER_DIRECT_MAP_ADR2,
    re_TRIGGER_DIRECT_MAP_ADR3,
    re_TRIGGER_DIRECT_MAP_ADR4,
    re_TRIGGER_DIRECT_MAP_CTRL,
    re_TRIGGER_DIRECT_MAP_CTX0,
    re_TRIGGER_DIRECT_MAP_CTX1,
    re_TRIGGER_DIRECT_MAP_CTX2,
    re_TRIGGER_DIRECT_MAP_CTX3,
    re_TRIGGER_DIRECT_MAP_CTX4,
    re_TRIGGER_STATS,




    // Config Access
    req,
    ack
    

);

import mby_ppe_trig_apply_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:0] MBY_PPE_TRIG_APPLY_MAP_OFFSET = {MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] TRIG_APPLY_SB_BAR = 3'b0;
parameter [7:0] TRIG_APPLY_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;

    // Clocks


    // Resets



    // Register Inputs
input TRIGGER_ACTION_CFG_1_t  handcode_reg_rdata_TRIGGER_ACTION_CFG_1;
input TRIGGER_ACTION_CFG_2_t  handcode_reg_rdata_TRIGGER_ACTION_CFG_2;
input TRIGGER_ACTION_GLORT_t  handcode_reg_rdata_TRIGGER_ACTION_GLORT;
input TRIGGER_ACTION_MIRROR_t  handcode_reg_rdata_TRIGGER_ACTION_MIRROR;
input TRIGGER_CONDITION_AMASK_1_t  handcode_reg_rdata_TRIGGER_CONDITION_AMASK_1;
input TRIGGER_CONDITION_AMASK_2_t  handcode_reg_rdata_TRIGGER_CONDITION_AMASK_2;
input TRIGGER_CONDITION_CFG_t  handcode_reg_rdata_TRIGGER_CONDITION_CFG;
input TRIGGER_CONDITION_CGRP_t  handcode_reg_rdata_TRIGGER_CONDITION_CGRP;
input TRIGGER_CONDITION_GLORT_t  handcode_reg_rdata_TRIGGER_CONDITION_GLORT;
input TRIGGER_CONDITION_PARAM_t  handcode_reg_rdata_TRIGGER_CONDITION_PARAM;
input TRIGGER_CONDITION_RX_t  handcode_reg_rdata_TRIGGER_CONDITION_RX;
input TRIGGER_DIRECT_MAP_ADM0_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM0;
input TRIGGER_DIRECT_MAP_ADM1_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM1;
input TRIGGER_DIRECT_MAP_ADM2_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM2;
input TRIGGER_DIRECT_MAP_ADM3_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM3;
input TRIGGER_DIRECT_MAP_ADM4_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM4;
input TRIGGER_DIRECT_MAP_ADR0_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR0;
input TRIGGER_DIRECT_MAP_ADR1_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR1;
input TRIGGER_DIRECT_MAP_ADR2_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR2;
input TRIGGER_DIRECT_MAP_ADR3_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR3;
input TRIGGER_DIRECT_MAP_ADR4_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR4;
input TRIGGER_DIRECT_MAP_CTRL_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTRL;
input TRIGGER_DIRECT_MAP_CTX0_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX0;
input TRIGGER_DIRECT_MAP_CTX1_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX1;
input TRIGGER_DIRECT_MAP_CTX2_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX2;
input TRIGGER_DIRECT_MAP_CTX3_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX3;
input TRIGGER_DIRECT_MAP_CTX4_t  handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX4;
input TRIGGER_STATS_t  handcode_reg_rdata_TRIGGER_STATS;

input handcode_rvalid_TRIGGER_ACTION_CFG_1_t  handcode_rvalid_TRIGGER_ACTION_CFG_1;
input handcode_rvalid_TRIGGER_ACTION_CFG_2_t  handcode_rvalid_TRIGGER_ACTION_CFG_2;
input handcode_rvalid_TRIGGER_ACTION_GLORT_t  handcode_rvalid_TRIGGER_ACTION_GLORT;
input handcode_rvalid_TRIGGER_ACTION_MIRROR_t  handcode_rvalid_TRIGGER_ACTION_MIRROR;
input handcode_rvalid_TRIGGER_CONDITION_AMASK_1_t  handcode_rvalid_TRIGGER_CONDITION_AMASK_1;
input handcode_rvalid_TRIGGER_CONDITION_AMASK_2_t  handcode_rvalid_TRIGGER_CONDITION_AMASK_2;
input handcode_rvalid_TRIGGER_CONDITION_CFG_t  handcode_rvalid_TRIGGER_CONDITION_CFG;
input handcode_rvalid_TRIGGER_CONDITION_CGRP_t  handcode_rvalid_TRIGGER_CONDITION_CGRP;
input handcode_rvalid_TRIGGER_CONDITION_GLORT_t  handcode_rvalid_TRIGGER_CONDITION_GLORT;
input handcode_rvalid_TRIGGER_CONDITION_PARAM_t  handcode_rvalid_TRIGGER_CONDITION_PARAM;
input handcode_rvalid_TRIGGER_CONDITION_RX_t  handcode_rvalid_TRIGGER_CONDITION_RX;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADM0_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADM0;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADM1_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADM1;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADM2_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADM2;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADM3_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADM3;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADM4_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADM4;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADR0_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADR0;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADR1_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADR1;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADR2_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADR2;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADR3_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADR3;
input handcode_rvalid_TRIGGER_DIRECT_MAP_ADR4_t  handcode_rvalid_TRIGGER_DIRECT_MAP_ADR4;
input handcode_rvalid_TRIGGER_DIRECT_MAP_CTRL_t  handcode_rvalid_TRIGGER_DIRECT_MAP_CTRL;
input handcode_rvalid_TRIGGER_DIRECT_MAP_CTX0_t  handcode_rvalid_TRIGGER_DIRECT_MAP_CTX0;
input handcode_rvalid_TRIGGER_DIRECT_MAP_CTX1_t  handcode_rvalid_TRIGGER_DIRECT_MAP_CTX1;
input handcode_rvalid_TRIGGER_DIRECT_MAP_CTX2_t  handcode_rvalid_TRIGGER_DIRECT_MAP_CTX2;
input handcode_rvalid_TRIGGER_DIRECT_MAP_CTX3_t  handcode_rvalid_TRIGGER_DIRECT_MAP_CTX3;
input handcode_rvalid_TRIGGER_DIRECT_MAP_CTX4_t  handcode_rvalid_TRIGGER_DIRECT_MAP_CTX4;
input handcode_rvalid_TRIGGER_STATS_t  handcode_rvalid_TRIGGER_STATS;

input handcode_wvalid_TRIGGER_ACTION_CFG_1_t  handcode_wvalid_TRIGGER_ACTION_CFG_1;
input handcode_wvalid_TRIGGER_ACTION_CFG_2_t  handcode_wvalid_TRIGGER_ACTION_CFG_2;
input handcode_wvalid_TRIGGER_ACTION_GLORT_t  handcode_wvalid_TRIGGER_ACTION_GLORT;
input handcode_wvalid_TRIGGER_ACTION_MIRROR_t  handcode_wvalid_TRIGGER_ACTION_MIRROR;
input handcode_wvalid_TRIGGER_CONDITION_AMASK_1_t  handcode_wvalid_TRIGGER_CONDITION_AMASK_1;
input handcode_wvalid_TRIGGER_CONDITION_AMASK_2_t  handcode_wvalid_TRIGGER_CONDITION_AMASK_2;
input handcode_wvalid_TRIGGER_CONDITION_CFG_t  handcode_wvalid_TRIGGER_CONDITION_CFG;
input handcode_wvalid_TRIGGER_CONDITION_CGRP_t  handcode_wvalid_TRIGGER_CONDITION_CGRP;
input handcode_wvalid_TRIGGER_CONDITION_GLORT_t  handcode_wvalid_TRIGGER_CONDITION_GLORT;
input handcode_wvalid_TRIGGER_CONDITION_PARAM_t  handcode_wvalid_TRIGGER_CONDITION_PARAM;
input handcode_wvalid_TRIGGER_CONDITION_RX_t  handcode_wvalid_TRIGGER_CONDITION_RX;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADM0_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADM0;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADM1_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADM1;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADM2_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADM2;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADM3_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADM3;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADM4_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADM4;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADR0_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADR0;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADR1_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADR1;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADR2_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADR2;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADR3_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADR3;
input handcode_wvalid_TRIGGER_DIRECT_MAP_ADR4_t  handcode_wvalid_TRIGGER_DIRECT_MAP_ADR4;
input handcode_wvalid_TRIGGER_DIRECT_MAP_CTRL_t  handcode_wvalid_TRIGGER_DIRECT_MAP_CTRL;
input handcode_wvalid_TRIGGER_DIRECT_MAP_CTX0_t  handcode_wvalid_TRIGGER_DIRECT_MAP_CTX0;
input handcode_wvalid_TRIGGER_DIRECT_MAP_CTX1_t  handcode_wvalid_TRIGGER_DIRECT_MAP_CTX1;
input handcode_wvalid_TRIGGER_DIRECT_MAP_CTX2_t  handcode_wvalid_TRIGGER_DIRECT_MAP_CTX2;
input handcode_wvalid_TRIGGER_DIRECT_MAP_CTX3_t  handcode_wvalid_TRIGGER_DIRECT_MAP_CTX3;
input handcode_wvalid_TRIGGER_DIRECT_MAP_CTX4_t  handcode_wvalid_TRIGGER_DIRECT_MAP_CTX4;
input handcode_wvalid_TRIGGER_STATS_t  handcode_wvalid_TRIGGER_STATS;

input handcode_error_TRIGGER_ACTION_CFG_1_t  handcode_error_TRIGGER_ACTION_CFG_1;
input handcode_error_TRIGGER_ACTION_CFG_2_t  handcode_error_TRIGGER_ACTION_CFG_2;
input handcode_error_TRIGGER_ACTION_GLORT_t  handcode_error_TRIGGER_ACTION_GLORT;
input handcode_error_TRIGGER_ACTION_MIRROR_t  handcode_error_TRIGGER_ACTION_MIRROR;
input handcode_error_TRIGGER_CONDITION_AMASK_1_t  handcode_error_TRIGGER_CONDITION_AMASK_1;
input handcode_error_TRIGGER_CONDITION_AMASK_2_t  handcode_error_TRIGGER_CONDITION_AMASK_2;
input handcode_error_TRIGGER_CONDITION_CFG_t  handcode_error_TRIGGER_CONDITION_CFG;
input handcode_error_TRIGGER_CONDITION_CGRP_t  handcode_error_TRIGGER_CONDITION_CGRP;
input handcode_error_TRIGGER_CONDITION_GLORT_t  handcode_error_TRIGGER_CONDITION_GLORT;
input handcode_error_TRIGGER_CONDITION_PARAM_t  handcode_error_TRIGGER_CONDITION_PARAM;
input handcode_error_TRIGGER_CONDITION_RX_t  handcode_error_TRIGGER_CONDITION_RX;
input handcode_error_TRIGGER_DIRECT_MAP_ADM0_t  handcode_error_TRIGGER_DIRECT_MAP_ADM0;
input handcode_error_TRIGGER_DIRECT_MAP_ADM1_t  handcode_error_TRIGGER_DIRECT_MAP_ADM1;
input handcode_error_TRIGGER_DIRECT_MAP_ADM2_t  handcode_error_TRIGGER_DIRECT_MAP_ADM2;
input handcode_error_TRIGGER_DIRECT_MAP_ADM3_t  handcode_error_TRIGGER_DIRECT_MAP_ADM3;
input handcode_error_TRIGGER_DIRECT_MAP_ADM4_t  handcode_error_TRIGGER_DIRECT_MAP_ADM4;
input handcode_error_TRIGGER_DIRECT_MAP_ADR0_t  handcode_error_TRIGGER_DIRECT_MAP_ADR0;
input handcode_error_TRIGGER_DIRECT_MAP_ADR1_t  handcode_error_TRIGGER_DIRECT_MAP_ADR1;
input handcode_error_TRIGGER_DIRECT_MAP_ADR2_t  handcode_error_TRIGGER_DIRECT_MAP_ADR2;
input handcode_error_TRIGGER_DIRECT_MAP_ADR3_t  handcode_error_TRIGGER_DIRECT_MAP_ADR3;
input handcode_error_TRIGGER_DIRECT_MAP_ADR4_t  handcode_error_TRIGGER_DIRECT_MAP_ADR4;
input handcode_error_TRIGGER_DIRECT_MAP_CTRL_t  handcode_error_TRIGGER_DIRECT_MAP_CTRL;
input handcode_error_TRIGGER_DIRECT_MAP_CTX0_t  handcode_error_TRIGGER_DIRECT_MAP_CTX0;
input handcode_error_TRIGGER_DIRECT_MAP_CTX1_t  handcode_error_TRIGGER_DIRECT_MAP_CTX1;
input handcode_error_TRIGGER_DIRECT_MAP_CTX2_t  handcode_error_TRIGGER_DIRECT_MAP_CTX2;
input handcode_error_TRIGGER_DIRECT_MAP_CTX3_t  handcode_error_TRIGGER_DIRECT_MAP_CTX3;
input handcode_error_TRIGGER_DIRECT_MAP_CTX4_t  handcode_error_TRIGGER_DIRECT_MAP_CTX4;
input handcode_error_TRIGGER_STATS_t  handcode_error_TRIGGER_STATS;


    // Register Outputs

    // Register signals for HandCoded registers
output TRIGGER_ACTION_CFG_1_t  handcode_reg_wdata_TRIGGER_ACTION_CFG_1;
output TRIGGER_ACTION_CFG_2_t  handcode_reg_wdata_TRIGGER_ACTION_CFG_2;
output TRIGGER_ACTION_GLORT_t  handcode_reg_wdata_TRIGGER_ACTION_GLORT;
output TRIGGER_ACTION_MIRROR_t  handcode_reg_wdata_TRIGGER_ACTION_MIRROR;
output TRIGGER_CONDITION_AMASK_1_t  handcode_reg_wdata_TRIGGER_CONDITION_AMASK_1;
output TRIGGER_CONDITION_AMASK_2_t  handcode_reg_wdata_TRIGGER_CONDITION_AMASK_2;
output TRIGGER_CONDITION_CFG_t  handcode_reg_wdata_TRIGGER_CONDITION_CFG;
output TRIGGER_CONDITION_CGRP_t  handcode_reg_wdata_TRIGGER_CONDITION_CGRP;
output TRIGGER_CONDITION_GLORT_t  handcode_reg_wdata_TRIGGER_CONDITION_GLORT;
output TRIGGER_CONDITION_PARAM_t  handcode_reg_wdata_TRIGGER_CONDITION_PARAM;
output TRIGGER_CONDITION_RX_t  handcode_reg_wdata_TRIGGER_CONDITION_RX;
output TRIGGER_DIRECT_MAP_ADM0_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM0;
output TRIGGER_DIRECT_MAP_ADM1_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM1;
output TRIGGER_DIRECT_MAP_ADM2_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM2;
output TRIGGER_DIRECT_MAP_ADM3_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM3;
output TRIGGER_DIRECT_MAP_ADM4_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM4;
output TRIGGER_DIRECT_MAP_ADR0_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR0;
output TRIGGER_DIRECT_MAP_ADR1_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR1;
output TRIGGER_DIRECT_MAP_ADR2_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR2;
output TRIGGER_DIRECT_MAP_ADR3_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR3;
output TRIGGER_DIRECT_MAP_ADR4_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR4;
output TRIGGER_DIRECT_MAP_CTRL_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTRL;
output TRIGGER_DIRECT_MAP_CTX0_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX0;
output TRIGGER_DIRECT_MAP_CTX1_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX1;
output TRIGGER_DIRECT_MAP_CTX2_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX2;
output TRIGGER_DIRECT_MAP_CTX3_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX3;
output TRIGGER_DIRECT_MAP_CTX4_t  handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX4;
output TRIGGER_STATS_t  handcode_reg_wdata_TRIGGER_STATS;

output we_TRIGGER_ACTION_CFG_1_t  we_TRIGGER_ACTION_CFG_1;
output we_TRIGGER_ACTION_CFG_2_t  we_TRIGGER_ACTION_CFG_2;
output we_TRIGGER_ACTION_GLORT_t  we_TRIGGER_ACTION_GLORT;
output we_TRIGGER_ACTION_MIRROR_t  we_TRIGGER_ACTION_MIRROR;
output we_TRIGGER_CONDITION_AMASK_1_t  we_TRIGGER_CONDITION_AMASK_1;
output we_TRIGGER_CONDITION_AMASK_2_t  we_TRIGGER_CONDITION_AMASK_2;
output we_TRIGGER_CONDITION_CFG_t  we_TRIGGER_CONDITION_CFG;
output we_TRIGGER_CONDITION_CGRP_t  we_TRIGGER_CONDITION_CGRP;
output we_TRIGGER_CONDITION_GLORT_t  we_TRIGGER_CONDITION_GLORT;
output we_TRIGGER_CONDITION_PARAM_t  we_TRIGGER_CONDITION_PARAM;
output we_TRIGGER_CONDITION_RX_t  we_TRIGGER_CONDITION_RX;
output we_TRIGGER_DIRECT_MAP_ADM0_t  we_TRIGGER_DIRECT_MAP_ADM0;
output we_TRIGGER_DIRECT_MAP_ADM1_t  we_TRIGGER_DIRECT_MAP_ADM1;
output we_TRIGGER_DIRECT_MAP_ADM2_t  we_TRIGGER_DIRECT_MAP_ADM2;
output we_TRIGGER_DIRECT_MAP_ADM3_t  we_TRIGGER_DIRECT_MAP_ADM3;
output we_TRIGGER_DIRECT_MAP_ADM4_t  we_TRIGGER_DIRECT_MAP_ADM4;
output we_TRIGGER_DIRECT_MAP_ADR0_t  we_TRIGGER_DIRECT_MAP_ADR0;
output we_TRIGGER_DIRECT_MAP_ADR1_t  we_TRIGGER_DIRECT_MAP_ADR1;
output we_TRIGGER_DIRECT_MAP_ADR2_t  we_TRIGGER_DIRECT_MAP_ADR2;
output we_TRIGGER_DIRECT_MAP_ADR3_t  we_TRIGGER_DIRECT_MAP_ADR3;
output we_TRIGGER_DIRECT_MAP_ADR4_t  we_TRIGGER_DIRECT_MAP_ADR4;
output we_TRIGGER_DIRECT_MAP_CTRL_t  we_TRIGGER_DIRECT_MAP_CTRL;
output we_TRIGGER_DIRECT_MAP_CTX0_t  we_TRIGGER_DIRECT_MAP_CTX0;
output we_TRIGGER_DIRECT_MAP_CTX1_t  we_TRIGGER_DIRECT_MAP_CTX1;
output we_TRIGGER_DIRECT_MAP_CTX2_t  we_TRIGGER_DIRECT_MAP_CTX2;
output we_TRIGGER_DIRECT_MAP_CTX3_t  we_TRIGGER_DIRECT_MAP_CTX3;
output we_TRIGGER_DIRECT_MAP_CTX4_t  we_TRIGGER_DIRECT_MAP_CTX4;
output we_TRIGGER_STATS_t  we_TRIGGER_STATS;

output re_TRIGGER_ACTION_CFG_1_t  re_TRIGGER_ACTION_CFG_1;
output re_TRIGGER_ACTION_CFG_2_t  re_TRIGGER_ACTION_CFG_2;
output re_TRIGGER_ACTION_GLORT_t  re_TRIGGER_ACTION_GLORT;
output re_TRIGGER_ACTION_MIRROR_t  re_TRIGGER_ACTION_MIRROR;
output re_TRIGGER_CONDITION_AMASK_1_t  re_TRIGGER_CONDITION_AMASK_1;
output re_TRIGGER_CONDITION_AMASK_2_t  re_TRIGGER_CONDITION_AMASK_2;
output re_TRIGGER_CONDITION_CFG_t  re_TRIGGER_CONDITION_CFG;
output re_TRIGGER_CONDITION_CGRP_t  re_TRIGGER_CONDITION_CGRP;
output re_TRIGGER_CONDITION_GLORT_t  re_TRIGGER_CONDITION_GLORT;
output re_TRIGGER_CONDITION_PARAM_t  re_TRIGGER_CONDITION_PARAM;
output re_TRIGGER_CONDITION_RX_t  re_TRIGGER_CONDITION_RX;
output re_TRIGGER_DIRECT_MAP_ADM0_t  re_TRIGGER_DIRECT_MAP_ADM0;
output re_TRIGGER_DIRECT_MAP_ADM1_t  re_TRIGGER_DIRECT_MAP_ADM1;
output re_TRIGGER_DIRECT_MAP_ADM2_t  re_TRIGGER_DIRECT_MAP_ADM2;
output re_TRIGGER_DIRECT_MAP_ADM3_t  re_TRIGGER_DIRECT_MAP_ADM3;
output re_TRIGGER_DIRECT_MAP_ADM4_t  re_TRIGGER_DIRECT_MAP_ADM4;
output re_TRIGGER_DIRECT_MAP_ADR0_t  re_TRIGGER_DIRECT_MAP_ADR0;
output re_TRIGGER_DIRECT_MAP_ADR1_t  re_TRIGGER_DIRECT_MAP_ADR1;
output re_TRIGGER_DIRECT_MAP_ADR2_t  re_TRIGGER_DIRECT_MAP_ADR2;
output re_TRIGGER_DIRECT_MAP_ADR3_t  re_TRIGGER_DIRECT_MAP_ADR3;
output re_TRIGGER_DIRECT_MAP_ADR4_t  re_TRIGGER_DIRECT_MAP_ADR4;
output re_TRIGGER_DIRECT_MAP_CTRL_t  re_TRIGGER_DIRECT_MAP_CTRL;
output re_TRIGGER_DIRECT_MAP_CTX0_t  re_TRIGGER_DIRECT_MAP_CTX0;
output re_TRIGGER_DIRECT_MAP_CTX1_t  re_TRIGGER_DIRECT_MAP_CTX1;
output re_TRIGGER_DIRECT_MAP_CTX2_t  re_TRIGGER_DIRECT_MAP_CTX2;
output re_TRIGGER_DIRECT_MAP_CTX3_t  re_TRIGGER_DIRECT_MAP_CTX3;
output re_TRIGGER_DIRECT_MAP_CTX4_t  re_TRIGGER_DIRECT_MAP_CTX4;
output re_TRIGGER_STATS_t  re_TRIGGER_STATS;




    // Config Access
input mby_ppe_trig_apply_map_cr_req_t  req;
output mby_ppe_trig_apply_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_trig_apply_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_TRIG_APPLY_MAP_MEM;
assign case_req_addr_MBY_PPE_TRIG_APPLY_MAP_MEM = req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_trig_apply;
always_comb begin : sb_fid_cond_trig_apply_BLOCK
    unique casez (req_fid) 
		TRIG_APPLY_SB_FID: sb_fid_cond_trig_apply = 1;
		default: sb_fid_cond_trig_apply = 0;
    endcase 
end


logic sb_bar_cond_trig_apply;
always_comb begin : sb_bar_cond_trig_apply_BLOCK
    unique casez (req_bar) 
		TRIG_APPLY_SB_BAR: sb_bar_cond_trig_apply = 1;
		default: sb_bar_cond_trig_apply = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// TRIGGER_CONDITION_CFG using HANDCODED_REG template.
logic addr_decode_TRIGGER_CONDITION_CFG;
logic write_req_TRIGGER_CONDITION_CFG;
logic read_req_TRIGGER_CONDITION_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b0?,4'h?,1'b?},
      {44'h2?,1'b?}:
          addr_decode_TRIGGER_CONDITION_CFG = req.valid;
      default: 
         addr_decode_TRIGGER_CONDITION_CFG = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_CONDITION_CFG = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_CONDITION_CFG ;
always_comb read_req_TRIGGER_CONDITION_CFG  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_CONDITION_CFG ;

always_comb we_TRIGGER_CONDITION_CFG = {8{write_req_TRIGGER_CONDITION_CFG}} & be;
always_comb re_TRIGGER_CONDITION_CFG = {8{read_req_TRIGGER_CONDITION_CFG}} & be;
always_comb handcode_reg_wdata_TRIGGER_CONDITION_CFG = write_data;


// ----------------------------------------------------------------------
// TRIGGER_CONDITION_PARAM using HANDCODED_REG template.
logic addr_decode_TRIGGER_CONDITION_PARAM;
logic write_req_TRIGGER_CONDITION_PARAM;
logic read_req_TRIGGER_CONDITION_PARAM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h3?,1'b?},
      {40'b10?,4'h?,1'b?}:
          addr_decode_TRIGGER_CONDITION_PARAM = req.valid;
      default: 
         addr_decode_TRIGGER_CONDITION_PARAM = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_CONDITION_PARAM = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_CONDITION_PARAM ;
always_comb read_req_TRIGGER_CONDITION_PARAM  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_CONDITION_PARAM ;

always_comb we_TRIGGER_CONDITION_PARAM = {8{write_req_TRIGGER_CONDITION_PARAM}} & be;
always_comb re_TRIGGER_CONDITION_PARAM = {8{read_req_TRIGGER_CONDITION_PARAM}} & be;
always_comb handcode_reg_wdata_TRIGGER_CONDITION_PARAM = write_data;


// ----------------------------------------------------------------------
// TRIGGER_CONDITION_CGRP using HANDCODED_REG template.
logic addr_decode_TRIGGER_CONDITION_CGRP;
logic write_req_TRIGGER_CONDITION_CGRP;
logic read_req_TRIGGER_CONDITION_CGRP;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b11?,4'h?,1'b?},
      {44'h8?,1'b?}:
          addr_decode_TRIGGER_CONDITION_CGRP = req.valid;
      default: 
         addr_decode_TRIGGER_CONDITION_CGRP = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_CONDITION_CGRP = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_CONDITION_CGRP ;
always_comb read_req_TRIGGER_CONDITION_CGRP  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_CONDITION_CGRP ;

always_comb we_TRIGGER_CONDITION_CGRP = {8{write_req_TRIGGER_CONDITION_CGRP}} & be;
always_comb re_TRIGGER_CONDITION_CGRP = {8{read_req_TRIGGER_CONDITION_CGRP}} & be;
always_comb handcode_reg_wdata_TRIGGER_CONDITION_CGRP = write_data;


// ----------------------------------------------------------------------
// TRIGGER_CONDITION_GLORT using HANDCODED_REG template.
logic addr_decode_TRIGGER_CONDITION_GLORT;
logic write_req_TRIGGER_CONDITION_GLORT;
logic read_req_TRIGGER_CONDITION_GLORT;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h9?,1'b?},
      {40'b101?,4'h?,1'b?}:
          addr_decode_TRIGGER_CONDITION_GLORT = req.valid;
      default: 
         addr_decode_TRIGGER_CONDITION_GLORT = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_CONDITION_GLORT = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_CONDITION_GLORT ;
always_comb read_req_TRIGGER_CONDITION_GLORT  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_CONDITION_GLORT ;

always_comb we_TRIGGER_CONDITION_GLORT = {8{write_req_TRIGGER_CONDITION_GLORT}} & be;
always_comb re_TRIGGER_CONDITION_GLORT = {8{read_req_TRIGGER_CONDITION_GLORT}} & be;
always_comb handcode_reg_wdata_TRIGGER_CONDITION_GLORT = write_data;


// ----------------------------------------------------------------------
// TRIGGER_CONDITION_RX using HANDCODED_REG template.
logic addr_decode_TRIGGER_CONDITION_RX;
logic write_req_TRIGGER_CONDITION_RX;
logic read_req_TRIGGER_CONDITION_RX;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'b110?,4'h?,1'b?},
      {44'hE?,1'b?}:
          addr_decode_TRIGGER_CONDITION_RX = req.valid;
      default: 
         addr_decode_TRIGGER_CONDITION_RX = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_CONDITION_RX = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_CONDITION_RX ;
always_comb read_req_TRIGGER_CONDITION_RX  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_CONDITION_RX ;

always_comb we_TRIGGER_CONDITION_RX = {8{write_req_TRIGGER_CONDITION_RX}} & be;
always_comb re_TRIGGER_CONDITION_RX = {8{read_req_TRIGGER_CONDITION_RX}} & be;
always_comb handcode_reg_wdata_TRIGGER_CONDITION_RX = write_data;


// ----------------------------------------------------------------------
// TRIGGER_CONDITION_AMASK_1 using HANDCODED_REG template.
logic addr_decode_TRIGGER_CONDITION_AMASK_1;
logic write_req_TRIGGER_CONDITION_AMASK_1;
logic read_req_TRIGGER_CONDITION_AMASK_1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'hF?,1'b?},
      {36'h1,4'b000?,4'h?,1'b?}:
          addr_decode_TRIGGER_CONDITION_AMASK_1 = req.valid;
      default: 
         addr_decode_TRIGGER_CONDITION_AMASK_1 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_CONDITION_AMASK_1 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_CONDITION_AMASK_1 ;
always_comb read_req_TRIGGER_CONDITION_AMASK_1  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_CONDITION_AMASK_1 ;

always_comb we_TRIGGER_CONDITION_AMASK_1 = {8{write_req_TRIGGER_CONDITION_AMASK_1}} & be;
always_comb re_TRIGGER_CONDITION_AMASK_1 = {8{read_req_TRIGGER_CONDITION_AMASK_1}} & be;
always_comb handcode_reg_wdata_TRIGGER_CONDITION_AMASK_1 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_CONDITION_AMASK_2 using HANDCODED_REG template.
logic addr_decode_TRIGGER_CONDITION_AMASK_2;
logic write_req_TRIGGER_CONDITION_AMASK_2;
logic read_req_TRIGGER_CONDITION_AMASK_2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h1,4'b001?,4'h?,1'b?},
      {44'h14?,1'b?}:
          addr_decode_TRIGGER_CONDITION_AMASK_2 = req.valid;
      default: 
         addr_decode_TRIGGER_CONDITION_AMASK_2 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_CONDITION_AMASK_2 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_CONDITION_AMASK_2 ;
always_comb read_req_TRIGGER_CONDITION_AMASK_2  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_CONDITION_AMASK_2 ;

always_comb we_TRIGGER_CONDITION_AMASK_2 = {8{write_req_TRIGGER_CONDITION_AMASK_2}} & be;
always_comb re_TRIGGER_CONDITION_AMASK_2 = {8{read_req_TRIGGER_CONDITION_AMASK_2}} & be;
always_comb handcode_reg_wdata_TRIGGER_CONDITION_AMASK_2 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_ACTION_CFG_1 using HANDCODED_REG template.
logic addr_decode_TRIGGER_ACTION_CFG_1;
logic write_req_TRIGGER_ACTION_CFG_1;
logic read_req_TRIGGER_ACTION_CFG_1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h15?,1'b?},
      {36'h1,4'b011?,4'h?,1'b?}:
          addr_decode_TRIGGER_ACTION_CFG_1 = req.valid;
      default: 
         addr_decode_TRIGGER_ACTION_CFG_1 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_ACTION_CFG_1 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_ACTION_CFG_1 ;
always_comb read_req_TRIGGER_ACTION_CFG_1  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_ACTION_CFG_1 ;

always_comb we_TRIGGER_ACTION_CFG_1 = {8{write_req_TRIGGER_ACTION_CFG_1}} & be;
always_comb re_TRIGGER_ACTION_CFG_1 = {8{read_req_TRIGGER_ACTION_CFG_1}} & be;
always_comb handcode_reg_wdata_TRIGGER_ACTION_CFG_1 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_ACTION_CFG_2 using HANDCODED_REG template.
logic addr_decode_TRIGGER_ACTION_CFG_2;
logic write_req_TRIGGER_ACTION_CFG_2;
logic read_req_TRIGGER_ACTION_CFG_2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h1,4'b100?,4'h?,1'b?},
      {44'h1A?,1'b?}:
          addr_decode_TRIGGER_ACTION_CFG_2 = req.valid;
      default: 
         addr_decode_TRIGGER_ACTION_CFG_2 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_ACTION_CFG_2 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_ACTION_CFG_2 ;
always_comb read_req_TRIGGER_ACTION_CFG_2  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_ACTION_CFG_2 ;

always_comb we_TRIGGER_ACTION_CFG_2 = {8{write_req_TRIGGER_ACTION_CFG_2}} & be;
always_comb re_TRIGGER_ACTION_CFG_2 = {8{read_req_TRIGGER_ACTION_CFG_2}} & be;
always_comb handcode_reg_wdata_TRIGGER_ACTION_CFG_2 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_ACTION_GLORT using HANDCODED_REG template.
logic addr_decode_TRIGGER_ACTION_GLORT;
logic write_req_TRIGGER_ACTION_GLORT;
logic read_req_TRIGGER_ACTION_GLORT;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h1B?,1'b?},
      {36'h1,4'b110?,4'h?,1'b?}:
          addr_decode_TRIGGER_ACTION_GLORT = req.valid;
      default: 
         addr_decode_TRIGGER_ACTION_GLORT = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_ACTION_GLORT = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_ACTION_GLORT ;
always_comb read_req_TRIGGER_ACTION_GLORT  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_ACTION_GLORT ;

always_comb we_TRIGGER_ACTION_GLORT = {8{write_req_TRIGGER_ACTION_GLORT}} & be;
always_comb re_TRIGGER_ACTION_GLORT = {8{read_req_TRIGGER_ACTION_GLORT}} & be;
always_comb handcode_reg_wdata_TRIGGER_ACTION_GLORT = write_data;


// ----------------------------------------------------------------------
// TRIGGER_ACTION_MIRROR using HANDCODED_REG template.
logic addr_decode_TRIGGER_ACTION_MIRROR;
logic write_req_TRIGGER_ACTION_MIRROR;
logic read_req_TRIGGER_ACTION_MIRROR;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h1,4'b111?,4'h?,1'b?},
      {44'h20?,1'b?}:
          addr_decode_TRIGGER_ACTION_MIRROR = req.valid;
      default: 
         addr_decode_TRIGGER_ACTION_MIRROR = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_ACTION_MIRROR = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_ACTION_MIRROR ;
always_comb read_req_TRIGGER_ACTION_MIRROR  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_ACTION_MIRROR ;

always_comb we_TRIGGER_ACTION_MIRROR = {8{write_req_TRIGGER_ACTION_MIRROR}} & be;
always_comb re_TRIGGER_ACTION_MIRROR = {8{read_req_TRIGGER_ACTION_MIRROR}} & be;
always_comb handcode_reg_wdata_TRIGGER_ACTION_MIRROR = write_data;


// ----------------------------------------------------------------------
// TRIGGER_STATS using HANDCODED_REG template.
logic addr_decode_TRIGGER_STATS;
logic write_req_TRIGGER_STATS;
logic read_req_TRIGGER_STATS;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h21?,1'b?},
      {36'h2,4'b001?,4'h?,1'b?}:
          addr_decode_TRIGGER_STATS = req.valid;
      default: 
         addr_decode_TRIGGER_STATS = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_STATS = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_STATS ;
always_comb read_req_TRIGGER_STATS  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_STATS ;

always_comb we_TRIGGER_STATS = {8{write_req_TRIGGER_STATS}} & be;
always_comb re_TRIGGER_STATS = {8{read_req_TRIGGER_STATS}} & be;
always_comb handcode_reg_wdata_TRIGGER_STATS = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_CTRL using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_CTRL;
logic write_req_TRIGGER_DIRECT_MAP_CTRL;
logic read_req_TRIGGER_DIRECT_MAP_CTRL;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h240,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_CTRL = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_CTRL = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_CTRL = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTRL ;
always_comb read_req_TRIGGER_DIRECT_MAP_CTRL  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTRL ;

always_comb we_TRIGGER_DIRECT_MAP_CTRL = {8{write_req_TRIGGER_DIRECT_MAP_CTRL}} & be;
always_comb re_TRIGGER_DIRECT_MAP_CTRL = {8{read_req_TRIGGER_DIRECT_MAP_CTRL}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTRL = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_CTX0 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_CTX0;
logic write_req_TRIGGER_DIRECT_MAP_CTX0;
logic read_req_TRIGGER_DIRECT_MAP_CTX0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h240,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX0 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX0 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_CTX0 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX0 ;
always_comb read_req_TRIGGER_DIRECT_MAP_CTX0  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX0 ;

always_comb we_TRIGGER_DIRECT_MAP_CTX0 = {8{write_req_TRIGGER_DIRECT_MAP_CTX0}} & be;
always_comb re_TRIGGER_DIRECT_MAP_CTX0 = {8{read_req_TRIGGER_DIRECT_MAP_CTX0}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX0 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_CTX1 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_CTX1;
logic write_req_TRIGGER_DIRECT_MAP_CTX1;
logic read_req_TRIGGER_DIRECT_MAP_CTX1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h241,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX1 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX1 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_CTX1 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX1 ;
always_comb read_req_TRIGGER_DIRECT_MAP_CTX1  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX1 ;

always_comb we_TRIGGER_DIRECT_MAP_CTX1 = {8{write_req_TRIGGER_DIRECT_MAP_CTX1}} & be;
always_comb re_TRIGGER_DIRECT_MAP_CTX1 = {8{read_req_TRIGGER_DIRECT_MAP_CTX1}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX1 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_CTX2 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_CTX2;
logic write_req_TRIGGER_DIRECT_MAP_CTX2;
logic read_req_TRIGGER_DIRECT_MAP_CTX2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h241,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX2 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX2 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_CTX2 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX2 ;
always_comb read_req_TRIGGER_DIRECT_MAP_CTX2  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX2 ;

always_comb we_TRIGGER_DIRECT_MAP_CTX2 = {8{write_req_TRIGGER_DIRECT_MAP_CTX2}} & be;
always_comb re_TRIGGER_DIRECT_MAP_CTX2 = {8{read_req_TRIGGER_DIRECT_MAP_CTX2}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX2 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_CTX3 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_CTX3;
logic write_req_TRIGGER_DIRECT_MAP_CTX3;
logic read_req_TRIGGER_DIRECT_MAP_CTX3;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h242,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX3 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX3 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_CTX3 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX3 ;
always_comb read_req_TRIGGER_DIRECT_MAP_CTX3  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX3 ;

always_comb we_TRIGGER_DIRECT_MAP_CTX3 = {8{write_req_TRIGGER_DIRECT_MAP_CTX3}} & be;
always_comb re_TRIGGER_DIRECT_MAP_CTX3 = {8{read_req_TRIGGER_DIRECT_MAP_CTX3}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX3 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_CTX4 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_CTX4;
logic write_req_TRIGGER_DIRECT_MAP_CTX4;
logic read_req_TRIGGER_DIRECT_MAP_CTX4;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h242,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX4 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_CTX4 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_CTX4 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX4 ;
always_comb read_req_TRIGGER_DIRECT_MAP_CTX4  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_CTX4 ;

always_comb we_TRIGGER_DIRECT_MAP_CTX4 = {8{write_req_TRIGGER_DIRECT_MAP_CTX4}} & be;
always_comb re_TRIGGER_DIRECT_MAP_CTX4 = {8{read_req_TRIGGER_DIRECT_MAP_CTX4}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_CTX4 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADM0 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADM0;
logic write_req_TRIGGER_DIRECT_MAP_ADM0;
logic read_req_TRIGGER_DIRECT_MAP_ADM0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h243,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM0 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM0 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADM0 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM0 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADM0  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM0 ;

always_comb we_TRIGGER_DIRECT_MAP_ADM0 = {8{write_req_TRIGGER_DIRECT_MAP_ADM0}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADM0 = {8{read_req_TRIGGER_DIRECT_MAP_ADM0}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM0 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADM1 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADM1;
logic write_req_TRIGGER_DIRECT_MAP_ADM1;
logic read_req_TRIGGER_DIRECT_MAP_ADM1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h243,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM1 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM1 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADM1 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM1 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADM1  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM1 ;

always_comb we_TRIGGER_DIRECT_MAP_ADM1 = {8{write_req_TRIGGER_DIRECT_MAP_ADM1}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADM1 = {8{read_req_TRIGGER_DIRECT_MAP_ADM1}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM1 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADM2 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADM2;
logic write_req_TRIGGER_DIRECT_MAP_ADM2;
logic read_req_TRIGGER_DIRECT_MAP_ADM2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h244,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM2 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM2 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADM2 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM2 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADM2  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM2 ;

always_comb we_TRIGGER_DIRECT_MAP_ADM2 = {8{write_req_TRIGGER_DIRECT_MAP_ADM2}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADM2 = {8{read_req_TRIGGER_DIRECT_MAP_ADM2}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM2 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADM3 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADM3;
logic write_req_TRIGGER_DIRECT_MAP_ADM3;
logic read_req_TRIGGER_DIRECT_MAP_ADM3;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h244,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM3 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM3 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADM3 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM3 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADM3  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM3 ;

always_comb we_TRIGGER_DIRECT_MAP_ADM3 = {8{write_req_TRIGGER_DIRECT_MAP_ADM3}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADM3 = {8{read_req_TRIGGER_DIRECT_MAP_ADM3}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM3 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADM4 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADM4;
logic write_req_TRIGGER_DIRECT_MAP_ADM4;
logic read_req_TRIGGER_DIRECT_MAP_ADM4;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h245,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM4 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADM4 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADM4 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM4 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADM4  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADM4 ;

always_comb we_TRIGGER_DIRECT_MAP_ADM4 = {8{write_req_TRIGGER_DIRECT_MAP_ADM4}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADM4 = {8{read_req_TRIGGER_DIRECT_MAP_ADM4}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADM4 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADR0 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADR0;
logic write_req_TRIGGER_DIRECT_MAP_ADR0;
logic read_req_TRIGGER_DIRECT_MAP_ADR0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h245,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR0 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR0 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADR0 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR0 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADR0  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR0 ;

always_comb we_TRIGGER_DIRECT_MAP_ADR0 = {8{write_req_TRIGGER_DIRECT_MAP_ADR0}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADR0 = {8{read_req_TRIGGER_DIRECT_MAP_ADR0}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR0 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADR1 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADR1;
logic write_req_TRIGGER_DIRECT_MAP_ADR1;
logic read_req_TRIGGER_DIRECT_MAP_ADR1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h246,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR1 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR1 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADR1 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR1 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADR1  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR1 ;

always_comb we_TRIGGER_DIRECT_MAP_ADR1 = {8{write_req_TRIGGER_DIRECT_MAP_ADR1}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADR1 = {8{read_req_TRIGGER_DIRECT_MAP_ADR1}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR1 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADR2 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADR2;
logic write_req_TRIGGER_DIRECT_MAP_ADR2;
logic read_req_TRIGGER_DIRECT_MAP_ADR2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h246,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR2 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR2 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADR2 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR2 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADR2  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR2 ;

always_comb we_TRIGGER_DIRECT_MAP_ADR2 = {8{write_req_TRIGGER_DIRECT_MAP_ADR2}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADR2 = {8{read_req_TRIGGER_DIRECT_MAP_ADR2}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR2 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADR3 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADR3;
logic write_req_TRIGGER_DIRECT_MAP_ADR3;
logic read_req_TRIGGER_DIRECT_MAP_ADR3;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h247,1'b0}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR3 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR3 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADR3 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR3 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADR3  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR3 ;

always_comb we_TRIGGER_DIRECT_MAP_ADR3 = {8{write_req_TRIGGER_DIRECT_MAP_ADR3}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADR3 = {8{read_req_TRIGGER_DIRECT_MAP_ADR3}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR3 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_DIRECT_MAP_ADR4 using HANDCODED_REG template.
logic addr_decode_TRIGGER_DIRECT_MAP_ADR4;
logic write_req_TRIGGER_DIRECT_MAP_ADR4;
logic read_req_TRIGGER_DIRECT_MAP_ADR4;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h247,1'b1}: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR4 = req.valid;
      default: 
         addr_decode_TRIGGER_DIRECT_MAP_ADR4 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_DIRECT_MAP_ADR4 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR4 ;
always_comb read_req_TRIGGER_DIRECT_MAP_ADR4  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_DIRECT_MAP_ADR4 ;

always_comb we_TRIGGER_DIRECT_MAP_ADR4 = {8{write_req_TRIGGER_DIRECT_MAP_ADR4}} & be;
always_comb re_TRIGGER_DIRECT_MAP_ADR4 = {8{read_req_TRIGGER_DIRECT_MAP_ADR4}} & be;
always_comb handcode_reg_wdata_TRIGGER_DIRECT_MAP_ADR4 = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_TRIG_APPLY_MAP_MEM) 
           {40'b0?,4'h?,1'b?},
           {44'h2?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_CONDITION_CFG;
                    ack.read_miss = handcode_error_TRIGGER_CONDITION_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h3?,1'b?},
           {40'b10?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_CONDITION_PARAM;
                    ack.read_miss = handcode_error_TRIGGER_CONDITION_PARAM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'b11?,4'h?,1'b?},
           {44'h8?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_CONDITION_CGRP;
                    ack.read_miss = handcode_error_TRIGGER_CONDITION_CGRP;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h9?,1'b?},
           {40'b101?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_CONDITION_GLORT;
                    ack.read_miss = handcode_error_TRIGGER_CONDITION_GLORT;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'b110?,4'h?,1'b?},
           {44'hE?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_CONDITION_RX;
                    ack.read_miss = handcode_error_TRIGGER_CONDITION_RX;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'hF?,1'b?},
           {36'h1,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_CONDITION_AMASK_1;
                    ack.read_miss = handcode_error_TRIGGER_CONDITION_AMASK_1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h1,4'b001?,4'h?,1'b?},
           {44'h14?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_CONDITION_AMASK_2;
                    ack.read_miss = handcode_error_TRIGGER_CONDITION_AMASK_2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h15?,1'b?},
           {36'h1,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_ACTION_CFG_1;
                    ack.read_miss = handcode_error_TRIGGER_ACTION_CFG_1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h1,4'b100?,4'h?,1'b?},
           {44'h1A?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_ACTION_CFG_2;
                    ack.read_miss = handcode_error_TRIGGER_ACTION_CFG_2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h1B?,1'b?},
           {36'h1,4'b110?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_ACTION_GLORT;
                    ack.read_miss = handcode_error_TRIGGER_ACTION_GLORT;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h1,4'b111?,4'h?,1'b?},
           {44'h20?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_ACTION_MIRROR;
                    ack.read_miss = handcode_error_TRIGGER_ACTION_MIRROR;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h21?,1'b?},
           {36'h2,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_STATS;
                    ack.read_miss = handcode_error_TRIGGER_STATS;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h240,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_CTRL;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_CTRL;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h240,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_CTX0;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h241,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_CTX1;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h241,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_CTX2;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h242,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_CTX3;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX3;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h242,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_CTX4;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX4;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h243,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADM0;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h243,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADM1;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h244,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADM2;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h244,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADM3;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM3;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h245,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADM4;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM4;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h245,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADR0;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h246,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADR1;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h246,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADR2;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h247,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADR3;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR3;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h247,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_DIRECT_MAP_ADR4;
                    ack.read_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR4;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_TRIG_APPLY_MAP_MEM) 
           {40'b0?,4'h?,1'b?},
           {44'h2?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_CONDITION_CFG;
                    ack.write_miss = handcode_error_TRIGGER_CONDITION_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h3?,1'b?},
           {40'b10?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_CONDITION_PARAM;
                    ack.write_miss = handcode_error_TRIGGER_CONDITION_PARAM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'b11?,4'h?,1'b?},
           {44'h8?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_CONDITION_CGRP;
                    ack.write_miss = handcode_error_TRIGGER_CONDITION_CGRP;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h9?,1'b?},
           {40'b101?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_CONDITION_GLORT;
                    ack.write_miss = handcode_error_TRIGGER_CONDITION_GLORT;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'b110?,4'h?,1'b?},
           {44'hE?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_CONDITION_RX;
                    ack.write_miss = handcode_error_TRIGGER_CONDITION_RX;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'hF?,1'b?},
           {36'h1,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_CONDITION_AMASK_1;
                    ack.write_miss = handcode_error_TRIGGER_CONDITION_AMASK_1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h1,4'b001?,4'h?,1'b?},
           {44'h14?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_CONDITION_AMASK_2;
                    ack.write_miss = handcode_error_TRIGGER_CONDITION_AMASK_2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h15?,1'b?},
           {36'h1,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_ACTION_CFG_1;
                    ack.write_miss = handcode_error_TRIGGER_ACTION_CFG_1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h1,4'b100?,4'h?,1'b?},
           {44'h1A?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_ACTION_CFG_2;
                    ack.write_miss = handcode_error_TRIGGER_ACTION_CFG_2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h1B?,1'b?},
           {36'h1,4'b110?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_ACTION_GLORT;
                    ack.write_miss = handcode_error_TRIGGER_ACTION_GLORT;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h1,4'b111?,4'h?,1'b?},
           {44'h20?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_ACTION_MIRROR;
                    ack.write_miss = handcode_error_TRIGGER_ACTION_MIRROR;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h21?,1'b?},
           {36'h2,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_STATS;
                    ack.write_miss = handcode_error_TRIGGER_STATS;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h240,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_CTRL;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_CTRL;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h240,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_CTX0;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h241,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_CTX1;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h241,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_CTX2;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h242,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_CTX3;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX3;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h242,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_CTX4;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_CTX4;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h243,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADM0;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h243,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADM1;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h244,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADM2;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h244,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADM3;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM3;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h245,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADM4;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADM4;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h245,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADR0;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h246,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADR1;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h246,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADR2;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h247,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADR3;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR3;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h247,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_DIRECT_MAP_ADR4;
                    ack.write_miss = handcode_error_TRIGGER_DIRECT_MAP_ADR4;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_TRIG_APPLY_MAP_MEM) 
           {40'b0?,4'h?,1'b?},
           {44'h2?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_CONDITION_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'h3?,1'b?},
           {40'b10?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_CONDITION_PARAM;
                 default: read_data = '0;
              endcase
           end
           {40'b11?,4'h?,1'b?},
           {44'h8?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_CONDITION_CGRP;
                 default: read_data = '0;
              endcase
           end
           {44'h9?,1'b?},
           {40'b101?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_CONDITION_GLORT;
                 default: read_data = '0;
              endcase
           end
           {40'b110?,4'h?,1'b?},
           {44'hE?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_CONDITION_RX;
                 default: read_data = '0;
              endcase
           end
           {44'hF?,1'b?},
           {36'h1,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_CONDITION_AMASK_1;
                 default: read_data = '0;
              endcase
           end
           {36'h1,4'b001?,4'h?,1'b?},
           {44'h14?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_CONDITION_AMASK_2;
                 default: read_data = '0;
              endcase
           end
           {44'h15?,1'b?},
           {36'h1,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_ACTION_CFG_1;
                 default: read_data = '0;
              endcase
           end
           {36'h1,4'b100?,4'h?,1'b?},
           {44'h1A?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_ACTION_CFG_2;
                 default: read_data = '0;
              endcase
           end
           {44'h1B?,1'b?},
           {36'h1,4'b110?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_ACTION_GLORT;
                 default: read_data = '0;
              endcase
           end
           {36'h1,4'b111?,4'h?,1'b?},
           {44'h20?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_ACTION_MIRROR;
                 default: read_data = '0;
              endcase
           end
           {44'h21?,1'b?},
           {36'h2,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_STATS;
                 default: read_data = '0;
              endcase
           end
           {44'h240,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTRL;
                 default: read_data = '0;
              endcase
           end
           {44'h240,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX0;
                 default: read_data = '0;
              endcase
           end
           {44'h241,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX1;
                 default: read_data = '0;
              endcase
           end
           {44'h241,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX2;
                 default: read_data = '0;
              endcase
           end
           {44'h242,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX3;
                 default: read_data = '0;
              endcase
           end
           {44'h242,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_CTX4;
                 default: read_data = '0;
              endcase
           end
           {44'h243,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM0;
                 default: read_data = '0;
              endcase
           end
           {44'h243,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM1;
                 default: read_data = '0;
              endcase
           end
           {44'h244,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM2;
                 default: read_data = '0;
              endcase
           end
           {44'h244,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM3;
                 default: read_data = '0;
              endcase
           end
           {44'h245,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADM4;
                 default: read_data = '0;
              endcase
           end
           {44'h245,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR0;
                 default: read_data = '0;
              endcase
           end
           {44'h246,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR1;
                 default: read_data = '0;
              endcase
           end
           {44'h246,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR2;
                 default: read_data = '0;
              endcase
           end
           {44'h247,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR3;
                 default: read_data = '0;
              endcase
           end
           {44'h247,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_SB_FID,TRIG_APPLY_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_DIRECT_MAP_ADR4;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {


// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
