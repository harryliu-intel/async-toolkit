// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

// INTEL TOP SECRET
// Copyright 2013 Intel Corporation. All Rights Reserved.
// $Id:  $

`ifndef NEW_ECC

// lintra -2056 "expression smaller than context"

package ecc_functions;

// Takes datain and tacks on the correct ecc in the correct position. 
function automatic logic [511:0] encode_ecc
  (input int           CBTS,        // number of ecc bits
   input int           WDTH,        // datapath bitwidth
   input logic [501:0] datain);     // datapath input
    logic [9:0]   chkout;
    logic [511:0] dataout;
    chkout = calculate_ecc(CBTS,datain);
    dataout[501:0] = datain;
    dataout[WDTH +: 10] = chkout;
    return(dataout);
endfunction


// The is a function that models the DW_ecc logic. Datapath and ecc
// bitwidths are set to the maximum supported by DW_ecc.
function automatic logic [9:0] calculate_ecc
  (input int           CBTS,      // number of ecc bits
   input logic [501:0] datain);   // data, rounded up to max bitwidth

    logic [9:0] chkout;

    // Vectors for 5 ecc bits
    if (CBTS==5) begin
      chkout[0] = ^(datain & 11'b11100101110) ^ 0;
      chkout[1] = ^(datain & 11'b10101010111) ^ 0;
      chkout[2] = ^(datain & 11'b11110011001) ^ 1;
      chkout[3] = ^(datain & 11'b01111100011) ^ 1;
      chkout[4] = ^(datain & 11'b00111111100) ^ 0;
    end
    else if (CBTS==6) begin
      chkout[0] = ^(datain & 26'b10101101110100101100101110) ^ 0;
      chkout[1] = ^(datain & 26'b11101011010001010101010111) ^ 0;
      chkout[2] = ^(datain & 26'b10100111111010011010011001) ^ 1;
      chkout[3] = ^(datain & 26'b10011110110011100011100011) ^ 1;
      chkout[4] = ^(datain & 26'b01111110011100000011111100) ^ 0;
      chkout[5] = ^(datain & 26'b11111110001111111100000000) ^ 0;
    end
    else if (CBTS==7) begin
      chkout[0] = ^(datain & 57'b101010011111010110110101010110100001011100100101111010001) ^ 0;
      chkout[1] = ^(datain & 57'b011101011011110101101000100010101010101110001010101010111) ^ 0;
      chkout[2] = ^(datain & 57'b010100111111010011011010110100110100110011010011010011001) ^ 1;
      chkout[3] = ^(datain & 57'b010011110111001111000110100111000111000110011100011100011) ^ 1;
      chkout[4] = ^(datain & 57'b001111110010111111000001111000000111111001100000011111100) ^ 0;
      chkout[5] = ^(datain & 57'b111111110001111111000000011111111000000001111111100000000) ^ 0;
      chkout[6] = ^(datain & 57'b111111110000000000111111111111111000000000000000011111111) ^ 0;
    end
    else if (CBTS==8) begin
      chkout[0] = ^(datain & 120'b101011010010101010101101111010100111010101010100111010101011010011010001101101001101000101001011001011100100101100101110) ^ 0;
      chkout[1] = ^(datain & 120'b111010101010001011101011010111010110100010111010110100010001010101010111000101010101011100010101010101110001010101010111) ^ 0;
      chkout[2] = ^(datain & 120'b101001100110101010100111110101001101101010101001101101011010011010011001101001101001100110100110100110011010011010011001) ^ 1;
      chkout[3] = ^(datain & 120'b100111100001101010011110110100111100011010100111100011010011100011100011001110001110001100111000111000110011100011100011) ^ 1;
      chkout[4] = ^(datain & 120'b011111100000011001111110010011111100000110011111100000111100000011111100110000001111110011000000111111001100000011111100) ^ 0;
      chkout[5] = ^(datain & 120'b111111100000000111111110001111111100000001111111100000001111111100000000111111110000000011111111000000001111111100000000) ^ 0;
      chkout[6] = ^(datain & 120'b000000011111111111111110000000000011111111111111100000001111111100000000000000001111111111111111000000000000000011111111) ^ 0;
      chkout[7] = ^(datain & 120'b000000011111111111111110001111111100000000000000011111110000000011111111111111110000000011111111000000000000000011111111) ^ 0;
    end
    else if (CBTS==9) begin
      chkout[0] = ^(datain & 247'b0110101010101101111010100111010100101011010010101101010011101010010101101001010110101001100101011010100101101010101011001001011110100011011010000101110101101000010111001001011110100011011010000101110010010111101000110110100001011100100101111010001) ^ 0;
      chkout[1] = ^(datain & 247'b0101000111101011010111010110100010111010101010001011101011010001011101010101000101110101010100010111010101010001111010100010101010101110001010101010111000101010101011100010101010101110001010101010111000101010101011100010101010101110001010101010111) ^ 0;
      chkout[2] = ^(datain & 247'b0011010110100111110101001101101010101001100110101010100110110101010100110011010101010011001101010101001100110101101001110100110100110011010011010011001101001101001100110100110100110011010011010011001101001101001100110100110100110011010011010011001) ^ 1;
      chkout[3] = ^(datain & 247'b0000110110011110110100111100011010100111100001101010011110001101010011110000110101001111000011010100111100001101100111100111000111000110011100011100011001110001110001100111000111000110011100011100011001110001110001100111000111000110011100011100011) ^ 1;
      chkout[4] = ^(datain & 247'b0000001101111110010011111100000110011111100000011001111110000011001111110000001100111111000000110011111100000011011111111000000111111001100000011111100110000001111110011000000111111001100000011111100110000001111110011000000111111001100000011111100) ^ 0;
      chkout[5] = ^(datain & 247'b0000000011111110001111111100000001111111100000000111111110000000111111110000000011111111111111110000000011111111000000000000000111111110000000011111111111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000) ^ 0;
      chkout[6] = ^(datain & 247'b1111111100000000001111111111111110000000000000000111111110000000111111111111111100000000000000001111111111111111000000000000000111111111111111100000000000000001111111111111111000000001111111100000000000000001111111111111111000000000000000011111111) ^ 0;
      chkout[7] = ^(datain & 247'b1111111100000000001111111100000001111111111111111000000001111111000000000000000011111111000000001111111111111111000000000000000111111111111111100000000111111110000000000000000111111110000000011111111111111110000000011111111000000000000000011111111) ^ 0;
      chkout[8] = ^(datain & 247'b1111111100000000001111111100000001111111111111111000000000000000111111111111111100000000111111110000000000000000111111111111111000000000000000011111111000000001111111111111111000000000000000011111111111111110000000011111111000000000000000011111111) ^ 0;
    end
    else if (CBTS==10) begin
      chkout[0] = ^(datain & 502'b1010110100101010101011011110101001110101010101001011010101010100111010101010100101101010101010010110101010101001011010101010100111010101010100101101010101010010110101010101001011010101010100101101010101010010110101010101001011010101010100111010101011010011010001101101001101000110110100110100011011010011010001101101001101000110110100110100011011010011010001101101001101000110110100110100011011010011010001101101001101000110110100110100011011010011010001101101001101000101001011001011100100101100101110) ^ 0;
      chkout[1] = ^(datain & 502'b1110101010100010111010110101110101101000101110101010100010111010110100010111010101010001011101010101000101110101010100010111010110100010111010101010001011101010101000101110101010100010111010101010001011101010101000101110101010100010111010110100010001010101010111000101010101011100010101010101110001010101010111000101010101011100010101010101110001010101010111000101010101011100010101010101110001010101010111000101010101011100010101010101110001010101010111000101010101011100010101010101110001010101010111) ^ 0;
      chkout[2] = ^(datain & 502'b1010011001101010101001111101010011011010101010011001101010101001101101010101001100110101010100110011010101010011001101010101001101101010101001100110101010100110011010101010011001101010101001100110101010100110011010101010011001101010101001101101011010011010011001101001101001100110100110100110011010011010011001101001101001100110100110100110011010011010011001101001101001100110100110100110011010011010011001101001101001100110100110100110011010011010011001101001101001100110100110100110011010011010011001) ^ 1;
      chkout[3] = ^(datain & 502'b1001111000011010100111101101001111000110101001111000011010100111100011010100111100001101010011110000110101001111000011010100111100011010100111100001101010011110000110101001111000011010100111100001101010011110000110101001111000011010100111100011010011100011100011001110001110001100111000111000110011100011100011001110001110001100111000111000110011100011100011001110001110001100111000111000110011100011100011001110001110001100111000111000110011100011100011001110001110001100111000111000110011100011100011) ^ 1;
      chkout[4] = ^(datain & 502'b0111111000000110011111100100111111000001100111111000000110011111100000110011111100000011001111110000001100111111000000110011111100000110011111100000011001111110000001100111111000000110011111100000011001111110000001100111111000000110011111100000111100000011111100110000001111110011000000111111001100000011111100110000001111110011000000111111001100000011111100110000001111110011000000111111001100000011111100110000001111110011000000111111001100000011111100110000001111110011000000111111001100000011111100) ^ 0;
      chkout[5] = ^(datain & 502'b1111111000000001111111100011111111000000011111111000000001111111100000001111111100000000000000001111111100000000111111111111111100000001111111100000000000000001111111100000000111111110000000011111111000000001111111111111111000000001111111100000001111111100000000111111110000000000000000111111110000000011111111000000001111111100000000111111111111111100000000111111110000000000000000111111110000000011111111111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000) ^ 0;
      chkout[6] = ^(datain & 502'b0000000111111111111111100000000000111111111111111000000001111111100000000000000011111111111111110000000000000000111111111111111100000000000000011111111111111110000000000000000111111110000000011111111111111110000000000000000111111111111111100000001111111100000000000000001111111111111111000000000000000011111111000000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000001111111100000000000000001111111111111111000000000000000011111111) ^ 0;
      chkout[7] = ^(datain & 502'b0000000111111111111111100011111111000000000000000111111110000000011111111111111100000000111111110000000000000000111111111111111100000000000000011111111000000001111111111111111000000001111111100000000000000001111111100000000111111111111111100000001111111100000000000000001111111100000000111111111111111100000000111111110000000000000000111111110000000011111111111111110000000000000000111111111111111100000000111111110000000000000000111111110000000011111111111111110000000011111111000000000000000011111111) ^ 0;
      chkout[8] = ^(datain & 502'b0000000111111111111111100011111111000000000000000111111111111111100000000000000011111111000000001111111111111111000000000000000011111111111111100000000111111110000000000000000111111111111111100000000000000001111111100000000111111111111111100000001111111100000000000000001111111100000000111111111111111100000000000000001111111111111111000000001111111100000000000000001111111111111111000000000000000011111111000000001111111111111111000000000000000011111111111111110000000011111111000000000000000011111111) ^ 0;
      chkout[9] = ^(datain & 502'b0000000111111111111111100011111111000000000000000111111111111111100000000000000011111111000000001111111111111111000000001111111100000000000000011111111000000001111111111111111000000000000000011111111111111110000000011111111000000000000000011111110000000011111111111111110000000011111111000000000000000011111111111111110000000000000000111111110000000011111111111111110000000011111111000000000000000011111111000000001111111111111111000000000000000011111111111111110000000011111111000000000000000011111111) ^ 0;
    end
    return(chkout);
endfunction

endpackage

// lintra +2056
   
`endif // !NEW_ECC
