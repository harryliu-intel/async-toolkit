///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_mesh_row_map.sv                                        
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_mesh_row_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_MESH_ROW_MAP_FF
`define RTLGEN_MBY_MESH_ROW_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_MESH_ROW_MAP_FF

`ifndef RTLGEN_MBY_MESH_ROW_MAP_EN_FF
`define RTLGEN_MBY_MESH_ROW_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_MESH_ROW_MAP_EN_FF

`ifndef RTLGEN_MBY_MESH_ROW_MAP_FF_RSTD
`define RTLGEN_MBY_MESH_ROW_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_MESH_ROW_MAP_FF_RSTD


module rtlgen_mby_mesh_row_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_MESH_ROW_MAP_EN_FF_RSTD
`define RTLGEN_MBY_MESH_ROW_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_mesh_row_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_MESH_ROW_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_MESH_ROW_MAP_FF_SYNCRST
`define RTLGEN_MBY_MESH_ROW_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_MESH_ROW_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_MESH_ROW_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_MESH_ROW_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_MESH_ROW_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_MESH_ROW_MAP_FF_BOTHRST
// `define RTLGEN_MBY_MESH_ROW_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_MESH_ROW_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_MESH_ROW_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_MESH_ROW_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_MESH_ROW_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_MESH_ROW_MAP_LATCH_LOW
`define RTLGEN_MBY_MESH_ROW_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_MESH_ROW_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_MESH_ROW_MAP_PH2_FF
`define RTLGEN_MBY_MESH_ROW_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_MESH_ROW_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_MESH_ROW_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_MESH_ROW_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_MESH_ROW_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_MESH_ROW_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_MESH_ROW_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_MESH_ROW_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_MESH_ROW_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_MESH_ROW_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_MESH_ROW_MAP_LATCH
`define RTLGEN_MBY_MESH_ROW_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_MESH_ROW_MAP_LATCH

`ifndef RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH
`define RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH

`ifndef RTLGEN_MBY_MESH_ROW_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_MESH_ROW_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_MESH_ROW_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_MESH_ROW_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_MESH_ROW_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_MESH_ROW_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_MESH_ROW_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_mesh_row_map ( //lintra s-2096
    // Clocks
    gated_clk,

    // Resets
    rst_n,


    // Register Inputs


    // Register Outputs
    MESH_ARB_RREQ_Y,
    MESH_ARB_RRSP_X,
    MESH_ARB_RRSP_Y,
    MESH_ARB_WREQ_Y,


    // Register signals for HandCoded registers



    // Config Access
    req,
    ack
    

);

import mby_mesh_row_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_MESH_ROW_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_MESH_ROW_MAP_MEM_ADDR_MSB:0] MBY_MESH_ROW_MAP_OFFSET = {MBY_MESH_ROW_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] MESH_SB_BAR = 3'b0;
parameter [7:0] MESH_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
`define MESH_ARB_RREQ_Y_CR_ADDR_def(INDEX) MESH_ARB_RREQ_Y_CR_ADDR``INDEX``[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_MESH_ROW_MAP_OFFSET[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
`define MESH_ARB_WREQ_Y_CR_ADDR_def(INDEX) MESH_ARB_WREQ_Y_CR_ADDR``INDEX``[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_MESH_ROW_MAP_OFFSET[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
`define MESH_ARB_RRSP_Y_CR_ADDR_def(INDEX) MESH_ARB_RRSP_Y_CR_ADDR``INDEX``[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_MESH_ROW_MAP_OFFSET[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
`define MESH_ARB_RRSP_X_CR_ADDR_def(INDEX) MESH_ARB_RRSP_X_CR_ADDR``INDEX``[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_MESH_ROW_MAP_OFFSET[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
localparam [7:0][MBY_MESH_ROW_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MESH_ARB_RREQ_Y_DECODE_ADDR = {`MESH_ARB_RREQ_Y_CR_ADDR_def([7]),`MESH_ARB_RREQ_Y_CR_ADDR_def([6]),`MESH_ARB_RREQ_Y_CR_ADDR_def([5]),`MESH_ARB_RREQ_Y_CR_ADDR_def([4]),`MESH_ARB_RREQ_Y_CR_ADDR_def([3]),`MESH_ARB_RREQ_Y_CR_ADDR_def([2]),`MESH_ARB_RREQ_Y_CR_ADDR_def([1]),`MESH_ARB_RREQ_Y_CR_ADDR_def([0])};
localparam [7:0][MBY_MESH_ROW_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MESH_ARB_WREQ_Y_DECODE_ADDR = {`MESH_ARB_WREQ_Y_CR_ADDR_def([7]),`MESH_ARB_WREQ_Y_CR_ADDR_def([6]),`MESH_ARB_WREQ_Y_CR_ADDR_def([5]),`MESH_ARB_WREQ_Y_CR_ADDR_def([4]),`MESH_ARB_WREQ_Y_CR_ADDR_def([3]),`MESH_ARB_WREQ_Y_CR_ADDR_def([2]),`MESH_ARB_WREQ_Y_CR_ADDR_def([1]),`MESH_ARB_WREQ_Y_CR_ADDR_def([0])};
localparam [7:0][MBY_MESH_ROW_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MESH_ARB_RRSP_Y_DECODE_ADDR = {`MESH_ARB_RRSP_Y_CR_ADDR_def([7]),`MESH_ARB_RRSP_Y_CR_ADDR_def([6]),`MESH_ARB_RRSP_Y_CR_ADDR_def([5]),`MESH_ARB_RRSP_Y_CR_ADDR_def([4]),`MESH_ARB_RRSP_Y_CR_ADDR_def([3]),`MESH_ARB_RRSP_Y_CR_ADDR_def([2]),`MESH_ARB_RRSP_Y_CR_ADDR_def([1]),`MESH_ARB_RRSP_Y_CR_ADDR_def([0])};
localparam [7:0][MBY_MESH_ROW_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MESH_ARB_RRSP_X_DECODE_ADDR = {`MESH_ARB_RRSP_X_CR_ADDR_def([7]),`MESH_ARB_RRSP_X_CR_ADDR_def([6]),`MESH_ARB_RRSP_X_CR_ADDR_def([5]),`MESH_ARB_RRSP_X_CR_ADDR_def([4]),`MESH_ARB_RRSP_X_CR_ADDR_def([3]),`MESH_ARB_RRSP_X_CR_ADDR_def([2]),`MESH_ARB_RRSP_X_CR_ADDR_def([1]),`MESH_ARB_RRSP_X_CR_ADDR_def([0])};

    // Clocks
input logic  gated_clk;

    // Resets
input logic  rst_n;


    // Register Inputs


    // Register Outputs
output MESH_ARB_RREQ_Y_t [7:0] MESH_ARB_RREQ_Y;
output MESH_ARB_RRSP_X_t [7:0] MESH_ARB_RRSP_X;
output MESH_ARB_RRSP_Y_t [7:0] MESH_ARB_RRSP_Y;
output MESH_ARB_WREQ_Y_t [7:0] MESH_ARB_WREQ_Y;


    // Register signals for HandCoded registers



    // Config Access
input mby_mesh_row_map_cr_req_t  req;
output mby_mesh_row_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_mesh_row_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_MESH_ROW_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_MESH_ROW_MAP_MEM;
assign case_req_addr_MBY_MESH_ROW_MAP_MEM = req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_mesh;
always_comb begin : sb_fid_cond_mesh_BLOCK
    unique casez (req_fid) 
		MESH_SB_FID: sb_fid_cond_mesh = 1;
		default: sb_fid_cond_mesh = 0;
    endcase 
end


logic sb_bar_cond_mesh;
always_comb begin : sb_bar_cond_mesh_BLOCK
    unique casez (req_bar) 
		MESH_SB_BAR: sb_bar_cond_mesh = 1;
		default: sb_bar_cond_mesh = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

//---------------------------------------------------------------------
// MESH_ARB_RREQ_Y Address Decode
logic [7:0] addr_decode_MESH_ARB_RREQ_Y;
logic [7:0] write_req_MESH_ARB_RREQ_Y;
always_comb begin
   addr_decode_MESH_ARB_RREQ_Y[0] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[0]) && req.valid ;
   addr_decode_MESH_ARB_RREQ_Y[1] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[1]) && req.valid ;
   addr_decode_MESH_ARB_RREQ_Y[2] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[2]) && req.valid ;
   addr_decode_MESH_ARB_RREQ_Y[3] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[3]) && req.valid ;
   addr_decode_MESH_ARB_RREQ_Y[4] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[4]) && req.valid ;
   addr_decode_MESH_ARB_RREQ_Y[5] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[5]) && req.valid ;
   addr_decode_MESH_ARB_RREQ_Y[6] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[6]) && req.valid ;
   addr_decode_MESH_ARB_RREQ_Y[7] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RREQ_Y_DECODE_ADDR[7]) && req.valid ;
   write_req_MESH_ARB_RREQ_Y[0] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[0] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RREQ_Y[1] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[1] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RREQ_Y[2] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[2] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RREQ_Y[3] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[3] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RREQ_Y[4] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[4] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RREQ_Y[5] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[5] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RREQ_Y[6] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[6] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RREQ_Y[7] = IsMEMWr && addr_decode_MESH_ARB_RREQ_Y[7] && sb_fid_cond_mesh && sb_bar_cond_mesh;
end

// ----------------------------------------------------------------------
// MESH_ARB_RREQ_Y.SB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RREQ_Y_SB_TO_SB;
always_comb begin
 up_MESH_ARB_RREQ_Y_SB_TO_SB[0] =
    ({1{write_req_MESH_ARB_RREQ_Y[0] }} &
    be[0:0]);
 up_MESH_ARB_RREQ_Y_SB_TO_SB[1] =
    ({1{write_req_MESH_ARB_RREQ_Y[1] }} &
    be[0:0]);
 up_MESH_ARB_RREQ_Y_SB_TO_SB[2] =
    ({1{write_req_MESH_ARB_RREQ_Y[2] }} &
    be[0:0]);
 up_MESH_ARB_RREQ_Y_SB_TO_SB[3] =
    ({1{write_req_MESH_ARB_RREQ_Y[3] }} &
    be[0:0]);
 up_MESH_ARB_RREQ_Y_SB_TO_SB[4] =
    ({1{write_req_MESH_ARB_RREQ_Y[4] }} &
    be[0:0]);
 up_MESH_ARB_RREQ_Y_SB_TO_SB[5] =
    ({1{write_req_MESH_ARB_RREQ_Y[5] }} &
    be[0:0]);
 up_MESH_ARB_RREQ_Y_SB_TO_SB[6] =
    ({1{write_req_MESH_ARB_RREQ_Y[6] }} &
    be[0:0]);
 up_MESH_ARB_RREQ_Y_SB_TO_SB[7] =
    ({1{write_req_MESH_ARB_RREQ_Y[7] }} &
    be[0:0]);
end

logic [7:0][7:0] nxt_MESH_ARB_RREQ_Y_SB_TO_SB;
always_comb begin
 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[0] = write_data[7:0];

 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[1] = write_data[7:0];

 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[2] = write_data[7:0];

 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[3] = write_data[7:0];

 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[4] = write_data[7:0];

 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[5] = write_data[7:0];

 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[6] = write_data[7:0];

 nxt_MESH_ARB_RREQ_Y_SB_TO_SB[7] = write_data[7:0];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[0][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[0][7:0], MESH_ARB_RREQ_Y[0].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[1][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[1][7:0], MESH_ARB_RREQ_Y[1].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[2][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[2][7:0], MESH_ARB_RREQ_Y[2].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[3][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[3][7:0], MESH_ARB_RREQ_Y[3].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[4][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[4][7:0], MESH_ARB_RREQ_Y[4].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[5][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[5][7:0], MESH_ARB_RREQ_Y[5].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[6][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[6][7:0], MESH_ARB_RREQ_Y[6].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_SB_TO_SB[7][0], nxt_MESH_ARB_RREQ_Y_SB_TO_SB[7][7:0], MESH_ARB_RREQ_Y[7].SB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RREQ_Y.EB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RREQ_Y_EB_TO_SB;
always_comb begin
 up_MESH_ARB_RREQ_Y_EB_TO_SB[0] =
    ({1{write_req_MESH_ARB_RREQ_Y[0] }} &
    be[1:1]);
 up_MESH_ARB_RREQ_Y_EB_TO_SB[1] =
    ({1{write_req_MESH_ARB_RREQ_Y[1] }} &
    be[1:1]);
 up_MESH_ARB_RREQ_Y_EB_TO_SB[2] =
    ({1{write_req_MESH_ARB_RREQ_Y[2] }} &
    be[1:1]);
 up_MESH_ARB_RREQ_Y_EB_TO_SB[3] =
    ({1{write_req_MESH_ARB_RREQ_Y[3] }} &
    be[1:1]);
 up_MESH_ARB_RREQ_Y_EB_TO_SB[4] =
    ({1{write_req_MESH_ARB_RREQ_Y[4] }} &
    be[1:1]);
 up_MESH_ARB_RREQ_Y_EB_TO_SB[5] =
    ({1{write_req_MESH_ARB_RREQ_Y[5] }} &
    be[1:1]);
 up_MESH_ARB_RREQ_Y_EB_TO_SB[6] =
    ({1{write_req_MESH_ARB_RREQ_Y[6] }} &
    be[1:1]);
 up_MESH_ARB_RREQ_Y_EB_TO_SB[7] =
    ({1{write_req_MESH_ARB_RREQ_Y[7] }} &
    be[1:1]);
end

logic [7:0][7:0] nxt_MESH_ARB_RREQ_Y_EB_TO_SB;
always_comb begin
 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[0] = write_data[15:8];

 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[1] = write_data[15:8];

 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[2] = write_data[15:8];

 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[3] = write_data[15:8];

 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[4] = write_data[15:8];

 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[5] = write_data[15:8];

 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[6] = write_data[15:8];

 nxt_MESH_ARB_RREQ_Y_EB_TO_SB[7] = write_data[15:8];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[0][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[0][7:0], MESH_ARB_RREQ_Y[0].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[1][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[1][7:0], MESH_ARB_RREQ_Y[1].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[2][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[2][7:0], MESH_ARB_RREQ_Y[2].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[3][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[3][7:0], MESH_ARB_RREQ_Y[3].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[4][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[4][7:0], MESH_ARB_RREQ_Y[4].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[5][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[5][7:0], MESH_ARB_RREQ_Y[5].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[6][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[6][7:0], MESH_ARB_RREQ_Y[6].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_SB[7][0], nxt_MESH_ARB_RREQ_Y_EB_TO_SB[7][7:0], MESH_ARB_RREQ_Y[7].EB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RREQ_Y.WB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RREQ_Y_WB_TO_SB;
always_comb begin
 up_MESH_ARB_RREQ_Y_WB_TO_SB[0] =
    ({1{write_req_MESH_ARB_RREQ_Y[0] }} &
    be[2:2]);
 up_MESH_ARB_RREQ_Y_WB_TO_SB[1] =
    ({1{write_req_MESH_ARB_RREQ_Y[1] }} &
    be[2:2]);
 up_MESH_ARB_RREQ_Y_WB_TO_SB[2] =
    ({1{write_req_MESH_ARB_RREQ_Y[2] }} &
    be[2:2]);
 up_MESH_ARB_RREQ_Y_WB_TO_SB[3] =
    ({1{write_req_MESH_ARB_RREQ_Y[3] }} &
    be[2:2]);
 up_MESH_ARB_RREQ_Y_WB_TO_SB[4] =
    ({1{write_req_MESH_ARB_RREQ_Y[4] }} &
    be[2:2]);
 up_MESH_ARB_RREQ_Y_WB_TO_SB[5] =
    ({1{write_req_MESH_ARB_RREQ_Y[5] }} &
    be[2:2]);
 up_MESH_ARB_RREQ_Y_WB_TO_SB[6] =
    ({1{write_req_MESH_ARB_RREQ_Y[6] }} &
    be[2:2]);
 up_MESH_ARB_RREQ_Y_WB_TO_SB[7] =
    ({1{write_req_MESH_ARB_RREQ_Y[7] }} &
    be[2:2]);
end

logic [7:0][7:0] nxt_MESH_ARB_RREQ_Y_WB_TO_SB;
always_comb begin
 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[0] = write_data[23:16];

 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[1] = write_data[23:16];

 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[2] = write_data[23:16];

 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[3] = write_data[23:16];

 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[4] = write_data[23:16];

 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[5] = write_data[23:16];

 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[6] = write_data[23:16];

 nxt_MESH_ARB_RREQ_Y_WB_TO_SB[7] = write_data[23:16];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[0][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[0][7:0], MESH_ARB_RREQ_Y[0].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[1][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[1][7:0], MESH_ARB_RREQ_Y[1].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[2][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[2][7:0], MESH_ARB_RREQ_Y[2].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[3][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[3][7:0], MESH_ARB_RREQ_Y[3].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[4][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[4][7:0], MESH_ARB_RREQ_Y[4].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[5][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[5][7:0], MESH_ARB_RREQ_Y[5].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[6][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[6][7:0], MESH_ARB_RREQ_Y[6].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_SB[7][0], nxt_MESH_ARB_RREQ_Y_WB_TO_SB[7][7:0], MESH_ARB_RREQ_Y[7].WB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RREQ_Y.NB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RREQ_Y_NB_TO_NB;
always_comb begin
 up_MESH_ARB_RREQ_Y_NB_TO_NB[0] =
    ({1{write_req_MESH_ARB_RREQ_Y[0] }} &
    be[3:3]);
 up_MESH_ARB_RREQ_Y_NB_TO_NB[1] =
    ({1{write_req_MESH_ARB_RREQ_Y[1] }} &
    be[3:3]);
 up_MESH_ARB_RREQ_Y_NB_TO_NB[2] =
    ({1{write_req_MESH_ARB_RREQ_Y[2] }} &
    be[3:3]);
 up_MESH_ARB_RREQ_Y_NB_TO_NB[3] =
    ({1{write_req_MESH_ARB_RREQ_Y[3] }} &
    be[3:3]);
 up_MESH_ARB_RREQ_Y_NB_TO_NB[4] =
    ({1{write_req_MESH_ARB_RREQ_Y[4] }} &
    be[3:3]);
 up_MESH_ARB_RREQ_Y_NB_TO_NB[5] =
    ({1{write_req_MESH_ARB_RREQ_Y[5] }} &
    be[3:3]);
 up_MESH_ARB_RREQ_Y_NB_TO_NB[6] =
    ({1{write_req_MESH_ARB_RREQ_Y[6] }} &
    be[3:3]);
 up_MESH_ARB_RREQ_Y_NB_TO_NB[7] =
    ({1{write_req_MESH_ARB_RREQ_Y[7] }} &
    be[3:3]);
end

logic [7:0][7:0] nxt_MESH_ARB_RREQ_Y_NB_TO_NB;
always_comb begin
 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[0] = write_data[31:24];

 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[1] = write_data[31:24];

 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[2] = write_data[31:24];

 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[3] = write_data[31:24];

 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[4] = write_data[31:24];

 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[5] = write_data[31:24];

 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[6] = write_data[31:24];

 nxt_MESH_ARB_RREQ_Y_NB_TO_NB[7] = write_data[31:24];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[0][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[0][7:0], MESH_ARB_RREQ_Y[0].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[1][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[1][7:0], MESH_ARB_RREQ_Y[1].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[2][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[2][7:0], MESH_ARB_RREQ_Y[2].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[3][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[3][7:0], MESH_ARB_RREQ_Y[3].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[4][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[4][7:0], MESH_ARB_RREQ_Y[4].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[5][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[5][7:0], MESH_ARB_RREQ_Y[5].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[6][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[6][7:0], MESH_ARB_RREQ_Y[6].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_NB_TO_NB[7][0], nxt_MESH_ARB_RREQ_Y_NB_TO_NB[7][7:0], MESH_ARB_RREQ_Y[7].NB_TO_NB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RREQ_Y.EB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RREQ_Y_EB_TO_NB;
always_comb begin
 up_MESH_ARB_RREQ_Y_EB_TO_NB[0] =
    ({1{write_req_MESH_ARB_RREQ_Y[0] }} &
    be[4:4]);
 up_MESH_ARB_RREQ_Y_EB_TO_NB[1] =
    ({1{write_req_MESH_ARB_RREQ_Y[1] }} &
    be[4:4]);
 up_MESH_ARB_RREQ_Y_EB_TO_NB[2] =
    ({1{write_req_MESH_ARB_RREQ_Y[2] }} &
    be[4:4]);
 up_MESH_ARB_RREQ_Y_EB_TO_NB[3] =
    ({1{write_req_MESH_ARB_RREQ_Y[3] }} &
    be[4:4]);
 up_MESH_ARB_RREQ_Y_EB_TO_NB[4] =
    ({1{write_req_MESH_ARB_RREQ_Y[4] }} &
    be[4:4]);
 up_MESH_ARB_RREQ_Y_EB_TO_NB[5] =
    ({1{write_req_MESH_ARB_RREQ_Y[5] }} &
    be[4:4]);
 up_MESH_ARB_RREQ_Y_EB_TO_NB[6] =
    ({1{write_req_MESH_ARB_RREQ_Y[6] }} &
    be[4:4]);
 up_MESH_ARB_RREQ_Y_EB_TO_NB[7] =
    ({1{write_req_MESH_ARB_RREQ_Y[7] }} &
    be[4:4]);
end

logic [7:0][7:0] nxt_MESH_ARB_RREQ_Y_EB_TO_NB;
always_comb begin
 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[0] = write_data[39:32];

 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[1] = write_data[39:32];

 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[2] = write_data[39:32];

 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[3] = write_data[39:32];

 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[4] = write_data[39:32];

 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[5] = write_data[39:32];

 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[6] = write_data[39:32];

 nxt_MESH_ARB_RREQ_Y_EB_TO_NB[7] = write_data[39:32];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[0][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[0][7:0], MESH_ARB_RREQ_Y[0].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[1][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[1][7:0], MESH_ARB_RREQ_Y[1].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[2][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[2][7:0], MESH_ARB_RREQ_Y[2].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[3][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[3][7:0], MESH_ARB_RREQ_Y[3].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[4][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[4][7:0], MESH_ARB_RREQ_Y[4].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[5][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[5][7:0], MESH_ARB_RREQ_Y[5].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[6][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[6][7:0], MESH_ARB_RREQ_Y[6].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_EB_TO_NB[7][0], nxt_MESH_ARB_RREQ_Y_EB_TO_NB[7][7:0], MESH_ARB_RREQ_Y[7].EB_TO_NB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RREQ_Y.WB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RREQ_Y_WB_TO_NB;
always_comb begin
 up_MESH_ARB_RREQ_Y_WB_TO_NB[0] =
    ({1{write_req_MESH_ARB_RREQ_Y[0] }} &
    be[5:5]);
 up_MESH_ARB_RREQ_Y_WB_TO_NB[1] =
    ({1{write_req_MESH_ARB_RREQ_Y[1] }} &
    be[5:5]);
 up_MESH_ARB_RREQ_Y_WB_TO_NB[2] =
    ({1{write_req_MESH_ARB_RREQ_Y[2] }} &
    be[5:5]);
 up_MESH_ARB_RREQ_Y_WB_TO_NB[3] =
    ({1{write_req_MESH_ARB_RREQ_Y[3] }} &
    be[5:5]);
 up_MESH_ARB_RREQ_Y_WB_TO_NB[4] =
    ({1{write_req_MESH_ARB_RREQ_Y[4] }} &
    be[5:5]);
 up_MESH_ARB_RREQ_Y_WB_TO_NB[5] =
    ({1{write_req_MESH_ARB_RREQ_Y[5] }} &
    be[5:5]);
 up_MESH_ARB_RREQ_Y_WB_TO_NB[6] =
    ({1{write_req_MESH_ARB_RREQ_Y[6] }} &
    be[5:5]);
 up_MESH_ARB_RREQ_Y_WB_TO_NB[7] =
    ({1{write_req_MESH_ARB_RREQ_Y[7] }} &
    be[5:5]);
end

logic [7:0][7:0] nxt_MESH_ARB_RREQ_Y_WB_TO_NB;
always_comb begin
 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[0] = write_data[47:40];

 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[1] = write_data[47:40];

 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[2] = write_data[47:40];

 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[3] = write_data[47:40];

 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[4] = write_data[47:40];

 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[5] = write_data[47:40];

 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[6] = write_data[47:40];

 nxt_MESH_ARB_RREQ_Y_WB_TO_NB[7] = write_data[47:40];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[0][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[0][7:0], MESH_ARB_RREQ_Y[0].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[1][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[1][7:0], MESH_ARB_RREQ_Y[1].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[2][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[2][7:0], MESH_ARB_RREQ_Y[2].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[3][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[3][7:0], MESH_ARB_RREQ_Y[3].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[4][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[4][7:0], MESH_ARB_RREQ_Y[4].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[5][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[5][7:0], MESH_ARB_RREQ_Y[5].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[6][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[6][7:0], MESH_ARB_RREQ_Y[6].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RREQ_Y_WB_TO_NB[7][0], nxt_MESH_ARB_RREQ_Y_WB_TO_NB[7][7:0], MESH_ARB_RREQ_Y[7].WB_TO_NB[7:0])

//---------------------------------------------------------------------
// MESH_ARB_WREQ_Y Address Decode
logic [7:0] addr_decode_MESH_ARB_WREQ_Y;
logic [7:0] write_req_MESH_ARB_WREQ_Y;
always_comb begin
   addr_decode_MESH_ARB_WREQ_Y[0] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[0]) && req.valid ;
   addr_decode_MESH_ARB_WREQ_Y[1] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[1]) && req.valid ;
   addr_decode_MESH_ARB_WREQ_Y[2] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[2]) && req.valid ;
   addr_decode_MESH_ARB_WREQ_Y[3] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[3]) && req.valid ;
   addr_decode_MESH_ARB_WREQ_Y[4] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[4]) && req.valid ;
   addr_decode_MESH_ARB_WREQ_Y[5] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[5]) && req.valid ;
   addr_decode_MESH_ARB_WREQ_Y[6] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[6]) && req.valid ;
   addr_decode_MESH_ARB_WREQ_Y[7] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_WREQ_Y_DECODE_ADDR[7]) && req.valid ;
   write_req_MESH_ARB_WREQ_Y[0] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[0] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_WREQ_Y[1] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[1] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_WREQ_Y[2] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[2] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_WREQ_Y[3] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[3] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_WREQ_Y[4] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[4] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_WREQ_Y[5] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[5] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_WREQ_Y[6] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[6] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_WREQ_Y[7] = IsMEMWr && addr_decode_MESH_ARB_WREQ_Y[7] && sb_fid_cond_mesh && sb_bar_cond_mesh;
end

// ----------------------------------------------------------------------
// MESH_ARB_WREQ_Y.SB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_WREQ_Y_SB_TO_SB;
always_comb begin
 up_MESH_ARB_WREQ_Y_SB_TO_SB[0] =
    ({1{write_req_MESH_ARB_WREQ_Y[0] }} &
    be[0:0]);
 up_MESH_ARB_WREQ_Y_SB_TO_SB[1] =
    ({1{write_req_MESH_ARB_WREQ_Y[1] }} &
    be[0:0]);
 up_MESH_ARB_WREQ_Y_SB_TO_SB[2] =
    ({1{write_req_MESH_ARB_WREQ_Y[2] }} &
    be[0:0]);
 up_MESH_ARB_WREQ_Y_SB_TO_SB[3] =
    ({1{write_req_MESH_ARB_WREQ_Y[3] }} &
    be[0:0]);
 up_MESH_ARB_WREQ_Y_SB_TO_SB[4] =
    ({1{write_req_MESH_ARB_WREQ_Y[4] }} &
    be[0:0]);
 up_MESH_ARB_WREQ_Y_SB_TO_SB[5] =
    ({1{write_req_MESH_ARB_WREQ_Y[5] }} &
    be[0:0]);
 up_MESH_ARB_WREQ_Y_SB_TO_SB[6] =
    ({1{write_req_MESH_ARB_WREQ_Y[6] }} &
    be[0:0]);
 up_MESH_ARB_WREQ_Y_SB_TO_SB[7] =
    ({1{write_req_MESH_ARB_WREQ_Y[7] }} &
    be[0:0]);
end

logic [7:0][7:0] nxt_MESH_ARB_WREQ_Y_SB_TO_SB;
always_comb begin
 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[0] = write_data[7:0];

 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[1] = write_data[7:0];

 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[2] = write_data[7:0];

 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[3] = write_data[7:0];

 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[4] = write_data[7:0];

 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[5] = write_data[7:0];

 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[6] = write_data[7:0];

 nxt_MESH_ARB_WREQ_Y_SB_TO_SB[7] = write_data[7:0];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[0][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[0][7:0], MESH_ARB_WREQ_Y[0].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[1][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[1][7:0], MESH_ARB_WREQ_Y[1].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[2][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[2][7:0], MESH_ARB_WREQ_Y[2].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[3][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[3][7:0], MESH_ARB_WREQ_Y[3].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[4][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[4][7:0], MESH_ARB_WREQ_Y[4].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[5][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[5][7:0], MESH_ARB_WREQ_Y[5].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[6][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[6][7:0], MESH_ARB_WREQ_Y[6].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_SB_TO_SB[7][0], nxt_MESH_ARB_WREQ_Y_SB_TO_SB[7][7:0], MESH_ARB_WREQ_Y[7].SB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_WREQ_Y.EB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_WREQ_Y_EB_TO_SB;
always_comb begin
 up_MESH_ARB_WREQ_Y_EB_TO_SB[0] =
    ({1{write_req_MESH_ARB_WREQ_Y[0] }} &
    be[1:1]);
 up_MESH_ARB_WREQ_Y_EB_TO_SB[1] =
    ({1{write_req_MESH_ARB_WREQ_Y[1] }} &
    be[1:1]);
 up_MESH_ARB_WREQ_Y_EB_TO_SB[2] =
    ({1{write_req_MESH_ARB_WREQ_Y[2] }} &
    be[1:1]);
 up_MESH_ARB_WREQ_Y_EB_TO_SB[3] =
    ({1{write_req_MESH_ARB_WREQ_Y[3] }} &
    be[1:1]);
 up_MESH_ARB_WREQ_Y_EB_TO_SB[4] =
    ({1{write_req_MESH_ARB_WREQ_Y[4] }} &
    be[1:1]);
 up_MESH_ARB_WREQ_Y_EB_TO_SB[5] =
    ({1{write_req_MESH_ARB_WREQ_Y[5] }} &
    be[1:1]);
 up_MESH_ARB_WREQ_Y_EB_TO_SB[6] =
    ({1{write_req_MESH_ARB_WREQ_Y[6] }} &
    be[1:1]);
 up_MESH_ARB_WREQ_Y_EB_TO_SB[7] =
    ({1{write_req_MESH_ARB_WREQ_Y[7] }} &
    be[1:1]);
end

logic [7:0][7:0] nxt_MESH_ARB_WREQ_Y_EB_TO_SB;
always_comb begin
 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[0] = write_data[15:8];

 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[1] = write_data[15:8];

 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[2] = write_data[15:8];

 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[3] = write_data[15:8];

 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[4] = write_data[15:8];

 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[5] = write_data[15:8];

 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[6] = write_data[15:8];

 nxt_MESH_ARB_WREQ_Y_EB_TO_SB[7] = write_data[15:8];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[0][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[0][7:0], MESH_ARB_WREQ_Y[0].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[1][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[1][7:0], MESH_ARB_WREQ_Y[1].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[2][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[2][7:0], MESH_ARB_WREQ_Y[2].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[3][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[3][7:0], MESH_ARB_WREQ_Y[3].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[4][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[4][7:0], MESH_ARB_WREQ_Y[4].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[5][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[5][7:0], MESH_ARB_WREQ_Y[5].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[6][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[6][7:0], MESH_ARB_WREQ_Y[6].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_SB[7][0], nxt_MESH_ARB_WREQ_Y_EB_TO_SB[7][7:0], MESH_ARB_WREQ_Y[7].EB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_WREQ_Y.WB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_WREQ_Y_WB_TO_SB;
always_comb begin
 up_MESH_ARB_WREQ_Y_WB_TO_SB[0] =
    ({1{write_req_MESH_ARB_WREQ_Y[0] }} &
    be[2:2]);
 up_MESH_ARB_WREQ_Y_WB_TO_SB[1] =
    ({1{write_req_MESH_ARB_WREQ_Y[1] }} &
    be[2:2]);
 up_MESH_ARB_WREQ_Y_WB_TO_SB[2] =
    ({1{write_req_MESH_ARB_WREQ_Y[2] }} &
    be[2:2]);
 up_MESH_ARB_WREQ_Y_WB_TO_SB[3] =
    ({1{write_req_MESH_ARB_WREQ_Y[3] }} &
    be[2:2]);
 up_MESH_ARB_WREQ_Y_WB_TO_SB[4] =
    ({1{write_req_MESH_ARB_WREQ_Y[4] }} &
    be[2:2]);
 up_MESH_ARB_WREQ_Y_WB_TO_SB[5] =
    ({1{write_req_MESH_ARB_WREQ_Y[5] }} &
    be[2:2]);
 up_MESH_ARB_WREQ_Y_WB_TO_SB[6] =
    ({1{write_req_MESH_ARB_WREQ_Y[6] }} &
    be[2:2]);
 up_MESH_ARB_WREQ_Y_WB_TO_SB[7] =
    ({1{write_req_MESH_ARB_WREQ_Y[7] }} &
    be[2:2]);
end

logic [7:0][7:0] nxt_MESH_ARB_WREQ_Y_WB_TO_SB;
always_comb begin
 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[0] = write_data[23:16];

 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[1] = write_data[23:16];

 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[2] = write_data[23:16];

 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[3] = write_data[23:16];

 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[4] = write_data[23:16];

 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[5] = write_data[23:16];

 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[6] = write_data[23:16];

 nxt_MESH_ARB_WREQ_Y_WB_TO_SB[7] = write_data[23:16];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[0][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[0][7:0], MESH_ARB_WREQ_Y[0].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[1][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[1][7:0], MESH_ARB_WREQ_Y[1].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[2][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[2][7:0], MESH_ARB_WREQ_Y[2].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[3][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[3][7:0], MESH_ARB_WREQ_Y[3].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[4][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[4][7:0], MESH_ARB_WREQ_Y[4].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[5][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[5][7:0], MESH_ARB_WREQ_Y[5].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[6][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[6][7:0], MESH_ARB_WREQ_Y[6].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_SB[7][0], nxt_MESH_ARB_WREQ_Y_WB_TO_SB[7][7:0], MESH_ARB_WREQ_Y[7].WB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_WREQ_Y.NB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_WREQ_Y_NB_TO_NB;
always_comb begin
 up_MESH_ARB_WREQ_Y_NB_TO_NB[0] =
    ({1{write_req_MESH_ARB_WREQ_Y[0] }} &
    be[3:3]);
 up_MESH_ARB_WREQ_Y_NB_TO_NB[1] =
    ({1{write_req_MESH_ARB_WREQ_Y[1] }} &
    be[3:3]);
 up_MESH_ARB_WREQ_Y_NB_TO_NB[2] =
    ({1{write_req_MESH_ARB_WREQ_Y[2] }} &
    be[3:3]);
 up_MESH_ARB_WREQ_Y_NB_TO_NB[3] =
    ({1{write_req_MESH_ARB_WREQ_Y[3] }} &
    be[3:3]);
 up_MESH_ARB_WREQ_Y_NB_TO_NB[4] =
    ({1{write_req_MESH_ARB_WREQ_Y[4] }} &
    be[3:3]);
 up_MESH_ARB_WREQ_Y_NB_TO_NB[5] =
    ({1{write_req_MESH_ARB_WREQ_Y[5] }} &
    be[3:3]);
 up_MESH_ARB_WREQ_Y_NB_TO_NB[6] =
    ({1{write_req_MESH_ARB_WREQ_Y[6] }} &
    be[3:3]);
 up_MESH_ARB_WREQ_Y_NB_TO_NB[7] =
    ({1{write_req_MESH_ARB_WREQ_Y[7] }} &
    be[3:3]);
end

logic [7:0][7:0] nxt_MESH_ARB_WREQ_Y_NB_TO_NB;
always_comb begin
 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[0] = write_data[31:24];

 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[1] = write_data[31:24];

 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[2] = write_data[31:24];

 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[3] = write_data[31:24];

 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[4] = write_data[31:24];

 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[5] = write_data[31:24];

 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[6] = write_data[31:24];

 nxt_MESH_ARB_WREQ_Y_NB_TO_NB[7] = write_data[31:24];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[0][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[0][7:0], MESH_ARB_WREQ_Y[0].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[1][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[1][7:0], MESH_ARB_WREQ_Y[1].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[2][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[2][7:0], MESH_ARB_WREQ_Y[2].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[3][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[3][7:0], MESH_ARB_WREQ_Y[3].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[4][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[4][7:0], MESH_ARB_WREQ_Y[4].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[5][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[5][7:0], MESH_ARB_WREQ_Y[5].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[6][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[6][7:0], MESH_ARB_WREQ_Y[6].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_NB_TO_NB[7][0], nxt_MESH_ARB_WREQ_Y_NB_TO_NB[7][7:0], MESH_ARB_WREQ_Y[7].NB_TO_NB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_WREQ_Y.EB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_WREQ_Y_EB_TO_NB;
always_comb begin
 up_MESH_ARB_WREQ_Y_EB_TO_NB[0] =
    ({1{write_req_MESH_ARB_WREQ_Y[0] }} &
    be[4:4]);
 up_MESH_ARB_WREQ_Y_EB_TO_NB[1] =
    ({1{write_req_MESH_ARB_WREQ_Y[1] }} &
    be[4:4]);
 up_MESH_ARB_WREQ_Y_EB_TO_NB[2] =
    ({1{write_req_MESH_ARB_WREQ_Y[2] }} &
    be[4:4]);
 up_MESH_ARB_WREQ_Y_EB_TO_NB[3] =
    ({1{write_req_MESH_ARB_WREQ_Y[3] }} &
    be[4:4]);
 up_MESH_ARB_WREQ_Y_EB_TO_NB[4] =
    ({1{write_req_MESH_ARB_WREQ_Y[4] }} &
    be[4:4]);
 up_MESH_ARB_WREQ_Y_EB_TO_NB[5] =
    ({1{write_req_MESH_ARB_WREQ_Y[5] }} &
    be[4:4]);
 up_MESH_ARB_WREQ_Y_EB_TO_NB[6] =
    ({1{write_req_MESH_ARB_WREQ_Y[6] }} &
    be[4:4]);
 up_MESH_ARB_WREQ_Y_EB_TO_NB[7] =
    ({1{write_req_MESH_ARB_WREQ_Y[7] }} &
    be[4:4]);
end

logic [7:0][7:0] nxt_MESH_ARB_WREQ_Y_EB_TO_NB;
always_comb begin
 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[0] = write_data[39:32];

 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[1] = write_data[39:32];

 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[2] = write_data[39:32];

 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[3] = write_data[39:32];

 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[4] = write_data[39:32];

 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[5] = write_data[39:32];

 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[6] = write_data[39:32];

 nxt_MESH_ARB_WREQ_Y_EB_TO_NB[7] = write_data[39:32];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[0][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[0][7:0], MESH_ARB_WREQ_Y[0].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[1][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[1][7:0], MESH_ARB_WREQ_Y[1].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[2][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[2][7:0], MESH_ARB_WREQ_Y[2].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[3][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[3][7:0], MESH_ARB_WREQ_Y[3].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[4][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[4][7:0], MESH_ARB_WREQ_Y[4].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[5][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[5][7:0], MESH_ARB_WREQ_Y[5].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[6][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[6][7:0], MESH_ARB_WREQ_Y[6].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_EB_TO_NB[7][0], nxt_MESH_ARB_WREQ_Y_EB_TO_NB[7][7:0], MESH_ARB_WREQ_Y[7].EB_TO_NB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_WREQ_Y.WB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_WREQ_Y_WB_TO_NB;
always_comb begin
 up_MESH_ARB_WREQ_Y_WB_TO_NB[0] =
    ({1{write_req_MESH_ARB_WREQ_Y[0] }} &
    be[5:5]);
 up_MESH_ARB_WREQ_Y_WB_TO_NB[1] =
    ({1{write_req_MESH_ARB_WREQ_Y[1] }} &
    be[5:5]);
 up_MESH_ARB_WREQ_Y_WB_TO_NB[2] =
    ({1{write_req_MESH_ARB_WREQ_Y[2] }} &
    be[5:5]);
 up_MESH_ARB_WREQ_Y_WB_TO_NB[3] =
    ({1{write_req_MESH_ARB_WREQ_Y[3] }} &
    be[5:5]);
 up_MESH_ARB_WREQ_Y_WB_TO_NB[4] =
    ({1{write_req_MESH_ARB_WREQ_Y[4] }} &
    be[5:5]);
 up_MESH_ARB_WREQ_Y_WB_TO_NB[5] =
    ({1{write_req_MESH_ARB_WREQ_Y[5] }} &
    be[5:5]);
 up_MESH_ARB_WREQ_Y_WB_TO_NB[6] =
    ({1{write_req_MESH_ARB_WREQ_Y[6] }} &
    be[5:5]);
 up_MESH_ARB_WREQ_Y_WB_TO_NB[7] =
    ({1{write_req_MESH_ARB_WREQ_Y[7] }} &
    be[5:5]);
end

logic [7:0][7:0] nxt_MESH_ARB_WREQ_Y_WB_TO_NB;
always_comb begin
 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[0] = write_data[47:40];

 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[1] = write_data[47:40];

 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[2] = write_data[47:40];

 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[3] = write_data[47:40];

 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[4] = write_data[47:40];

 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[5] = write_data[47:40];

 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[6] = write_data[47:40];

 nxt_MESH_ARB_WREQ_Y_WB_TO_NB[7] = write_data[47:40];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[0][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[0][7:0], MESH_ARB_WREQ_Y[0].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[1][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[1][7:0], MESH_ARB_WREQ_Y[1].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[2][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[2][7:0], MESH_ARB_WREQ_Y[2].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[3][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[3][7:0], MESH_ARB_WREQ_Y[3].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[4][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[4][7:0], MESH_ARB_WREQ_Y[4].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[5][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[5][7:0], MESH_ARB_WREQ_Y[5].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[6][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[6][7:0], MESH_ARB_WREQ_Y[6].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_WREQ_Y_WB_TO_NB[7][0], nxt_MESH_ARB_WREQ_Y_WB_TO_NB[7][7:0], MESH_ARB_WREQ_Y[7].WB_TO_NB[7:0])

//---------------------------------------------------------------------
// MESH_ARB_RRSP_Y Address Decode
logic [7:0] addr_decode_MESH_ARB_RRSP_Y;
logic [7:0] write_req_MESH_ARB_RRSP_Y;
always_comb begin
   addr_decode_MESH_ARB_RRSP_Y[0] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[0]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_Y[1] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[1]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_Y[2] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[2]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_Y[3] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[3]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_Y[4] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[4]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_Y[5] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[5]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_Y[6] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[6]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_Y[7] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_Y_DECODE_ADDR[7]) && req.valid ;
   write_req_MESH_ARB_RRSP_Y[0] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[0] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_Y[1] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[1] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_Y[2] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[2] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_Y[3] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[3] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_Y[4] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[4] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_Y[5] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[5] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_Y[6] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[6] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_Y[7] = IsMEMWr && addr_decode_MESH_ARB_RRSP_Y[7] && sb_fid_cond_mesh && sb_bar_cond_mesh;
end

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.MEM_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_MEM_TO_SB;
always_comb begin
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_Y_MEM_TO_SB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[0:0]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_MEM_TO_SB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[0] = write_data[7:0];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[1] = write_data[7:0];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[2] = write_data[7:0];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[3] = write_data[7:0];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[4] = write_data[7:0];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[5] = write_data[7:0];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[6] = write_data[7:0];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[7] = write_data[7:0];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[0][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[0][7:0], MESH_ARB_RRSP_Y[0].MEM_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[1][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[1][7:0], MESH_ARB_RRSP_Y[1].MEM_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[2][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[2][7:0], MESH_ARB_RRSP_Y[2].MEM_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[3][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[3][7:0], MESH_ARB_RRSP_Y[3].MEM_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[4][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[4][7:0], MESH_ARB_RRSP_Y[4].MEM_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[5][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[5][7:0], MESH_ARB_RRSP_Y[5].MEM_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[6][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[6][7:0], MESH_ARB_RRSP_Y[6].MEM_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_SB[7][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_SB[7][7:0], MESH_ARB_RRSP_Y[7].MEM_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.SB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_SB_TO_SB;
always_comb begin
 up_MESH_ARB_RRSP_Y_SB_TO_SB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_Y_SB_TO_SB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_Y_SB_TO_SB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_Y_SB_TO_SB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_Y_SB_TO_SB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_Y_SB_TO_SB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_Y_SB_TO_SB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_Y_SB_TO_SB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[1:1]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_SB_TO_SB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[0] = write_data[15:8];

 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[1] = write_data[15:8];

 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[2] = write_data[15:8];

 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[3] = write_data[15:8];

 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[4] = write_data[15:8];

 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[5] = write_data[15:8];

 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[6] = write_data[15:8];

 nxt_MESH_ARB_RRSP_Y_SB_TO_SB[7] = write_data[15:8];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[0][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[0][7:0], MESH_ARB_RRSP_Y[0].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[1][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[1][7:0], MESH_ARB_RRSP_Y[1].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[2][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[2][7:0], MESH_ARB_RRSP_Y[2].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[3][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[3][7:0], MESH_ARB_RRSP_Y[3].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[4][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[4][7:0], MESH_ARB_RRSP_Y[4].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[5][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[5][7:0], MESH_ARB_RRSP_Y[5].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[6][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[6][7:0], MESH_ARB_RRSP_Y[6].SB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_SB_TO_SB[7][0], nxt_MESH_ARB_RRSP_Y_SB_TO_SB[7][7:0], MESH_ARB_RRSP_Y[7].SB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.EB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_EB_TO_SB;
always_comb begin
 up_MESH_ARB_RRSP_Y_EB_TO_SB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_Y_EB_TO_SB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_Y_EB_TO_SB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_Y_EB_TO_SB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_Y_EB_TO_SB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_Y_EB_TO_SB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_Y_EB_TO_SB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_Y_EB_TO_SB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[2:2]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_EB_TO_SB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[0] = write_data[23:16];

 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[1] = write_data[23:16];

 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[2] = write_data[23:16];

 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[3] = write_data[23:16];

 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[4] = write_data[23:16];

 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[5] = write_data[23:16];

 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[6] = write_data[23:16];

 nxt_MESH_ARB_RRSP_Y_EB_TO_SB[7] = write_data[23:16];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[0][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[0][7:0], MESH_ARB_RRSP_Y[0].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[1][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[1][7:0], MESH_ARB_RRSP_Y[1].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[2][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[2][7:0], MESH_ARB_RRSP_Y[2].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[3][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[3][7:0], MESH_ARB_RRSP_Y[3].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[4][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[4][7:0], MESH_ARB_RRSP_Y[4].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[5][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[5][7:0], MESH_ARB_RRSP_Y[5].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[6][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[6][7:0], MESH_ARB_RRSP_Y[6].EB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_SB[7][0], nxt_MESH_ARB_RRSP_Y_EB_TO_SB[7][7:0], MESH_ARB_RRSP_Y[7].EB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.WB_TO_SB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_WB_TO_SB;
always_comb begin
 up_MESH_ARB_RRSP_Y_WB_TO_SB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_Y_WB_TO_SB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_Y_WB_TO_SB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_Y_WB_TO_SB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_Y_WB_TO_SB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_Y_WB_TO_SB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_Y_WB_TO_SB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_Y_WB_TO_SB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[3:3]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_WB_TO_SB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[0] = write_data[31:24];

 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[1] = write_data[31:24];

 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[2] = write_data[31:24];

 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[3] = write_data[31:24];

 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[4] = write_data[31:24];

 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[5] = write_data[31:24];

 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[6] = write_data[31:24];

 nxt_MESH_ARB_RRSP_Y_WB_TO_SB[7] = write_data[31:24];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[0][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[0][7:0], MESH_ARB_RRSP_Y[0].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[1][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[1][7:0], MESH_ARB_RRSP_Y[1].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[2][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[2][7:0], MESH_ARB_RRSP_Y[2].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[3][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[3][7:0], MESH_ARB_RRSP_Y[3].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[4][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[4][7:0], MESH_ARB_RRSP_Y[4].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[5][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[5][7:0], MESH_ARB_RRSP_Y[5].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[6][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[6][7:0], MESH_ARB_RRSP_Y[6].WB_TO_SB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_SB[7][0], nxt_MESH_ARB_RRSP_Y_WB_TO_SB[7][7:0], MESH_ARB_RRSP_Y[7].WB_TO_SB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.MEM_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_MEM_TO_NB;
always_comb begin
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_Y_MEM_TO_NB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[4:4]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_MEM_TO_NB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[0] = write_data[39:32];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[1] = write_data[39:32];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[2] = write_data[39:32];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[3] = write_data[39:32];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[4] = write_data[39:32];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[5] = write_data[39:32];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[6] = write_data[39:32];

 nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[7] = write_data[39:32];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[0][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[0][7:0], MESH_ARB_RRSP_Y[0].MEM_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[1][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[1][7:0], MESH_ARB_RRSP_Y[1].MEM_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[2][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[2][7:0], MESH_ARB_RRSP_Y[2].MEM_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[3][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[3][7:0], MESH_ARB_RRSP_Y[3].MEM_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[4][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[4][7:0], MESH_ARB_RRSP_Y[4].MEM_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[5][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[5][7:0], MESH_ARB_RRSP_Y[5].MEM_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[6][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[6][7:0], MESH_ARB_RRSP_Y[6].MEM_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_MEM_TO_NB[7][0], nxt_MESH_ARB_RRSP_Y_MEM_TO_NB[7][7:0], MESH_ARB_RRSP_Y[7].MEM_TO_NB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.NB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_NB_TO_NB;
always_comb begin
 up_MESH_ARB_RRSP_Y_NB_TO_NB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_Y_NB_TO_NB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_Y_NB_TO_NB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_Y_NB_TO_NB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_Y_NB_TO_NB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_Y_NB_TO_NB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_Y_NB_TO_NB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_Y_NB_TO_NB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[5:5]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_NB_TO_NB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[0] = write_data[47:40];

 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[1] = write_data[47:40];

 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[2] = write_data[47:40];

 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[3] = write_data[47:40];

 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[4] = write_data[47:40];

 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[5] = write_data[47:40];

 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[6] = write_data[47:40];

 nxt_MESH_ARB_RRSP_Y_NB_TO_NB[7] = write_data[47:40];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[0][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[0][7:0], MESH_ARB_RRSP_Y[0].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[1][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[1][7:0], MESH_ARB_RRSP_Y[1].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[2][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[2][7:0], MESH_ARB_RRSP_Y[2].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[3][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[3][7:0], MESH_ARB_RRSP_Y[3].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[4][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[4][7:0], MESH_ARB_RRSP_Y[4].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[5][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[5][7:0], MESH_ARB_RRSP_Y[5].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[6][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[6][7:0], MESH_ARB_RRSP_Y[6].NB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_NB_TO_NB[7][0], nxt_MESH_ARB_RRSP_Y_NB_TO_NB[7][7:0], MESH_ARB_RRSP_Y[7].NB_TO_NB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.EB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_EB_TO_NB;
always_comb begin
 up_MESH_ARB_RRSP_Y_EB_TO_NB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_Y_EB_TO_NB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_Y_EB_TO_NB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_Y_EB_TO_NB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_Y_EB_TO_NB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_Y_EB_TO_NB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_Y_EB_TO_NB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_Y_EB_TO_NB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[6:6]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_EB_TO_NB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[0] = write_data[55:48];

 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[1] = write_data[55:48];

 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[2] = write_data[55:48];

 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[3] = write_data[55:48];

 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[4] = write_data[55:48];

 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[5] = write_data[55:48];

 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[6] = write_data[55:48];

 nxt_MESH_ARB_RRSP_Y_EB_TO_NB[7] = write_data[55:48];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[0][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[0][7:0], MESH_ARB_RRSP_Y[0].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[1][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[1][7:0], MESH_ARB_RRSP_Y[1].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[2][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[2][7:0], MESH_ARB_RRSP_Y[2].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[3][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[3][7:0], MESH_ARB_RRSP_Y[3].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[4][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[4][7:0], MESH_ARB_RRSP_Y[4].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[5][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[5][7:0], MESH_ARB_RRSP_Y[5].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[6][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[6][7:0], MESH_ARB_RRSP_Y[6].EB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_EB_TO_NB[7][0], nxt_MESH_ARB_RRSP_Y_EB_TO_NB[7][7:0], MESH_ARB_RRSP_Y[7].EB_TO_NB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_Y.WB_TO_NB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_Y_WB_TO_NB;
always_comb begin
 up_MESH_ARB_RRSP_Y_WB_TO_NB[0] =
    ({1{write_req_MESH_ARB_RRSP_Y[0] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_Y_WB_TO_NB[1] =
    ({1{write_req_MESH_ARB_RRSP_Y[1] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_Y_WB_TO_NB[2] =
    ({1{write_req_MESH_ARB_RRSP_Y[2] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_Y_WB_TO_NB[3] =
    ({1{write_req_MESH_ARB_RRSP_Y[3] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_Y_WB_TO_NB[4] =
    ({1{write_req_MESH_ARB_RRSP_Y[4] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_Y_WB_TO_NB[5] =
    ({1{write_req_MESH_ARB_RRSP_Y[5] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_Y_WB_TO_NB[6] =
    ({1{write_req_MESH_ARB_RRSP_Y[6] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_Y_WB_TO_NB[7] =
    ({1{write_req_MESH_ARB_RRSP_Y[7] }} &
    be[7:7]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_Y_WB_TO_NB;
always_comb begin
 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[0] = write_data[63:56];

 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[1] = write_data[63:56];

 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[2] = write_data[63:56];

 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[3] = write_data[63:56];

 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[4] = write_data[63:56];

 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[5] = write_data[63:56];

 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[6] = write_data[63:56];

 nxt_MESH_ARB_RRSP_Y_WB_TO_NB[7] = write_data[63:56];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[0][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[0][7:0], MESH_ARB_RRSP_Y[0].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[1][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[1][7:0], MESH_ARB_RRSP_Y[1].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[2][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[2][7:0], MESH_ARB_RRSP_Y[2].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[3][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[3][7:0], MESH_ARB_RRSP_Y[3].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[4][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[4][7:0], MESH_ARB_RRSP_Y[4].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[5][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[5][7:0], MESH_ARB_RRSP_Y[5].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[6][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[6][7:0], MESH_ARB_RRSP_Y[6].WB_TO_NB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_Y_WB_TO_NB[7][0], nxt_MESH_ARB_RRSP_Y_WB_TO_NB[7][7:0], MESH_ARB_RRSP_Y[7].WB_TO_NB[7:0])

//---------------------------------------------------------------------
// MESH_ARB_RRSP_X Address Decode
logic [7:0] addr_decode_MESH_ARB_RRSP_X;
logic [7:0] write_req_MESH_ARB_RRSP_X;
always_comb begin
   addr_decode_MESH_ARB_RRSP_X[0] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[0]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_X[1] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[1]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_X[2] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[2]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_X[3] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[3]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_X[4] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[4]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_X[5] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[5]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_X[6] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[6]) && req.valid ;
   addr_decode_MESH_ARB_RRSP_X[7] = (req_addr[MBY_MESH_ROW_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MESH_ARB_RRSP_X_DECODE_ADDR[7]) && req.valid ;
   write_req_MESH_ARB_RRSP_X[0] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[0] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_X[1] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[1] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_X[2] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[2] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_X[3] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[3] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_X[4] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[4] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_X[5] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[5] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_X[6] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[6] && sb_fid_cond_mesh && sb_bar_cond_mesh;
   write_req_MESH_ARB_RRSP_X[7] = IsMEMWr && addr_decode_MESH_ARB_RRSP_X[7] && sb_fid_cond_mesh && sb_bar_cond_mesh;
end

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.MEM_TO_EB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_MEM_TO_EB;
always_comb begin
 up_MESH_ARB_RRSP_X_MEM_TO_EB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_X_MEM_TO_EB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_X_MEM_TO_EB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_X_MEM_TO_EB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_X_MEM_TO_EB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_X_MEM_TO_EB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_X_MEM_TO_EB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[0:0]);
 up_MESH_ARB_RRSP_X_MEM_TO_EB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[0:0]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_MEM_TO_EB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[0] = write_data[7:0];

 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[1] = write_data[7:0];

 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[2] = write_data[7:0];

 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[3] = write_data[7:0];

 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[4] = write_data[7:0];

 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[5] = write_data[7:0];

 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[6] = write_data[7:0];

 nxt_MESH_ARB_RRSP_X_MEM_TO_EB[7] = write_data[7:0];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[0][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[0][7:0], MESH_ARB_RRSP_X[0].MEM_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[1][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[1][7:0], MESH_ARB_RRSP_X[1].MEM_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[2][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[2][7:0], MESH_ARB_RRSP_X[2].MEM_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[3][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[3][7:0], MESH_ARB_RRSP_X[3].MEM_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[4][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[4][7:0], MESH_ARB_RRSP_X[4].MEM_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[5][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[5][7:0], MESH_ARB_RRSP_X[5].MEM_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[6][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[6][7:0], MESH_ARB_RRSP_X[6].MEM_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_EB[7][0], nxt_MESH_ARB_RRSP_X_MEM_TO_EB[7][7:0], MESH_ARB_RRSP_X[7].MEM_TO_EB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.EB_TO_EB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_EB_TO_EB;
always_comb begin
 up_MESH_ARB_RRSP_X_EB_TO_EB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_X_EB_TO_EB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_X_EB_TO_EB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_X_EB_TO_EB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_X_EB_TO_EB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_X_EB_TO_EB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_X_EB_TO_EB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[1:1]);
 up_MESH_ARB_RRSP_X_EB_TO_EB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[1:1]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_EB_TO_EB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_EB_TO_EB[0] = write_data[15:8];

 nxt_MESH_ARB_RRSP_X_EB_TO_EB[1] = write_data[15:8];

 nxt_MESH_ARB_RRSP_X_EB_TO_EB[2] = write_data[15:8];

 nxt_MESH_ARB_RRSP_X_EB_TO_EB[3] = write_data[15:8];

 nxt_MESH_ARB_RRSP_X_EB_TO_EB[4] = write_data[15:8];

 nxt_MESH_ARB_RRSP_X_EB_TO_EB[5] = write_data[15:8];

 nxt_MESH_ARB_RRSP_X_EB_TO_EB[6] = write_data[15:8];

 nxt_MESH_ARB_RRSP_X_EB_TO_EB[7] = write_data[15:8];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[0][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[0][7:0], MESH_ARB_RRSP_X[0].EB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[1][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[1][7:0], MESH_ARB_RRSP_X[1].EB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[2][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[2][7:0], MESH_ARB_RRSP_X[2].EB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[3][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[3][7:0], MESH_ARB_RRSP_X[3].EB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[4][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[4][7:0], MESH_ARB_RRSP_X[4].EB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[5][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[5][7:0], MESH_ARB_RRSP_X[5].EB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[6][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[6][7:0], MESH_ARB_RRSP_X[6].EB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_EB_TO_EB[7][0], nxt_MESH_ARB_RRSP_X_EB_TO_EB[7][7:0], MESH_ARB_RRSP_X[7].EB_TO_EB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.SB_TO_EB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_SB_TO_EB;
always_comb begin
 up_MESH_ARB_RRSP_X_SB_TO_EB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_X_SB_TO_EB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_X_SB_TO_EB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_X_SB_TO_EB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_X_SB_TO_EB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_X_SB_TO_EB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_X_SB_TO_EB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[2:2]);
 up_MESH_ARB_RRSP_X_SB_TO_EB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[2:2]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_SB_TO_EB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_SB_TO_EB[0] = write_data[23:16];

 nxt_MESH_ARB_RRSP_X_SB_TO_EB[1] = write_data[23:16];

 nxt_MESH_ARB_RRSP_X_SB_TO_EB[2] = write_data[23:16];

 nxt_MESH_ARB_RRSP_X_SB_TO_EB[3] = write_data[23:16];

 nxt_MESH_ARB_RRSP_X_SB_TO_EB[4] = write_data[23:16];

 nxt_MESH_ARB_RRSP_X_SB_TO_EB[5] = write_data[23:16];

 nxt_MESH_ARB_RRSP_X_SB_TO_EB[6] = write_data[23:16];

 nxt_MESH_ARB_RRSP_X_SB_TO_EB[7] = write_data[23:16];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[0][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[0][7:0], MESH_ARB_RRSP_X[0].SB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[1][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[1][7:0], MESH_ARB_RRSP_X[1].SB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[2][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[2][7:0], MESH_ARB_RRSP_X[2].SB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[3][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[3][7:0], MESH_ARB_RRSP_X[3].SB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[4][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[4][7:0], MESH_ARB_RRSP_X[4].SB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[5][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[5][7:0], MESH_ARB_RRSP_X[5].SB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[6][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[6][7:0], MESH_ARB_RRSP_X[6].SB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_EB[7][0], nxt_MESH_ARB_RRSP_X_SB_TO_EB[7][7:0], MESH_ARB_RRSP_X[7].SB_TO_EB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.NB_TO_EB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_NB_TO_EB;
always_comb begin
 up_MESH_ARB_RRSP_X_NB_TO_EB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_X_NB_TO_EB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_X_NB_TO_EB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_X_NB_TO_EB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_X_NB_TO_EB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_X_NB_TO_EB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_X_NB_TO_EB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[3:3]);
 up_MESH_ARB_RRSP_X_NB_TO_EB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[3:3]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_NB_TO_EB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_NB_TO_EB[0] = write_data[31:24];

 nxt_MESH_ARB_RRSP_X_NB_TO_EB[1] = write_data[31:24];

 nxt_MESH_ARB_RRSP_X_NB_TO_EB[2] = write_data[31:24];

 nxt_MESH_ARB_RRSP_X_NB_TO_EB[3] = write_data[31:24];

 nxt_MESH_ARB_RRSP_X_NB_TO_EB[4] = write_data[31:24];

 nxt_MESH_ARB_RRSP_X_NB_TO_EB[5] = write_data[31:24];

 nxt_MESH_ARB_RRSP_X_NB_TO_EB[6] = write_data[31:24];

 nxt_MESH_ARB_RRSP_X_NB_TO_EB[7] = write_data[31:24];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[0][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[0][7:0], MESH_ARB_RRSP_X[0].NB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[1][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[1][7:0], MESH_ARB_RRSP_X[1].NB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[2][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[2][7:0], MESH_ARB_RRSP_X[2].NB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[3][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[3][7:0], MESH_ARB_RRSP_X[3].NB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[4][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[4][7:0], MESH_ARB_RRSP_X[4].NB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[5][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[5][7:0], MESH_ARB_RRSP_X[5].NB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[6][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[6][7:0], MESH_ARB_RRSP_X[6].NB_TO_EB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_EB[7][0], nxt_MESH_ARB_RRSP_X_NB_TO_EB[7][7:0], MESH_ARB_RRSP_X[7].NB_TO_EB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.MEM_TO_WB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_MEM_TO_WB;
always_comb begin
 up_MESH_ARB_RRSP_X_MEM_TO_WB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_X_MEM_TO_WB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_X_MEM_TO_WB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_X_MEM_TO_WB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_X_MEM_TO_WB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_X_MEM_TO_WB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_X_MEM_TO_WB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[4:4]);
 up_MESH_ARB_RRSP_X_MEM_TO_WB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[4:4]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_MEM_TO_WB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[0] = write_data[39:32];

 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[1] = write_data[39:32];

 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[2] = write_data[39:32];

 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[3] = write_data[39:32];

 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[4] = write_data[39:32];

 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[5] = write_data[39:32];

 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[6] = write_data[39:32];

 nxt_MESH_ARB_RRSP_X_MEM_TO_WB[7] = write_data[39:32];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[0][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[0][7:0], MESH_ARB_RRSP_X[0].MEM_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[1][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[1][7:0], MESH_ARB_RRSP_X[1].MEM_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[2][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[2][7:0], MESH_ARB_RRSP_X[2].MEM_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[3][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[3][7:0], MESH_ARB_RRSP_X[3].MEM_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[4][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[4][7:0], MESH_ARB_RRSP_X[4].MEM_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[5][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[5][7:0], MESH_ARB_RRSP_X[5].MEM_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[6][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[6][7:0], MESH_ARB_RRSP_X[6].MEM_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_MEM_TO_WB[7][0], nxt_MESH_ARB_RRSP_X_MEM_TO_WB[7][7:0], MESH_ARB_RRSP_X[7].MEM_TO_WB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.WB_TO_WB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_WB_TO_WB;
always_comb begin
 up_MESH_ARB_RRSP_X_WB_TO_WB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_X_WB_TO_WB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_X_WB_TO_WB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_X_WB_TO_WB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_X_WB_TO_WB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_X_WB_TO_WB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_X_WB_TO_WB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[5:5]);
 up_MESH_ARB_RRSP_X_WB_TO_WB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[5:5]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_WB_TO_WB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_WB_TO_WB[0] = write_data[47:40];

 nxt_MESH_ARB_RRSP_X_WB_TO_WB[1] = write_data[47:40];

 nxt_MESH_ARB_RRSP_X_WB_TO_WB[2] = write_data[47:40];

 nxt_MESH_ARB_RRSP_X_WB_TO_WB[3] = write_data[47:40];

 nxt_MESH_ARB_RRSP_X_WB_TO_WB[4] = write_data[47:40];

 nxt_MESH_ARB_RRSP_X_WB_TO_WB[5] = write_data[47:40];

 nxt_MESH_ARB_RRSP_X_WB_TO_WB[6] = write_data[47:40];

 nxt_MESH_ARB_RRSP_X_WB_TO_WB[7] = write_data[47:40];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[0][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[0][7:0], MESH_ARB_RRSP_X[0].WB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[1][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[1][7:0], MESH_ARB_RRSP_X[1].WB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[2][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[2][7:0], MESH_ARB_RRSP_X[2].WB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[3][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[3][7:0], MESH_ARB_RRSP_X[3].WB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[4][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[4][7:0], MESH_ARB_RRSP_X[4].WB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[5][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[5][7:0], MESH_ARB_RRSP_X[5].WB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[6][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[6][7:0], MESH_ARB_RRSP_X[6].WB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_WB_TO_WB[7][0], nxt_MESH_ARB_RRSP_X_WB_TO_WB[7][7:0], MESH_ARB_RRSP_X[7].WB_TO_WB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.SB_TO_WB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_SB_TO_WB;
always_comb begin
 up_MESH_ARB_RRSP_X_SB_TO_WB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_X_SB_TO_WB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_X_SB_TO_WB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_X_SB_TO_WB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_X_SB_TO_WB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_X_SB_TO_WB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_X_SB_TO_WB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[6:6]);
 up_MESH_ARB_RRSP_X_SB_TO_WB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[6:6]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_SB_TO_WB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_SB_TO_WB[0] = write_data[55:48];

 nxt_MESH_ARB_RRSP_X_SB_TO_WB[1] = write_data[55:48];

 nxt_MESH_ARB_RRSP_X_SB_TO_WB[2] = write_data[55:48];

 nxt_MESH_ARB_RRSP_X_SB_TO_WB[3] = write_data[55:48];

 nxt_MESH_ARB_RRSP_X_SB_TO_WB[4] = write_data[55:48];

 nxt_MESH_ARB_RRSP_X_SB_TO_WB[5] = write_data[55:48];

 nxt_MESH_ARB_RRSP_X_SB_TO_WB[6] = write_data[55:48];

 nxt_MESH_ARB_RRSP_X_SB_TO_WB[7] = write_data[55:48];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[0][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[0][7:0], MESH_ARB_RRSP_X[0].SB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[1][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[1][7:0], MESH_ARB_RRSP_X[1].SB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[2][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[2][7:0], MESH_ARB_RRSP_X[2].SB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[3][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[3][7:0], MESH_ARB_RRSP_X[3].SB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[4][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[4][7:0], MESH_ARB_RRSP_X[4].SB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[5][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[5][7:0], MESH_ARB_RRSP_X[5].SB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[6][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[6][7:0], MESH_ARB_RRSP_X[6].SB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_SB_TO_WB[7][0], nxt_MESH_ARB_RRSP_X_SB_TO_WB[7][7:0], MESH_ARB_RRSP_X[7].SB_TO_WB[7:0])

// ----------------------------------------------------------------------
// MESH_ARB_RRSP_X.NB_TO_WB x8 RW, using RW template.
logic [7:0][0:0] up_MESH_ARB_RRSP_X_NB_TO_WB;
always_comb begin
 up_MESH_ARB_RRSP_X_NB_TO_WB[0] =
    ({1{write_req_MESH_ARB_RRSP_X[0] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_X_NB_TO_WB[1] =
    ({1{write_req_MESH_ARB_RRSP_X[1] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_X_NB_TO_WB[2] =
    ({1{write_req_MESH_ARB_RRSP_X[2] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_X_NB_TO_WB[3] =
    ({1{write_req_MESH_ARB_RRSP_X[3] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_X_NB_TO_WB[4] =
    ({1{write_req_MESH_ARB_RRSP_X[4] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_X_NB_TO_WB[5] =
    ({1{write_req_MESH_ARB_RRSP_X[5] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_X_NB_TO_WB[6] =
    ({1{write_req_MESH_ARB_RRSP_X[6] }} &
    be[7:7]);
 up_MESH_ARB_RRSP_X_NB_TO_WB[7] =
    ({1{write_req_MESH_ARB_RRSP_X[7] }} &
    be[7:7]);
end

logic [7:0][7:0] nxt_MESH_ARB_RRSP_X_NB_TO_WB;
always_comb begin
 nxt_MESH_ARB_RRSP_X_NB_TO_WB[0] = write_data[63:56];

 nxt_MESH_ARB_RRSP_X_NB_TO_WB[1] = write_data[63:56];

 nxt_MESH_ARB_RRSP_X_NB_TO_WB[2] = write_data[63:56];

 nxt_MESH_ARB_RRSP_X_NB_TO_WB[3] = write_data[63:56];

 nxt_MESH_ARB_RRSP_X_NB_TO_WB[4] = write_data[63:56];

 nxt_MESH_ARB_RRSP_X_NB_TO_WB[5] = write_data[63:56];

 nxt_MESH_ARB_RRSP_X_NB_TO_WB[6] = write_data[63:56];

 nxt_MESH_ARB_RRSP_X_NB_TO_WB[7] = write_data[63:56];

end


`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[0][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[0][7:0], MESH_ARB_RRSP_X[0].NB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[1][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[1][7:0], MESH_ARB_RRSP_X[1].NB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[2][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[2][7:0], MESH_ARB_RRSP_X[2].NB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[3][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[3][7:0], MESH_ARB_RRSP_X[3].NB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[4][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[4][7:0], MESH_ARB_RRSP_X[4].NB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[5][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[5][7:0], MESH_ARB_RRSP_X[5].NB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[6][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[6][7:0], MESH_ARB_RRSP_X[6].NB_TO_WB[7:0])
`RTLGEN_MBY_MESH_ROW_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MESH_ARB_RRSP_X_NB_TO_WB[7][0], nxt_MESH_ARB_RRSP_X_NB_TO_WB[7][7:0], MESH_ARB_RRSP_X[7].NB_TO_WB[7:0])

// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_MESH_ROW_MAP_MEM) 
           MESH_ARB_RREQ_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_MESH_ROW_MAP_MEM) 
           MESH_ARB_RREQ_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_MESH_ROW_MAP_MEM) 
           MESH_ARB_RREQ_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[0]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[1]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[2]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[3]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[4]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[5]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[6]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RREQ_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RREQ_Y[7]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[0]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[1]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[2]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[3]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[4]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[5]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[6]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_WREQ_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_WREQ_Y[7]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[0]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[1]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[2]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[3]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[4]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[5]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[6]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_Y_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_Y[7]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[0]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[1]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[2]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[3]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[4]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[5]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[6]};
                 default: read_data = '0;
              endcase
           end
           MESH_ARB_RRSP_X_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {MESH_SB_FID,MESH_SB_BAR}: read_data = {MESH_ARB_RRSP_X[7]};
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    MESH_ARB_RREQ_Y[0].reserved0 = '0;
    MESH_ARB_RREQ_Y[1].reserved0 = '0;
    MESH_ARB_RREQ_Y[2].reserved0 = '0;
    MESH_ARB_RREQ_Y[3].reserved0 = '0;
    MESH_ARB_RREQ_Y[4].reserved0 = '0;
    MESH_ARB_RREQ_Y[5].reserved0 = '0;
    MESH_ARB_RREQ_Y[6].reserved0 = '0;
    MESH_ARB_RREQ_Y[7].reserved0 = '0;
    MESH_ARB_WREQ_Y[0].reserved0 = '0;
    MESH_ARB_WREQ_Y[1].reserved0 = '0;
    MESH_ARB_WREQ_Y[2].reserved0 = '0;
    MESH_ARB_WREQ_Y[3].reserved0 = '0;
    MESH_ARB_WREQ_Y[4].reserved0 = '0;
    MESH_ARB_WREQ_Y[5].reserved0 = '0;
    MESH_ARB_WREQ_Y[6].reserved0 = '0;
    MESH_ARB_WREQ_Y[7].reserved0 = '0;
end

// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
