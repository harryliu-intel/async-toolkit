///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///
// -------------------------------------------------------------------
// -- Intel Proprietary
// -- Copyright (C) 2018 Intel Corporation
// -- All Rights Reserved
// -------------------------------------------------------------------
// -- Author : Jon Bagge <jon.bagge@intel.com>
// -- Project Name : Madison Bay
// -- Description : Ingress to RX PPE interface
// --
// -------------------------------------------------------------------

interface igr_rx_ppe_if
import shared_pkg::*;
();
igr_rx_ppe_tail_t   intf0_tail;     //tail information for interface 0
igr_rx_ppe_head_t   intf0_head;     //head segment for interface 0
logic               intf0_ack;      //segment acknowledge for interface 0

igr_rx_ppe_tail_t   intf1_tail;     //tail information for interface 1
igr_rx_ppe_head_t   intf1_head;     //head segment for interface 1
logic               intf1_ack;      //segment acknowledge for interface 1

modport igr(
    output  intf0_tail,
    output  intf0_head,
    input   intf0_ack,
    output  intf1_tail,
    output  intf1_head,
    input   intf1_ack
);

modport ppe(
    input   intf0_tail,
    input   intf0_head,
    output  intf0_ack,
    input   intf1_tail,
    input   intf1_head,
    output  intf1_ack
);

endinterface: igr_rx_ppe_if
