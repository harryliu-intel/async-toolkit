begin
delay_cclk(1);
end
