// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0


///
///  INTEL CONFIDENTIAL
///
///  Copyright 2015 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///
//-----------------------------------------------------------------------------
// Title         : 
// Project       : Fox River
//-----------------------------------------------------------------------------
// File          : fxr_10b_ecc_cor.sv
// Author        : neuman.paul  <paul.neuman@intel.com>
// Created       : 17.06.2015  d.m.y
//-----------------------------------------------------------------------------
// Description :  !)b ECC Gen
//-----------------------------------------------------------------------------
// Intel Proprietary
// Copyright (C) 2015 Intel Corporation
// All Rights Reserved
//------------------------------------------------------------------------------

module fxr_10b_ecc_cor (
  input  logic [255:0]     data_in, 
  input  logic [9:0]       chk_in,
  input  logic [3:0]       par_in,
  input  logic             ecc_val,
  output logic [255:0]     data_out,
  output logic [9:0]       chk_out,
  output logic [9:0]       syn,
  output                   sbe,
  output                   mbe
);

  typedef struct packed {
    logic [9:0]  id;
  }  ten_bit;

  logic [255:0]            datain;
  logic [9:0]              syndrome_x;
  logic [9:0]              syndrome;
  logic [255:0]            correctionvector;
  logic [1:0]              parity_err;
  logic [255:0]            data_mask;
  logic                    syn_sbe;
  
  assign datain = data_in ;
  
  fxr_10b_ecc_gen fxr_10b_ecc_gen0(
     .data  (data_in),  
     .chk   (syndrome_x)
  );
  
  assign parity_err[0] =  (par_in[1] ^ (^datain[127:64])) | (par_in[0] ^ (^datain[63:0])) ;
  assign parity_err[1] =  (par_in[3] ^ (^datain[255:192])) | (par_in[2] ^ (^datain[191:128])) ;
  
  assign syndrome = (syndrome_x ^ chk_in) & {10{ecc_val}};

  assign syn = syndrome ;
  
  assign chk_out = syn_sbe ? (chk_in ^ syndrome) : chk_in ;
  
  assign syn_sbe = ((syndrome == 10'h200) | (syndrome == 10'h100) | (syndrome == 10'h080) | (syndrome == 10'h040) | (syndrome == 10'h020) | 
                    (syndrome == 10'h010) | (syndrome == 10'h008) | (syndrome == 10'h004) | (syndrome == 10'h002) | (syndrome == 10'h001)) ;
  
  assign sbe = (^syndrome) & (parity_err[1] | parity_err[0] | syn_sbe);
  
  assign mbe = (|syndrome) & ~((^syndrome) & (parity_err[1] | parity_err[0] | syn_sbe)) ;
  
  assign correctionvector = data_mask ;
        
  assign data_out = ((sbe == 1'b1) & (syn_sbe == 1'b0)) ? (datain ^ correctionvector) : datain ;
  
  always_comb
  unique case(syndrome)
      10'b0001100001 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000001 ; 
      10'b0011000010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000002 ; 
      10'b0110000100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000004 ; 
      10'b1100001000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000008 ;
      10'b1000110000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000010 ; 
      10'b0010100001 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000020 ; 
      10'b0101000010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000040 ; 
      10'b1010000100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000080 ;
      10'b0100101000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000100 ; 
      10'b1001010000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000200 ; 
      10'b0000100011 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000400 ; 
      10'b0001000110 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000800 ;
      10'b0010001100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000001000 ; 
      10'b0100011000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000002000 ; 
      10'b1000010001 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000004000 ; 
      10'b0000100101 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000008000 ;
      10'b0001001010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000010000 ; 
      10'b0010010100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000020000 ; 
      10'b0100001001 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000040000 ; 
      10'b1000010010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000080000 ;
      10'b0001100111 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000100000 ; 
      10'b0011001011 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000200000 ; 
      10'b0110010011 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000400000 ; 
      10'b1100001101 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000800000 ;
      10'b1000110101 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000001000000 ; 
      10'b0010111001 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000002000000 ; 
      10'b0101001110 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000004000000 ; 
      10'b1010010110 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000008000000 ;
      10'b0100111010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000010000000 ; 
      10'b1001011100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000020000000 ; 
      10'b0011100011 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000040000000 ; 
      10'b0101100110 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000080000000 ;
      10'b1001101100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000100000000 ; 
      10'b0110111000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000200000000 ; 
      10'b1010110001 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000400000000 ; 
      10'b1100100101 : data_mask = 256'h0000000000000000000000000000000000000000000000000000000800000000 ;
      10'b0111001010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000001000000000 ; 
      10'b1011010100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000002000000000 ; 
      10'b1101001001 : data_mask = 256'h0000000000000000000000000000000000000000000000000000004000000000 ; 
      10'b1110010010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000008000000000 ;
      10'b0000001101 : data_mask = 256'h0000000000000000000000000000000000000000000000000000010000000000 ; 
      10'b0000010011 : data_mask = 256'h0000000000000000000000000000000000000000000000000000020000000000 ; 
      10'b0110100000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000040000000000 ; 
      10'b1001100000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000080000000000 ;
      10'b1111000010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000100000000000 ; 
      10'b0001100010 : data_mask = 256'h0000000000000000000000000000000000000000000000000000200000000000 ; 
      10'b0011000100 : data_mask = 256'h0000000000000000000000000000000000000000000000000000400000000000 ; 
      10'b0110001000 : data_mask = 256'h0000000000000000000000000000000000000000000000000000800000000000 ;
      10'b1100010000 : data_mask = 256'h0000000000000000000000000000000000000000000000000001000000000000 ; 
      10'b1000100001 : data_mask = 256'h0000000000000000000000000000000000000000000000000002000000000000 ; 
      10'b0010100010 : data_mask = 256'h0000000000000000000000000000000000000000000000000004000000000000 ; 
      10'b0101000100 : data_mask = 256'h0000000000000000000000000000000000000000000000000008000000000000 ;
      10'b1010001000 : data_mask = 256'h0000000000000000000000000000000000000000000000000010000000000000 ; 
      10'b0100110000 : data_mask = 256'h0000000000000000000000000000000000000000000000000020000000000000 ; 
      10'b1001000001 : data_mask = 256'h0000000000000000000000000000000000000000000000000040000000000000 ; 
      10'b0001000011 : data_mask = 256'h0000000000000000000000000000000000000000000000000080000000000000 ;
      10'b0010000110 : data_mask = 256'h0000000000000000000000000000000000000000000000000100000000000000 ; 
      10'b0100001100 : data_mask = 256'h0000000000000000000000000000000000000000000000000200000000000000 ; 
      10'b1000011000 : data_mask = 256'h0000000000000000000000000000000000000000000000000400000000000000 ; 
      10'b0000110001 : data_mask = 256'h0000000000000000000000000000000000000000000000000800000000000000 ;
      10'b0001000101 : data_mask = 256'h0000000000000000000000000000000000000000000000001000000000000000 ; 
      10'b0010001010 : data_mask = 256'h0000000000000000000000000000000000000000000000002000000000000000 ; 
      10'b0100010100 : data_mask = 256'h0000000000000000000000000000000000000000000000004000000000000000 ; 
      10'b1000001001 : data_mask = 256'h0000000000000000000000000000000000000000000000008000000000000000 ;
      10'b0000110010 : data_mask = 256'h0000000000000000000000000000000000000000000000010000000000000000 ; 
      10'b0011000111 : data_mask = 256'h0000000000000000000000000000000000000000000000020000000000000000 ; 
      10'b0110001011 : data_mask = 256'h0000000000000000000000000000000000000000000000040000000000000000 ; 
      10'b1100010011 : data_mask = 256'h0000000000000000000000000000000000000000000000080000000000000000 ;
      10'b1000101101 : data_mask = 256'h0000000000000000000000000000000000000000000000100000000000000000 ; 
      10'b0001110101 : data_mask = 256'h0000000000000000000000000000000000000000000000200000000000000000 ; 
      10'b0101011001 : data_mask = 256'h0000000000000000000000000000000000000000000000400000000000000000 ; 
      10'b1010001110 : data_mask = 256'h0000000000000000000000000000000000000000000000800000000000000000 ;
      10'b0100110110 : data_mask = 256'h0000000000000000000000000000000000000000000001000000000000000000 ; 
      10'b1001011010 : data_mask = 256'h0000000000000000000000000000000000000000000002000000000000000000 ; 
      10'b0010111100 : data_mask = 256'h0000000000000000000000000000000000000000000004000000000000000000 ; 
      10'b0011100110 : data_mask = 256'h0000000000000000000000000000000000000000000008000000000000000000 ;
      10'b0101101100 : data_mask = 256'h0000000000000000000000000000000000000000000010000000000000000000 ; 
      10'b1001111000 : data_mask = 256'h0000000000000000000000000000000000000000000020000000000000000000 ; 
      10'b0110110001 : data_mask = 256'h0000000000000000000000000000000000000000000040000000000000000000 ; 
      10'b1010100011 : data_mask = 256'h0000000000000000000000000000000000000000000080000000000000000000 ;
      10'b1100101010 : data_mask = 256'h0000000000000000000000000000000000000000000100000000000000000000 ; 
      10'b0111010100 : data_mask = 256'h0000000000000000000000000000000000000000000200000000000000000000 ; 
      10'b1011001001 : data_mask = 256'h0000000000000000000000000000000000000000000400000000000000000000 ; 
      10'b1101010010 : data_mask = 256'h0000000000000000000000000000000000000000000800000000000000000000 ;
      10'b1110000101 : data_mask = 256'h0000000000000000000000000000000000000000001000000000000000000000 ; 
      10'b0000001011 : data_mask = 256'h0000000000000000000000000000000000000000002000000000000000000000 ; 
      10'b0000011100 : data_mask = 256'h0000000000000000000000000000000000000000004000000000000000000000 ; 
      10'b0101100000 : data_mask = 256'h0000000000000000000000000000000000000000008000000000000000000000 ;
      10'b1110000000 : data_mask = 256'h0000000000000000000000000000000000000000010000000000000000000000 ;
      10'b1011110000 : data_mask = 256'h0000000000000000000000000000000000000000020000000000000000000000 ; 
      10'b0001100100 : data_mask = 256'h0000000000000000000000000000000000000000040000000000000000000000 ; 
      10'b0011001000 : data_mask = 256'h0000000000000000000000000000000000000000080000000000000000000000 ;
      10'b0110010000 : data_mask = 256'h0000000000000000000000000000000000000000100000000000000000000000 ; 
      10'b1100000001 : data_mask = 256'h0000000000000000000000000000000000000000200000000000000000000000 ; 
      10'b1000100010 : data_mask = 256'h0000000000000000000000000000000000000000400000000000000000000000 ; 
      10'b0010100100 : data_mask = 256'h0000000000000000000000000000000000000000800000000000000000000000 ;
      10'b0101001000 : data_mask = 256'h0000000000000000000000000000000000000001000000000000000000000000 ; 
      10'b1010010000 : data_mask = 256'h0000000000000000000000000000000000000002000000000000000000000000 ; 
      10'b0100100001 : data_mask = 256'h0000000000000000000000000000000000000004000000000000000000000000 ; 
      10'b1001000010 : data_mask = 256'h0000000000000000000000000000000000000008000000000000000000000000 ;
      10'b0010000011 : data_mask = 256'h0000000000000000000000000000000000000010000000000000000000000000 ; 
      10'b0100000110 : data_mask = 256'h0000000000000000000000000000000000000020000000000000000000000000 ; 
      10'b1000001100 : data_mask = 256'h0000000000000000000000000000000000000040000000000000000000000000 ; 
      10'b0000111000 : data_mask = 256'h0000000000000000000000000000000000000080000000000000000000000000 ;
      10'b0001010001 : data_mask = 256'h0000000000000000000000000000000000000100000000000000000000000000 ; 
      10'b0010000101 : data_mask = 256'h0000000000000000000000000000000000000200000000000000000000000000 ; 
      10'b0100001010 : data_mask = 256'h0000000000000000000000000000000000000400000000000000000000000000 ; 
      10'b1000010100 : data_mask = 256'h0000000000000000000000000000000000000800000000000000000000000000 ;
      10'b0000101001 : data_mask = 256'h0000000000000000000000000000000000001000000000000000000000000000 ; 
      10'b0001010010 : data_mask = 256'h0000000000000000000000000000000000002000000000000000000000000000 ; 
      10'b0110000111 : data_mask = 256'h0000000000000000000000000000000000004000000000000000000000000000 ; 
      10'b1100001011 : data_mask = 256'h0000000000000000000000000000000000008000000000000000000000000000 ;
      10'b1000110011 : data_mask = 256'h0000000000000000000000000000000000010000000000000000000000000000 ; 
      10'b0001101101 : data_mask = 256'h0000000000000000000000000000000000020000000000000000000000000000 ; 
      10'b0011010101 : data_mask = 256'h0000000000000000000000000000000000040000000000000000000000000000 ; 
      10'b1010011001 : data_mask = 256'h0000000000000000000000000000000000080000000000000000000000000000 ;
      10'b0100101110 : data_mask = 256'h0000000000000000000000000000000000100000000000000000000000000000 ; 
      10'b1001010110 : data_mask = 256'h0000000000000000000000000000000000200000000000000000000000000000 ; 
      10'b0010111010 : data_mask = 256'h0000000000000000000000000000000000400000000000000000000000000000 ; 
      10'b0101011100 : data_mask = 256'h0000000000000000000000000000000000800000000000000000000000000000 ;
      10'b0011101100 : data_mask = 256'h0000000000000000000000000000000001000000000000000000000000000000 ; 
      10'b0101111000 : data_mask = 256'h0000000000000000000000000000000002000000000000000000000000000000 ; 
      10'b1001110001 : data_mask = 256'h0000000000000000000000000000000004000000000000000000000000000000 ; 
      10'b0110100011 : data_mask = 256'h0000000000000000000000000000000008000000000000000000000000000000 ;
      10'b1010100110 : data_mask = 256'h0000000000000000000000000000000010000000000000000000000000000000 ; 
      10'b1100110100 : data_mask = 256'h0000000000000000000000000000000020000000000000000000000000000000 ; 
      10'b0111001001 : data_mask = 256'h0000000000000000000000000000000040000000000000000000000000000000 ; 
      10'b1011010010 : data_mask = 256'h0000000000000000000000000000000080000000000000000000000000000000 ;
      10'b1101000101 : data_mask = 256'h0000000000000000000000000000000100000000000000000000000000000000 ; 
      10'b1110001010 : data_mask = 256'h0000000000000000000000000000000200000000000000000000000000000000 ; 
      10'b0000011010 : data_mask = 256'h0000000000000000000000000000000400000000000000000000000000000000 ; 
      10'b0000000111 : data_mask = 256'h0000000000000000000000000000000800000000000000000000000000000000 ;
      10'b1101000000 : data_mask = 256'h0000000000000000000000000000001000000000000000000000000000000000 ; 
      10'b0011100000 : data_mask = 256'h0000000000000000000000000000002000000000000000000000000000000000 ; 
      10'b1110100100 : data_mask = 256'h0000000000000000000000000000004000000000000000000000000000000000 ; 
      10'b0001101000 : data_mask = 256'h0000000000000000000000000000008000000000000000000000000000000000 ;
      10'b0011010000 : data_mask = 256'h0000000000000000000000000000010000000000000000000000000000000000 ; 
      10'b0110000001 : data_mask = 256'h0000000000000000000000000000020000000000000000000000000000000000 ; 
      10'b1100000010 : data_mask = 256'h0000000000000000000000000000040000000000000000000000000000000000 ; 
      10'b1000100100 : data_mask = 256'h0000000000000000000000000000080000000000000000000000000000000000 ;
      10'b0010101000 : data_mask = 256'h0000000000000000000000000000100000000000000000000000000000000000 ; 
      10'b0101010000 : data_mask = 256'h0000000000000000000000000000200000000000000000000000000000000000 ; 
      10'b1010000001 : data_mask = 256'h0000000000000000000000000000400000000000000000000000000000000000 ; 
      10'b0100100010 : data_mask = 256'h0000000000000000000000000000800000000000000000000000000000000000 ;
      10'b1001000100 : data_mask = 256'h0000000000000000000000000001000000000000000000000000000000000000 ; 
      10'b0100000011 : data_mask = 256'h0000000000000000000000000002000000000000000000000000000000000000 ; 
      10'b1000000110 : data_mask = 256'h0000000000000000000000000004000000000000000000000000000000000000 ; 
      10'b0000101100 : data_mask = 256'h0000000000000000000000000008000000000000000000000000000000000000 ;
      10'b0001011000 : data_mask = 256'h0000000000000000000000000010000000000000000000000000000000000000 ; 
      10'b0010010001 : data_mask = 256'h0000000000000000000000000020000000000000000000000000000000000000 ; 
      10'b0100000101 : data_mask = 256'h0000000000000000000000000040000000000000000000000000000000000000 ; 
      10'b1000001010 : data_mask = 256'h0000000000000000000000000080000000000000000000000000000000000000 ;
      10'b0000110100 : data_mask = 256'h0000000000000000000000000100000000000000000000000000000000000000 ; 
      10'b0001001001 : data_mask = 256'h0000000000000000000000000200000000000000000000000000000000000000 ; 
      10'b0010010010 : data_mask = 256'h0000000000000000000000000400000000000000000000000000000000000000 ; 
      10'b1100000111 : data_mask = 256'h0000000000000000000000000800000000000000000000000000000000000000 ;
      10'b1000101011 : data_mask = 256'h0000000000000000000000001000000000000000000000000000000000000000 ; 
      10'b0001110011 : data_mask = 256'h0000000000000000000000002000000000000000000000000000000000000000 ; 
      10'b0011001101 : data_mask = 256'h0000000000000000000000004000000000000000000000000000000000000000 ; 
      10'b0110010101 : data_mask = 256'h0000000000000000000000008000000000000000000000000000000000000000 ;
      10'b0100111001 : data_mask = 256'h0000000000000000000000010000000000000000000000000000000000000000 ; 
      10'b1001001110 : data_mask = 256'h0000000000000000000000020000000000000000000000000000000000000000 ; 
      10'b0010110110 : data_mask = 256'h0000000000000000000000040000000000000000000000000000000000000000 ; 
      10'b0101011010 : data_mask = 256'h0000000000000000000000080000000000000000000000000000000000000000 ;
      10'b1010011100 : data_mask = 256'h0000000000000000000000100000000000000000000000000000000000000000 ; 
      10'b0011111000 : data_mask = 256'h0000000000000000000000200000000000000000000000000000000000000000 ; 
      10'b0101110001 : data_mask = 256'h0000000000000000000000400000000000000000000000000000000000000000 ; 
      10'b1001100011 : data_mask = 256'h0000000000000000000000800000000000000000000000000000000000000000 ;
      10'b0110100110 : data_mask = 256'h0000000000000000000001000000000000000000000000000000000000000000 ; 
      10'b1010101100 : data_mask = 256'h0000000000000000000002000000000000000000000000000000000000000000 ; 
      10'b1100101001 : data_mask = 256'h0000000000000000000004000000000000000000000000000000000000000000 ; 
      10'b0111010010 : data_mask = 256'h0000000000000000000008000000000000000000000000000000000000000000 ;
      10'b1011000101 : data_mask = 256'h0000000000000000000010000000000000000000000000000000000000000000 ; 
      10'b1101001010 : data_mask = 256'h0000000000000000000020000000000000000000000000000000000000000000 ; 
      10'b1110010100 : data_mask = 256'h0000000000000000000040000000000000000000000000000000000000000000 ; 
      10'b0000010110 : data_mask = 256'h0000000000000000000080000000000000000000000000000000000000000000 ;
      10'b0000011001 : data_mask = 256'h0000000000000000000100000000000000000000000000000000000000000000 ; 
      10'b1011000000 : data_mask = 256'h0000000000000000000200000000000000000000000000000000000000000000 ; 
      10'b1100100000 : data_mask = 256'h0000000000000000000400000000000000000000000000000000000000000000 ; 
      10'b0001001111 : data_mask = 256'h0000000000000000000800000000000000000000000000000000000000000000 ;
      10'b0001110000 : data_mask = 256'h0000000000000000001000000000000000000000000000000000000000000000 ; 
      10'b0011000001 : data_mask = 256'h0000000000000000002000000000000000000000000000000000000000000000 ; 
      10'b0110000010 : data_mask = 256'h0000000000000000004000000000000000000000000000000000000000000000 ; 
      10'b1100000100 : data_mask = 256'h0000000000000000008000000000000000000000000000000000000000000000 ;
      10'b1000101000 : data_mask = 256'h0000000000000000010000000000000000000000000000000000000000000000 ; 
      10'b0010110000 : data_mask = 256'h0000000000000000020000000000000000000000000000000000000000000000 ; 
      10'b0101000001 : data_mask = 256'h0000000000000000040000000000000000000000000000000000000000000000 ; 
      10'b1010000010 : data_mask = 256'h0000000000000000080000000000000000000000000000000000000000000000 ;
      10'b0100100100 : data_mask = 256'h0000000000000000100000000000000000000000000000000000000000000000 ; 
      10'b1001001000 : data_mask = 256'h0000000000000000200000000000000000000000000000000000000000000000 ; 
      10'b1000000011 : data_mask = 256'h0000000000000000400000000000000000000000000000000000000000000000 ; 
      10'b0000100110 : data_mask = 256'h0000000000000000800000000000000000000000000000000000000000000000 ;
      10'b0001001100 : data_mask = 256'h0000000000000001000000000000000000000000000000000000000000000000 ; 
      10'b0010011000 : data_mask = 256'h0000000000000002000000000000000000000000000000000000000000000000 ; 
      10'b0100010001 : data_mask = 256'h0000000000000004000000000000000000000000000000000000000000000000 ; 
      10'b1000000101 : data_mask = 256'h0000000000000008000000000000000000000000000000000000000000000000 ;
      10'b0000101010 : data_mask = 256'h0000000000000010000000000000000000000000000000000000000000000000 ; 
      10'b0001010100 : data_mask = 256'h0000000000000020000000000000000000000000000000000000000000000000 ; 
      10'b0010001001 : data_mask = 256'h0000000000000040000000000000000000000000000000000000000000000000 ; 
      10'b0100010010 : data_mask = 256'h0000000000000080000000000000000000000000000000000000000000000000 ;
      10'b1000100111 : data_mask = 256'h0000000000000100000000000000000000000000000000000000000000000000 ; 
      10'b0001101011 : data_mask = 256'h0000000000000200000000000000000000000000000000000000000000000000 ; 
      10'b0011010011 : data_mask = 256'h0000000000000400000000000000000000000000000000000000000000000000 ; 
      10'b0110001101 : data_mask = 256'h0000000000000800000000000000000000000000000000000000000000000000 ;
      10'b1100010101 : data_mask = 256'h0000000000001000000000000000000000000000000000000000000000000000 ; 
      10'b1001011001 : data_mask = 256'h0000000000002000000000000000000000000000000000000000000000000000 ; 
      10'b0010101110 : data_mask = 256'h0000000000004000000000000000000000000000000000000000000000000000 ; 
      10'b0101010110 : data_mask = 256'h0000000000008000000000000000000000000000000000000000000000000000 ;
      10'b1010011010 : data_mask = 256'h0000000000010000000000000000000000000000000000000000000000000000 ; 
      10'b0100111100 : data_mask = 256'h0000000000020000000000000000000000000000000000000000000000000000 ; 
      10'b0011110001 : data_mask = 256'h0000000000040000000000000000000000000000000000000000000000000000 ; 
      10'b0101100011 : data_mask = 256'h0000000000080000000000000000000000000000000000000000000000000000 ;
      10'b1001100110 : data_mask = 256'h0000000000100000000000000000000000000000000000000000000000000000 ; 
      10'b0110101100 : data_mask = 256'h0000000000200000000000000000000000000000000000000000000000000000 ; 
      10'b1010111000 : data_mask = 256'h0000000000400000000000000000000000000000000000000000000000000000 ; 
      10'b1100110010 : data_mask = 256'h0000000000800000000000000000000000000000000000000000000000000000 ;
      10'b0111000101 : data_mask = 256'h0000000001000000000000000000000000000000000000000000000000000000 ; 
      10'b1011001010 : data_mask = 256'h0000000002000000000000000000000000000000000000000000000000000000 ; 
      10'b1101010100 : data_mask = 256'h0000000004000000000000000000000000000000000000000000000000000000 ; 
      10'b1110001001 : data_mask = 256'h0000000008000000000000000000000000000000000000000000000000000000 ;
      10'b0000010101 : data_mask = 256'h0000000010000000000000000000000000000000000000000000000000000000 ; 
      10'b0000001110 : data_mask = 256'h0000000020000000000000000000000000000000000000000000000000000000 ; 
      10'b1010100000 : data_mask = 256'h0000000040000000000000000000000000000000000000000000000000000000 ; 
      10'b0111000000 : data_mask = 256'h0000000080000000000000000000000000000000000000000000000000000000 ;
      10'b0100011011 : data_mask = 256'h0000000100000000000000000000000000000000000000000000000000000000 ; 
      10'b0111100001 : data_mask = 256'h0000000200000000000000000000000000000000000000000000000000000000 ; 
      10'b0111100100 : data_mask = 256'h0000000400000000000000000000000000000000000000000000000000000000 ; 
      10'b0111101000 : data_mask = 256'h0000000800000000000000000000000000000000000000000000000000000000 ;
      10'b0111110000 : data_mask = 256'h0000001000000000000000000000000000000000000000000000000000000000 ; 
      10'b1011100001 : data_mask = 256'h0000002000000000000000000000000000000000000000000000000000000000 ; 
      10'b1011100100 : data_mask = 256'h0000004000000000000000000000000000000000000000000000000000000000 ; 
      10'b1011101000 : data_mask = 256'h0000008000000000000000000000000000000000000000000000000000000000 ;
      10'b1101100001 : data_mask = 256'h0000010000000000000000000000000000000000000000000000000000000000 ; 
      10'b1101100010 : data_mask = 256'h0000020000000000000000000000000000000000000000000000000000000000 ; 
      10'b1101100100 : data_mask = 256'h0000040000000000000000000000000000000000000000000000000000000000 ; 
      10'b1101110000 : data_mask = 256'h0000080000000000000000000000000000000000000000000000000000000000 ;
      10'b1110101000 : data_mask = 256'h0000100000000000000000000000000000000000000000000000000000000000 ; 
      10'b1110110000 : data_mask = 256'h0000200000000000000000000000000000000000000000000000000000000000 ; 
      10'b1111000100 : data_mask = 256'h0000400000000000000000000000000000000000000000000000000000000000 ; 
      10'b1111010000 : data_mask = 256'h0000800000000000000000000000000000000000000000000000000000000000 ;
      10'b0000101111 : data_mask = 256'h0001000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0010001111 : data_mask = 256'h0002000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0100001111 : data_mask = 256'h0004000000000000000000000000000000000000000000000000000000000000 ; 
      10'b1000001111 : data_mask = 256'h0008000000000000000000000000000000000000000000000000000000000000 ;
      10'b0000110111 : data_mask = 256'h0010000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0001010111 : data_mask = 256'h0020000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0010010111 : data_mask = 256'h0040000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0000111011 : data_mask = 256'h0080000000000000000000000000000000000000000000000000000000000000 ;
      10'b0001011011 : data_mask = 256'h0100000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0010011011 : data_mask = 256'h0200000000000000000000000000000000000000000000000000000000000000 ; 
      10'b1000011011 : data_mask = 256'h0400000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0100011101 : data_mask = 256'h0800000000000000000000000000000000000000000000000000000000000000 ;
      10'b1000011101 : data_mask = 256'h1000000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0010011110 : data_mask = 256'h2000000000000000000000000000000000000000000000000000000000000000 ; 
      10'b0100011110 : data_mask = 256'h4000000000000000000000000000000000000000000000000000000000000000 ; 
      10'b1000011110 : data_mask = 256'h8000000000000000000000000000000000000000000000000000000000000000 ;
      default        : data_mask = 256'h0000000000000000000000000000000000000000000000000000000000000000 ;
  endcase
  
/*  
  ten_bit [25:0]           h_matrix;

  assign h_matrix[000] = 10'b0001100001 ; 
  assign h_matrix[001] = 10'b0011000010 ; 
  assign h_matrix[002] = 10'b0110000100 ; 
  assign h_matrix[003] = 10'b1100001000 ;
  assign h_matrix[004] = 10'b1000110000 ; 
  assign h_matrix[005] = 10'b0010100001 ; 
  assign h_matrix[006] = 10'b0101000010 ; 
  assign h_matrix[007] = 10'b1010000100 ;
  assign h_matrix[008] = 10'b0100101000 ; 
  assign h_matrix[009] = 10'b1001010000 ; 
  assign h_matrix[010] = 10'b0000100011 ; 
  assign h_matrix[011] = 10'b0001000110 ;
  assign h_matrix[012] = 10'b0010001100 ; 
  assign h_matrix[013] = 10'b0100011000 ; 
  assign h_matrix[014] = 10'b1000010001 ; 
  assign h_matrix[015] = 10'b0000100101 ;
  assign h_matrix[016] = 10'b0001001010 ; 
  assign h_matrix[017] = 10'b0010010100 ; 
  assign h_matrix[018] = 10'b0100001001 ; 
  assign h_matrix[019] = 10'b1000010010 ;
  assign h_matrix[020] = 10'b0001100111 ; 
  assign h_matrix[021] = 10'b0011001011 ; 
  assign h_matrix[022] = 10'b0110010011 ; 
  assign h_matrix[023] = 10'b1100001101 ;
  assign h_matrix[024] = 10'b1000110101 ; 
  assign h_matrix[025] = 10'b0010111001 ; 
  assign h_matrix[026] = 10'b0101001110 ; 
  assign h_matrix[027] = 10'b1010010110 ;
  assign h_matrix[028] = 10'b0100111010 ; 
  assign h_matrix[029] = 10'b1001011100 ; 
  assign h_matrix[030] = 10'b0011100011 ; 
  assign h_matrix[031] = 10'b0101100110 ;
  assign h_matrix[032] = 10'b1001101100 ; 
  assign h_matrix[033] = 10'b0110111000 ; 
  assign h_matrix[034] = 10'b1010110001 ; 
  assign h_matrix[035] = 10'b1100100101 ;
  assign h_matrix[036] = 10'b0111001010 ; 
  assign h_matrix[037] = 10'b1011010100 ; 
  assign h_matrix[038] = 10'b1101001001 ; 
  assign h_matrix[039] = 10'b1110010010 ;
  assign h_matrix[040] = 10'b0000001101 ; 
  assign h_matrix[041] = 10'b0000010011 ; 
  assign h_matrix[042] = 10'b0110100000 ; 
  assign h_matrix[043] = 10'b1001100000 ;
  assign h_matrix[044] = 10'b1111000010 ; 
  assign h_matrix[045] = 10'b0001100010 ; 
  assign h_matrix[046] = 10'b0011000100 ; 
  assign h_matrix[047] = 10'b0110001000 ;
  assign h_matrix[048] = 10'b1100010000 ; 
  assign h_matrix[049] = 10'b1000100001 ; 
  assign h_matrix[050] = 10'b0010100010 ; 
  assign h_matrix[051] = 10'b0101000100 ;
  assign h_matrix[052] = 10'b1010001000 ; 
  assign h_matrix[053] = 10'b0100110000 ; 
  assign h_matrix[054] = 10'b1001000001 ; 
  assign h_matrix[055] = 10'b0001000011 ;
  assign h_matrix[056] = 10'b0010000110 ; 
  assign h_matrix[057] = 10'b0100001100 ; 
  assign h_matrix[058] = 10'b1000011000 ; 
  assign h_matrix[059] = 10'b0000110001 ;
  assign h_matrix[060] = 10'b0001000101 ; 
  assign h_matrix[061] = 10'b0010001010 ; 
  assign h_matrix[062] = 10'b0100010100 ; 
  assign h_matrix[063] = 10'b1000001001 ;
  assign h_matrix[064] = 10'b0000110010 ; 
  assign h_matrix[065] = 10'b0011000111 ; 
  assign h_matrix[060] = 10'b0110001011 ; 
  assign h_matrix[067] = 10'b1100010011 ;
  assign h_matrix[068] = 10'b1000101101 ; 
  assign h_matrix[069] = 10'b0001110101 ; 
  assign h_matrix[070] = 10'b0101011001 ; 
  assign h_matrix[071] = 10'b1010001110 ;
  assign h_matrix[072] = 10'b0100110110 ; 
  assign h_matrix[073] = 10'b1001011010 ; 
  assign h_matrix[074] = 10'b0010111100 ; 
  assign h_matrix[075] = 10'b0011100110 ;
  assign h_matrix[076] = 10'b0101101100 ; 
  assign h_matrix[077] = 10'b1001111000 ; 
  assign h_matrix[078] = 10'b0110110001 ; 
  assign h_matrix[079] = 10'b1010100011 ;
  assign h_matrix[080] = 10'b1100101010 ; 
  assign h_matrix[081] = 10'b0111010100 ; 
  assign h_matrix[082] = 10'b1011001001 ; 
  assign h_matrix[083] = 10'b1101010010 ;
  assign h_matrix[084] = 10'b1110000101 ; 
  assign h_matrix[085] = 10'b0000001011 ; 
  assign h_matrix[086] = 10'b0000011100 ; 
  assign h_matrix[087] = 10'b0101100000 ;
  assign h_matrix[088] = 10'b1110000000 ;
  assign h_matrix[089] = 10'b1011110000 ; 
  assign h_matrix[090] = 10'b0001100100 ; 
  assign h_matrix[091] = 10'b0011001000 ;
  assign h_matrix[092] = 10'b0110010000 ; 
  assign h_matrix[093] = 10'b1100000001 ; 
  assign h_matrix[094] = 10'b1000100010 ; 
  assign h_matrix[095] = 10'b0010100100 ;
  assign h_matrix[096] = 10'b0101001000 ; 
  assign h_matrix[097] = 10'b1010010000 ; 
  assign h_matrix[098] = 10'b0100100001 ; 
  assign h_matrix[099] = 10'b1001000010 ;
  assign h_matrix[100] = 10'b0010000011 ; 
  assign h_matrix[101] = 10'b0100000110 ; 
  assign h_matrix[102] = 10'b1000001100 ; 
  assign h_matrix[103] = 10'b0000111000 ;
  assign h_matrix[104] = 10'b0001010001 ; 
  assign h_matrix[105] = 10'b0010000101 ; 
  assign h_matrix[106] = 10'b0100001010 ; 
  assign h_matrix[107] = 10'b1000010100 ;
  assign h_matrix[108] = 10'b0000101001 ; 
  assign h_matrix[109] = 10'b0001010010 ; 
  assign h_matrix[110] = 10'b0110000111 ; 
  assign h_matrix[111] = 10'b1100001011 ;
  assign h_matrix[112] = 10'b1000110011 ; 
  assign h_matrix[113] = 10'b0001101101 ; 
  assign h_matrix[114] = 10'b0011010101 ; 
  assign h_matrix[115] = 10'b1010011001 ;
  assign h_matrix[116] = 10'b0100101110 ; 
  assign h_matrix[117] = 10'b1001010110 ; 
  assign h_matrix[118] = 10'b0010111010 ; 
  assign h_matrix[119] = 10'b0101011100 ;
  assign h_matrix[120] = 10'b0011101100 ; 
  assign h_matrix[121] = 10'b0101111000 ; 
  assign h_matrix[122] = 10'b1001110001 ; 
  assign h_matrix[123] = 10'b0110100011 ;
  assign h_matrix[124] = 10'b1010100110 ; 
  assign h_matrix[125] = 10'b1100110100 ; 
  assign h_matrix[126] = 10'b0111001001 ; 
  assign h_matrix[127] = 10'b1011010010 ;
  assign h_matrix[128] = 10'b1101000101 ; 
  assign h_matrix[129] = 10'b1110001010 ; 
  assign h_matrix[130] = 10'b0000011010 ; 
  assign h_matrix[131] = 10'b0000000111 ;
  assign h_matrix[132] = 10'b1101000000 ; 
  assign h_matrix[133] = 10'b0011100000 ; 
  assign h_matrix[134] = 10'b1110100100 ; 
  assign h_matrix[135] = 10'b0001101000 ;
  assign h_matrix[136] = 10'b0011010000 ; 
  assign h_matrix[137] = 10'b0110000001 ; 
  assign h_matrix[138] = 10'b1100000010 ; 
  assign h_matrix[139] = 10'b1000100100 ;
  assign h_matrix[140] = 10'b0010101000 ; 
  assign h_matrix[141] = 10'b0101010000 ; 
  assign h_matrix[142] = 10'b1010000001 ; 
  assign h_matrix[143] = 10'b0100100010 ;
  assign h_matrix[144] = 10'b1001000100 ; 
  assign h_matrix[145] = 10'b0100000011 ; 
  assign h_matrix[146] = 10'b1000000110 ; 
  assign h_matrix[147] = 10'b0000101100 ;
  assign h_matrix[148] = 10'b0001011000 ; 
  assign h_matrix[149] = 10'b0010010001 ; 
  assign h_matrix[150] = 10'b0100000101 ; 
  assign h_matrix[151] = 10'b1000001010 ;
  assign h_matrix[152] = 10'b0000110100 ; 
  assign h_matrix[153] = 10'b0001001001 ; 
  assign h_matrix[154] = 10'b0010010010 ; 
  assign h_matrix[155] = 10'b1100000111 ;
  assign h_matrix[156] = 10'b1000101011 ; 
  assign h_matrix[157] = 10'b0001110011 ; 
  assign h_matrix[158] = 10'b0011001101 ; 
  assign h_matrix[159] = 10'b0110010101 ;
  assign h_matrix[160] = 10'b0100111001 ; 
  assign h_matrix[161] = 10'b1001001110 ; 
  assign h_matrix[162] = 10'b0010110110 ; 
  assign h_matrix[163] = 10'b0101011010 ;
  assign h_matrix[164] = 10'b1010011100 ; 
  assign h_matrix[165] = 10'b0011111000 ; 
  assign h_matrix[166] = 10'b0101110001 ; 
  assign h_matrix[167] = 10'b1001100011 ;
  assign h_matrix[168] = 10'b0110100110 ; 
  assign h_matrix[169] = 10'b1010101100 ; 
  assign h_matrix[170] = 10'b1100101001 ; 
  assign h_matrix[171] = 10'b0111010010 ;
  assign h_matrix[172] = 10'b1011000101 ; 
  assign h_matrix[173] = 10'b1101001010 ; 
  assign h_matrix[174] = 10'b1110010100 ; 
  assign h_matrix[175] = 10'b0000010110 ;
  assign h_matrix[176] = 10'b0000011001 ; 
  assign h_matrix[177] = 10'b1011000000 ; 
  assign h_matrix[178] = 10'b1100100000 ; 
  assign h_matrix[179] = 10'b0001001111 ;
  assign h_matrix[180] = 10'b0001110000 ; 
  assign h_matrix[181] = 10'b0011000001 ; 
  assign h_matrix[182] = 10'b0110000010 ; 
  assign h_matrix[183] = 10'b1100000100 ;
  assign h_matrix[184] = 10'b1000101000 ; 
  assign h_matrix[185] = 10'b0010110000 ; 
  assign h_matrix[186] = 10'b0101000001 ; 
  assign h_matrix[187] = 10'b1010000010 ;
  assign h_matrix[188] = 10'b0100100100 ; 
  assign h_matrix[189] = 10'b1001001000 ; 
  assign h_matrix[190] = 10'b1000000011 ; 
  assign h_matrix[191] = 10'b0000100110 ;
  assign h_matrix[192] = 10'b0001001100 ; 
  assign h_matrix[193] = 10'b0010011000 ; 
  assign h_matrix[194] = 10'b0100010001 ; 
  assign h_matrix[195] = 10'b1000000101 ;
  assign h_matrix[196] = 10'b0000101010 ; 
  assign h_matrix[197] = 10'b0001010100 ; 
  assign h_matrix[198] = 10'b0010001001 ; 
  assign h_matrix[199] = 10'b0100010010 ;
  assign h_matrix[200] = 10'b1000100111 ; 
  assign h_matrix[201] = 10'b0001101011 ; 
  assign h_matrix[202] = 10'b0011010011 ; 
  assign h_matrix[203] = 10'b0110001101 ;
  assign h_matrix[204] = 10'b1100010101 ; 
  assign h_matrix[205] = 10'b1001011001 ; 
  assign h_matrix[206] = 10'b0010101110 ; 
  assign h_matrix[207] = 10'b0101010110 ;
  assign h_matrix[208] = 10'b1010011010 ; 
  assign h_matrix[209] = 10'b0100111100 ; 
  assign h_matrix[210] = 10'b0011110001 ; 
  assign h_matrix[211] = 10'b0101100011 ;
  assign h_matrix[212] = 10'b1001100110 ; 
  assign h_matrix[213] = 10'b0110101100 ; 
  assign h_matrix[214] = 10'b1010111000 ; 
  assign h_matrix[215] = 10'b1100110010 ;
  assign h_matrix[216] = 10'b0111000101 ; 
  assign h_matrix[217] = 10'b1011001010 ; 
  assign h_matrix[218] = 10'b1101010100 ; 
  assign h_matrix[219] = 10'b1110001001 ;
  assign h_matrix[220] = 10'b0000010101 ; 
  assign h_matrix[221] = 10'b0000001110 ; 
  assign h_matrix[222] = 10'b1010100000 ; 
  assign h_matrix[223] = 10'b0111000000 ;
  assign h_matrix[224] = 10'b0100011011 ; 
  assign h_matrix[225] = 10'b0111100001 ; 
  assign h_matrix[226] = 10'b0111100100 ; 
  assign h_matrix[227] = 10'b0111101000 ;
  assign h_matrix[228] = 10'b0111110000 ; 
  assign h_matrix[229] = 10'b1011100001 ; 
  assign h_matrix[230] = 10'b1011100100 ; 
  assign h_matrix[231] = 10'b1011101000 ;
  assign h_matrix[232] = 10'b1101100001 ; 
  assign h_matrix[233] = 10'b1101100010 ; 
  assign h_matrix[234] = 10'b1101100100 ; 
  assign h_matrix[235] = 10'b1101110000 ;
  assign h_matrix[236] = 10'b1110101000 ; 
  assign h_matrix[237] = 10'b1110110000 ; 
  assign h_matrix[238] = 10'b1111000100 ; 
  assign h_matrix[239] = 10'b1111010000 ;
  assign h_matrix[240] = 10'b0000101111 ; 
  assign h_matrix[241] = 10'b0010001111 ; 
  assign h_matrix[242] = 10'b0100001111 ; 
  assign h_matrix[243] = 10'b1000001111 ;
  assign h_matrix[244] = 10'b0000110111 ; 
  assign h_matrix[245] = 10'b0001010111 ; 
  assign h_matrix[246] = 10'b0010010111 ; 
  assign h_matrix[247] = 10'b0000111011 ;
  assign h_matrix[248] = 10'b0001011011 ; 
  assign h_matrix[249] = 10'b0010011011 ; 
  assign h_matrix[250] = 10'b1000011011 ; 
  assign h_matrix[251] = 10'b0100011101 ;
  assign h_matrix[252] = 10'b1000011101 ; 
  assign h_matrix[253] = 10'b0010011110 ; 
  assign h_matrix[254] = 10'b0100011110 ; 
  assign h_matrix[255] = 10'b1000011110 ;
*/
/*
/////////////////////////////////////////////////////////////////////////////////////////////// 
//IS this the same??
  logic         bit0 ;
  logic         bit1 ;
  logic         bit2 ;
  logic         bit3 ;
  logic         bit4 ;
  logic         bit5 ;
  logic         bit6 ;
  logic         bit7 ;
  logic         bit8 ;
  logic         bit9 ;
  logic [9:0]   chk2 ;
  logic [9:0]   synd ;
  logic [3:0]   sum;
  logic         sbe_x;
  logic         mbe_x;
  
  logic [255:0] data_out_x ;
  
  logic [255:0] vecx0  ;
  logic [255:0] vecx1  ;
  logic [255:0] vecx2  ;    
  logic [255:0] vecx3  ;
  logic [255:0] vecx4  ;
  logic [255:0] vecx5  ;
  logic [255:0] vecx6  ;
  logic [255:0] vecx7  ;
  logic [255:0] vecx8  ;
  logic [255:0] vecx9  ; 
  
  logic [255:0] zero ;
  
  logic [255:0] vec0  ;
  logic [255:0] vec1  ;
  logic [255:0] vec2  ;    
  logic [255:0] vec3  ;
  logic [255:0] vec4  ;
  logic [255:0] vec5  ;
  logic [255:0] vec6  ;
  logic [255:0] vec7  ;
  logic [255:0] vec8  ;
  logic [255:0] vec9  ; 
  
    assign zero  =  256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
  
    assign vecx0 =  256'h1fff0123190c3f4c442914c1fa6242094c0fd3142034c07d98c2034c43f4c421;
    assign vecx1 =  256'he7ff02012299c790c848a98e3c86840e9871e43840298b8f21843290dc790c42;
    assign vecx2 =  256'hf87f44443532d9299088d316c94d084931b64a6084521db253084129ad929884;
    assign vecx3 =  256'hff8f10892a636a532109263b5298108643da94c1086536d4a610815336a53108;
    assign vecx4 =  256'hfff0a81114c7b4a60211c87da5302104a6ed2982124a67694c2102a63b4a6210;
    assign vecx5 =  256'h00913ffe40fe4310931407e5310898e03f531084c681fd3108262c0fd3108531;
    assign vecx6 =  256'h0120cffe871ca621243a38ea621121b1c7a621090e8e3a6210c87871e4310a43;
    assign vecx7 =  256'h2242f0fecb654c420a625b34c4205362d94c42129b16cc862114d4b64a6210a6;
    assign vecx8 =  256'h4804ff1f8daa988414c46d498842a6536a90c425319b514c422994da94c4214c;
    assign vecx9 =  256'h9408ffe04ed131086986769218854c53b429884a631da298845318ed29884298;
    
  fxr_10b_ecc_gen fxr_10b_ecc_gen0(
     .data  (data_in),  
     .chk   (chk2)
  );
   
    assign synd = chk_in ^ chk2 ;
  
    assign syn = synd ;
  
    assign sum = {3'b0,synd[0]} + {3'b0,synd[1]} + {3'b0,synd[2]} + {3'b0,synd[3]} + {3'b0,synd[4]} +
               {3'b0,synd[5]} + {3'b0,synd[6]} + {3'b0,synd[7]} + {3'b0,synd[8]} + {3'b0,synd[9]} ; 
  
//  always_comb begin 
//    if(synd == 10'h0) begin
//      sbe_x = 1'b0 ;
//      mbe_x = 1'b0 ;
//    end  
//    else if((sum == 4'h1) | (sum == 4'h3)  | (sum == 4'h4) | (sum == 4'h5)) begin   //??
//      sbe_x = 1'b1 ;
//      mbe_x = 1'b0 ;
//    end
//    else begin
//      sbe_x = 1'b0 ;
//      mbe_x = 1'b1 ;
//    end 
//  end  
  
//    assign sbe = sbe_x ;
  
//    assign mbe = mbe_x ;
  
//  always_comb begin 
//    if(sum == 4'h1)
//      chk_out = chk2 ;
//    else
//      chk_out = chk_in ;
//  end 
  
    assign vec0 = (synd[0] == 1'b1) ? vecx0 : zero ;
    assign vec1 = (synd[1] == 1'b1) ? vecx1 : zero ;
    assign vec2 = (synd[2] == 1'b1) ? vecx2 : zero ;
    assign vec3 = (synd[3] == 1'b1) ? vecx3 : zero ;
    assign vec4 = (synd[4] == 1'b1) ? vecx4 : zero ;
    assign vec5 = (synd[5] == 1'b1) ? vecx5 : zero ;
    assign vec6 = (synd[6] == 1'b1) ? vecx6 : zero ;
    assign vec7 = (synd[7] == 1'b1) ? vecx7 : zero ;
    assign vec8 = (synd[8] == 1'b1) ? vecx8 : zero ;
    assign vec9 = (synd[9] == 1'b1) ? vecx9 : zero ;
  
//                     (SBE on check bit)       (SBE in data)
    assign data_out_x = (sum == 4'h1) ? data_in : (vec0 & vec1 & vec2 & vec3 & vec4 & vec5 & vec6 & vec7 & vec8 & vec9) ^ data_in ;
  
//    assign   data_out = data_out_x ;
//    assign data_out = data_in ;
*/        

/*  
  logic [255:0] vec0  ;
  logic [255:0] vec1  ;
  logic [255:0] vec2  ;    
  logic [255:0] vec3  ;
  logic [255:0] vec4  ;
  logic [255:0] vec5  ;
  logic [255:0] vec6  ;
  logic [255:0] vec7  ;
  logic [255:0] vec8  ;
  logic [255:0] vec9  ;  
  
    assign vec0 = (2**0)+(2**5)+(2**10)+(2**14)+(2**15)+(2**18)+(2**20)+(2**21)+(2**22)+(2**23)+(2**24)+(2**25)+(2**30)+(2**34)+(2**35)+(2**38)+(2**40)+(2**41)+(2**49)+(2**54)+(2**55)+(2**59)+(2**60)+(2**63)+(2**64)+(2**66)+(2**67)+(2**68)+(2**69)+(2**70)+(2**78)+(2**79)+(2**82)+(2**84)+(2**85)+(2**93)+(2**98)+(2**100)+(2**104)+(2**105)+(2**108)+(2**110)+(2**111)+(2**112)+(2**113)+(2**114)+(2**115)+(2**122)+(2**123)+(2**126)+(2**128)+(2**131)+(2**137)+(2**142)+(2**145)+(2**149)+(2**150)+(2**153)+(2**155)+(2**156)+(2**157)+(2**158)+(2**159)+(2**160)+(2**166)+(2**167)+(2**170)+(2**172)+(2**176)+(2**179)+(2**181)+(2**186)+(2**190)+(2**194)+(2**195)+(2**198)+(2**200)+(2**201)+(2**202)+(2**203)+(2**204)+(2**205)+(2**210)+(2**211)+(2**216)+(2**219)+(2**220)+(2**224)+(2**225)+(2**229)+(2**232)+(2**240)+(2**241)+(2**242)+(2**243)+(2**244)+(2**245)+(2**246)+(2**247)+(2**248)+(2**249)+(2**250)+(2**251)+(2**252);
    assign vec1 = (2**1)+(2**6)+(2**10)+(2**11)+(2**16)+(2**19)+(2**20)+(2**21)+(2**22)+(2**26)+(2**27)+(2**28)+(2**30)+(2**31)+(2**36)+(2**39)+(2**41)+(2**44)+(2**45)+(2**50)+(2**55)+(2**56)+(2**61)+(2**64)+(2**65)+(2**66)+(2**67)+(2**71)+(2**72)+(2**73)+(2**75)+(2**79)+(2**80)+(2**83)+(2**85)+(2**94)+(2**99)+(2**100)+(2**101)+(2**106)+(2**109)+(2**110)+(2**111)+(2**112)+(2**116)+(2**117)+(2**118)+(2**123)+(2**124)+(2**127)+(2**129)+(2**130)+(2**131)+(2**138)+(2**143)+(2**145)+(2**146)+(2**151)+(2**154)+(2**155)+(2**156)+(2**157)+(2**161)+(2**162)+(2**163)+(2**167)+(2**168)+(2**171)+(2**173)+(2**175)+(2**179)+(2**182)+(2**187)+(2**190)+(2**191)+(2**196)+(2**199)+(2**200)+(2**201)+(2**202)+(2**206)+(2**207)+(2**208)+(2**211)+(2**212)+(2**215)+(2**217)+(2**221)+(2**224)+(2**233)+(2**240)+(2**241)+(2**242)+(2**243)+(2**244)+(2**245)+(2**246)+(2**247)+(2**248)+(2**249)+(2**250)+(2** 253)+(2**254)+(2**255);
    assign vec2 = (2**2)+(2**7)+(2**11)+(2**12)+(2**15)+(2**17)+(2**20)+(2**23)+(2**24)+(2**26)+(2**27)+(2**29)+(2**31)+(2**32)+(2**35)+(2**37)+(2**40)+(2**46)+(2**51)+(2**56)+(2**57)+(2**60)+(2**62)+(2**65)+(2**68)+(2**69)+(2**71)+(2**72)+(2**74)+(2**75)+(2**76)+(2**81)+(2**84)+(2**86)+(2**90)+(2**95)+(2**101)+(2**102)+(2**105)+(2**107)+(2**110)+(2**113)+(2**114)+(2**116)+(2**117)+(2**119)+(2**120)+(2**124)+(2**125)+(2**128)+(2**131)+(2**134)+(2**139)+(2**144)+(2**146)+(2**147)+(2**150)+(2**152)+(2**155)+(2**158)+(2**159)+(2**161)+(2**162)+(2**164)+(2**168)+(2**169)+(2**172)+(2**174)+(2**175)+(2**179)+(2**183)+(2**188)+(2**191)+(2**192)+(2**195)+(2**197)+(2**200)+(2**203)+(2**204)+(2**206)+(2**207)+(2**209)+(2**212)+(2**213)+(2**216)+(2**218)+(2**220)+(2**221)+(2**226)+(2**230)+(2**234)+(2**238)+(2**240)+(2**241)+(2**242)+(2**243)+(2**244)+(2**245)+(2**246)+(2**251)+(2**252)+(2**253)+(2**254)+(2**255);
    assign vec3 = (2**3)+(2**8)+(2**12)+(2**13)+(2**16)+(2**18)+(2**21)+(2**23)+(2**25)+(2**26)+(2**28)+(2**29)+(2**32)+(2**33)+(2**36)+(2**38)+(2**40)+(2**47)+(2**52)+(2**57)+(2**58)+(2**61)+(2**63)+(2** 66)+(2**68)+(2**70)+(2**71)+(2**73)+(2**74)+(2**76)+(2**77)+(2**80)+(2**82)+(2**85)+(2**86)+(2**91)+(2**96)+(2**102)+(2**103)+(2**106)+(2**108)+(2**111)+(2**113)+(2**115)+(2**116)+(2**118)+(2**119)+(2**120)+(2**121)+(2**126)+(2**129)+(2**130)+(2**135)+(2**140)+(2**147)+(2**148)+(2**151)+(2**153)+(2**156)+(2**158)+(2**160)+(2**161)+(2**163)+(2**164)+(2**165)+(2**169)+(2**170)+(2**173)+(2**176)+(2**179)+(2**184)+(2**189)+(2**192)+(2**193)+(2**196)+(2**198)+(2**201)+(2**203)+(2**205)+(2**206)+(2**208)+(2**209)+(2**213)+(2**214)+(2**217)+(2**219)+(2**221)+(2**224)+(2**227)+(2**231)+(2**236)+(2**240)+(2**241)+(2**242)+(2**243)+(2**247)+(2**248)+(2**249)+(2**250)+(2**251)+(2**252)+(2**253)+(2**254)+(2**255);
    assign vec4 = (2**4)+(2**9)+(2**13)+(2**14)+(2**17)+(2**19)+(2**22)+(2**24)+(2**25)+(2**27)+(2**28)+(2**29)+(2**33)+(2**34)+(2**37)+(2**39)+(2**41)+(2**48)+(2**53)+(2**58)+(2**59)+(2**62)+(2**64)+(2**67)+(2**69)+(2**70)+(2**72)+(2**73)+(2**74)+(2**77)+(2**78)+(2**81)+(2**83)+(2**86)+(2**89)+(2**92)+(2**97)+(2**103)+(2**104)+(2**107)+(2**109)+(2**112)+(2**114)+(2**115)+(2**117)+(2**118)+(2**119)+(2**121)+(2**122)+(2**125)+(2**127)+(2**130)+(2**136)+(2**141)+(2**148)+(2**149)+(2**152)+(2**154)+(2**157)+(2**159)+(2**160)+(2**162)+(2**163)+(2**164)+(2**165)+(2**166)+(2**171)+(2**174)+(2**175)+(2**176)+(2**180)+(2**185)+(2**193)+(2**194)+(2**197)+(2**199)+(2**202)+(2**204)+(2**205)+(2**207)+(2**208)+(2**209)+(2**210)+(2**214)+(2**215)+(2**218)+(2**220)+(2**224)+(2**228)+(2**235)+(2**237)+(2**239)+(2**244)+(2**245)+(2**246)+(2**247)+(2**248)+(2**249)+(2**250)+(2**251)+(2**252)+(2**253)+(2**254)+(2**255);
    assign vec5 = (2**0)+(2**4)+(2**5)+(2**8)+(2**10)+(2**15)+(2**20)+(2**24)+(2**25)+(2**28)+(2**30)+(2**31)+(2**32)+(2**33)+(2**34)+(2**35)+(2**42)+(2**43)+(2**45)+(2**49)+(2**50)+(2**53)+(2**59)+(2**64)+(2**68)+(2**69)+(2**72)+(2**74)+(2**75)+(2**76)+(2**77)+(2**78)+(2**79)+(2**80)+(2**87)+(2**89)+(2**90)+(2**94)+(2**95)+(2**98)+(2**103)+(2**108)+(2**112)+(2**113)+(2**116)+(2**118)+(2**120)+(2**121)+(2**122)+(2**123)+(2**124)+(2**125)+(2**133)+(2**134)+(2**135)+(2**139)+(2**140)+(2**143)+(2**147)+(2**152)+(2**156)+(2**157)+(2**160)+(2**162)+(2**165)+(2**166)+(2**167)+(2**168)+(2**169)+(2**170)+(2**178)+(2**180)+(2**184)+(2**185)+(2**188)+(2**191)+(2**196)+(2**200)+(2**201)+(2**206)+(2**209)+(2**210)+(2**211)+(2**212)+(2**213)+(2**214)+(2**215)+(2**222)+(2**225)+(2**226)+(2**227)+(2**228)+(2**229)+(2**230)+(2**231)+(2**232)+(2**233)+(2**234)+(2**235)+(2**236)+(2**237)+(2**240)+(2**244)+(2**247);
    assign vec6 = (2**0)+(2**1)+(2**6)+(2**9)+(2**11)+(2**16)+(2**20)+(2**21)+(2**26)+(2**29)+(2**30)+(2**31)+(2**32)+(2**36)+(2**37)+(2**38)+(2**43)+(2**44)+(2**45)+(2**46)+(2**51)+(2**54)+(2**55)+(2**60)+(2**65)+(2**69)+(2**70)+(2**73)+(2**75)+(2**76)+(2**77)+(2**81)+(2**82)+(2**83)+(2**87)+(2**89)+(2**90)+(2**91)+(2**96)+(2**99)+(2**104)+(2**109)+(2**113)+(2**114)+(2**117)+(2**119)+(2**120)+(2**121)+(2**122)+(2**126)+(2**127)+(2**128)+(2**132)+(2**133)+(2**135)+(2**136)+(2**141)+(2**144)+(2**148)+(2**153)+(2**157)+(2**158)+(2**161)+(2**163)+(2**165)+(2**166)+(2**167)+(2**171)+(2**172)+(2**173)+(2**177)+(2**179)+(2**180)+(2**181)+(2**186)+(2**189)+(2**192)+(2**197)+(2**201)+(2**202)+(2**205)+(2**207)+(2**210)+(2**211)+(2**212)+(2**216)+(2**217)+(2**218)+(2**223)+(2**225)+(2**226)+(2**227)+(2**228)+(2**229)+(2**230)+(2**231)+(2**232)+(2**233)+(2**234)+(2**235)+(2**238)+(2**239)+(2**245)+(2**248);
    assign vec7 = (2**1)+(2**2)+(2**5)+(2**7)+(2**12)+(2**17)+(2**21)+(2**22)+(2**25)+(2**27)+(2**30)+(2**33)+(2**34)+(2**36)+(2**37)+(2**39)+(2**42)+(2**44)+(2**46)+(2**47)+(2**50)+(2**52)+(2**56)+(2**61)+(2**65)+(2**66)+(2**71)+(2**74)+(2**75)+(2**78)+(2**79)+(2**81)+(2**82)+(2**84)+(2**88)+(2**89)+(2**91)+(2**92)+(2**95)+(2**97)+(2**100)+(2**105)+(2**110)+(2**114)+(2**115)+(2**118)+(2**120)+(2**123)+(2**124)+(2**126)+(2**127)+(2**129)+(2**133)+(2**134)+(2**136)+(2**137)+(2**140)+(2**142)+(2**149)+(2**154)+(2**158)+(2**159)+(2**162)+(2**164)+(2**165)+(2**168)+(2**169)+(2**171)+(2**172)+(2**174)+(2**177)+(2**181)+(2**182)+(2**185)+(2**187)+(2**193)+(2**198)+(2**202)+(2**203)+(2**206)+(2**208)+(2**210)+(2**213)+(2**214)+(2**216)+(2**217)+(2**219)+(2**222)+(2**223)+(2**225)+(2**226)+(2**227)+(2**228)+(2**229)+(2**230)+(2**231)+(2**236)+(2**237)+(2**238)+(2**239)+(2**241)+(2**246)+(2**249)+(2**253);
    assign vec8 = (2**2)+(2**3)+(2**6)+(2**8)+(2**13)+(2**18)+(2**22)+(2**23)+(2**26)+(2**28)+(2**31)+(2**33)+(2**35)+(2**36)+(2**38)+(2**39)+(2**42)+(2**44)+(2**47)+(2**48)+(2**51)+(2**53)+(2**57)+(2**62)+(2**66)+(2**67)+(2**70)+(2**72)+(2**76)+(2**78)+(2**80)+(2**81)+(2**83)+(2**84)+(2**87)+(2**88)+(2**92)+(2**93)+(2**96)+(2**98)+(2**101)+(2**106)+(2**110)+(2**111)+(2**116)+(2**119)+(2**121)+(2**123)+(2**125)+(2**126)+(2**128)+(2**129)+(2**132)+(2**134)+(2**137)+(2**138)+(2**141)+(2**143)+(2**145)+(2**150)+(2**155)+(2**159)+(2**160)+(2**163)+(2**166)+(2**168)+(2**170)+(2**171)+(2**173)+(2**174)+(2**178)+(2**182)+(2**183)+(2**186)+(2**188)+(2**194)+(2**199)+(2**203)+(2**204)+(2**207)+(2**209)+(2**211)+(2**213)+(2**215)+(2**216)+(2**218)+(2**219)+(2**223)+(2**224)+(2**225)+(2**226)+(2**227)+(2**228)+(2**232)+(2**233)+(2**234)+(2**235)+(2**236)+(2**237)+(2**238)+(2**239)+(2**242)+(2**251)+(2**254);
    assign vec9 = (2**3)+(2**4)+(2**7)+(2**9)+(2**14)+(2**19)+(2**23)+(2**24)+(2**27)+(2**29)+(2**32)+(2**34)+(2**35)+(2**37)+(2**38)+(2**39)+(2**43)+(2**44)+(2**48)+(2**49)+(2**52)+(2**54)+(2**58)+(2**63)+(2**67)+(2**68)+(2**71)+(2**73)+(2**77)+(2**79)+(2**80)+(2**82)+(2**83)+(2**84)+(2**88)+(2**89)+(2**93)+(2**94)+(2**97)+(2**99)+(2**102)+(2**107)+(2**111)+(2**112)+(2**115)+(2**117)+(2**122)+(2**124)+(2**125)+(2**127)+(2**128)+(2**129)+(2**132)+(2**134)+(2**138)+(2**139)+(2**142)+(2**144)+(2**146)+(2**151)+(2**155)+(2**156)+(2**161)+(2**164)+(2**167)+(2**169)+(2**170)+(2**172)+(2**173)+(2**174)+(2**177)+(2**178)+(2**183)+(2**184)+(2**187)+(2**189)+(2**190)+(2**195)+(2**200)+(2**204)+(2**205)+(2**208)+(2**212)+(2**214)+(2**215)+(2**217)+(2**218)+(2**219)+(2**222)+(2**229)+(2**230)+(2**231)+(2**232)+(2**233)+(2**234)+(2**235)+(2**236)+(2**237)+(2**238)+(2**239)+(2**243)+(2**250)+(2**252)+(2**255);
  
  
  logic [255:0] vecx0  ;
  logic [255:0] vecx1  ;
  logic [255:0] vecx2  ;    
  logic [255:0] vecx3  ;
  logic [255:0] vecx4  ;
  logic [255:0] vecx5  ;
  logic [255:0] vecx6  ;
  logic [255:0] vecx7  ;
  logic [255:0] vecx8  ;
  logic [255:0] vecx9  ; 
  
    assign vecx0 =  256'h1fff0123190c3f4c442914c1fa6242094c0fd3142034c07d98c2034c43f4c421;
    assign vecx1 =  256'he7ff02012299c790c848a98e3c86840e9871e43840298b8f21843290dc790c42;
    assign vecx2 =  256'hf87f44443532d9299088d316c94d084931b64a6084521db253084129ad929884;
    assign vecx3 =  256'hff8f10892a636a532109263b5298108643da94c1086536d4a610815336a53108;
    assign vecx4 =  256'hfff0a81114c7b4a60211c87da5302104a6ed2982124a67694c2102a63b4a6210;
    assign vecx5 =  256'h00913ffe40fe4310931407e5310898e03f531084c681fd3108262c0fd3108531;
    assign vecx6 =  256'h0120cffe871ca621243a38ea621121b1c7a621090e8e3a6210c87871e4310a43;
    assign vecx7 =  256'h2242f0fecb654c420a625b34c4205362d94c42129b16cc862114d4b64a6210a6;
    assign vecx8 =  256'h4804ff1f8daa988414c46d498842a6536a90c425319b514c422994da94c4214c;
    assign vecx9 =  256'h9408ffe04ed131086986769218854c53b429884a631da298845318ed29884298 ;
  
  logic [9:0] tes;
  
    assign tes[0] = (vec0 == vecx0) ;
    assign tes[1] = (vec1 == vecx1) ;
    assign tes[2] = (vec2 == vecx2) ;
    assign tes[3] = (vec3 == vecx3) ;
    assign tes[4] = (vec4 == vecx4) ;
    assign tes[5] = (vec5 == vecx5) ;
    assign tes[6] = (vec6 == vecx6) ;
    assign tes[7] = (vec7 == vecx7) ;
    assign tes[8] = (vec8 == vecx8) ;
    assign tes[9] = (vec9 == vecx9) ;
*/
  
endmodule // fxr_10b_ecc_cor
