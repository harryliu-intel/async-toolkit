magic
tech scmos
timestamp 965070645
<< ndiffusion >>
rect 198 660 206 661
rect 198 656 206 657
rect 198 647 206 648
rect 198 643 206 644
rect 198 634 206 635
rect 198 630 206 631
rect 198 621 206 622
rect 198 617 206 618
rect 198 608 206 609
rect 198 604 206 605
rect 198 595 206 596
rect 198 591 206 592
rect 198 582 206 583
rect 198 578 206 579
rect 198 569 206 570
rect 198 565 206 566
<< pdiffusion >>
rect 222 650 230 651
rect 222 642 230 647
rect 222 638 230 639
rect 222 629 230 630
rect 222 621 230 626
rect 222 617 230 618
rect 222 608 230 609
rect 222 600 230 605
rect 222 596 230 597
rect 222 587 230 588
rect 222 579 230 584
rect 222 575 230 576
<< ntransistor >>
rect 198 657 206 660
rect 198 644 206 647
rect 198 631 206 634
rect 198 618 206 621
rect 198 605 206 608
rect 198 592 206 595
rect 198 579 206 582
rect 198 566 206 569
<< ptransistor >>
rect 222 647 230 650
rect 222 639 230 642
rect 222 626 230 629
rect 222 618 230 621
rect 222 605 230 608
rect 222 597 230 600
rect 222 584 230 587
rect 222 576 230 579
<< polysilicon >>
rect 194 657 198 660
rect 206 657 220 660
rect 217 650 220 657
rect 217 647 222 650
rect 230 647 234 650
rect 194 644 198 647
rect 206 644 211 647
rect 208 642 211 644
rect 208 639 222 642
rect 230 639 234 642
rect 194 631 198 634
rect 206 631 211 634
rect 208 629 211 631
rect 208 626 222 629
rect 230 626 234 629
rect 194 618 198 621
rect 206 618 222 621
rect 230 618 234 621
rect 194 605 198 608
rect 206 605 222 608
rect 230 605 234 608
rect 208 597 222 600
rect 230 597 234 600
rect 208 595 211 597
rect 194 592 198 595
rect 206 592 211 595
rect 208 584 222 587
rect 230 584 234 587
rect 208 582 211 584
rect 194 579 198 582
rect 206 579 211 582
rect 217 576 222 579
rect 230 576 234 579
rect 217 569 220 576
rect 194 566 198 569
rect 206 566 220 569
<< ndcontact >>
rect 198 661 206 669
rect 198 648 206 656
rect 198 635 206 643
rect 198 622 206 630
rect 198 609 206 617
rect 198 596 206 604
rect 198 583 206 591
rect 198 570 206 578
rect 198 557 206 565
<< pdcontact >>
rect 222 651 230 659
rect 222 630 230 638
rect 222 609 230 617
rect 222 588 230 596
rect 222 567 230 575
<< polycontact >>
rect 186 644 194 652
rect 234 647 242 655
rect 186 618 194 626
rect 234 626 242 634
rect 234 605 242 613
rect 186 592 194 600
rect 234 584 242 592
rect 186 566 194 574
<< metal1 >>
rect 198 661 206 669
rect 186 644 194 652
rect 198 648 218 656
rect 222 651 230 659
rect 187 626 193 644
rect 198 635 206 643
rect 210 638 218 648
rect 234 647 242 655
rect 210 630 230 638
rect 235 634 241 647
rect 186 618 194 626
rect 198 622 218 630
rect 234 626 242 634
rect 187 600 193 618
rect 198 609 206 617
rect 210 604 218 622
rect 222 609 230 617
rect 235 613 241 626
rect 234 605 242 613
rect 186 592 194 600
rect 198 596 218 604
rect 187 574 193 592
rect 198 583 206 591
rect 210 588 230 596
rect 235 592 241 605
rect 210 578 218 588
rect 234 584 242 592
rect 186 566 194 574
rect 198 570 218 578
rect 222 567 230 575
rect 198 557 206 565
<< labels >>
rlabel metal1 202 600 202 600 1 x
rlabel polysilicon 197 606 197 606 1 b
rlabel polysilicon 197 593 197 593 1 a
rlabel polysilicon 197 567 197 567 1 a
rlabel polysilicon 197 580 197 580 1 b
rlabel metal1 202 652 202 652 1 x
rlabel polysilicon 197 658 197 658 1 b
rlabel polysilicon 197 645 197 645 1 a
rlabel metal1 202 626 202 626 5 x
rlabel polysilicon 197 619 197 619 1 a
rlabel polysilicon 197 632 197 632 1 b
rlabel polysilicon 231 606 231 606 7 b
rlabel polysilicon 231 598 231 598 7 a
rlabel polysilicon 231 585 231 585 7 b
rlabel polysilicon 231 577 231 577 7 a
rlabel metal1 226 592 226 592 5 x
rlabel polysilicon 231 619 231 619 7 a
rlabel polysilicon 231 627 231 627 7 b
rlabel polysilicon 231 640 231 640 7 a
rlabel polysilicon 231 648 231 648 7 b
rlabel metal1 226 634 226 634 5 x
rlabel metal1 202 574 202 574 5 x
rlabel metal1 202 665 202 665 5 GND!
rlabel metal1 202 639 202 639 1 GND!
rlabel metal1 202 613 202 613 1 GND!
rlabel metal1 202 587 202 587 1 GND!
rlabel metal1 202 561 202 561 1 GND!
rlabel metal1 226 571 226 571 1 Vdd!
rlabel metal1 226 613 226 613 1 Vdd!
rlabel metal1 226 655 226 655 1 Vdd!
rlabel space 185 556 199 670 7 ^n
rlabel space 229 566 243 660 3 ^p
<< end >>
