magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -19 50 -15 51
rect -1 50 3 51
rect -19 44 -15 48
rect -1 44 3 48
rect -19 38 -15 42
rect -33 30 -29 35
rect -19 35 -15 36
rect -19 30 -15 31
rect -1 38 3 42
rect -1 35 3 36
rect -1 30 3 31
rect -33 25 -29 28
rect -19 24 -15 28
rect -1 24 3 28
rect -19 18 -15 22
rect -1 18 3 22
rect -19 15 -15 16
rect -1 15 3 16
<< pdiffusion >>
rect 15 44 19 45
rect 33 44 39 45
rect 48 44 60 45
rect 15 38 19 42
rect 33 38 39 42
rect 48 41 60 42
rect 48 38 56 41
rect 15 35 19 36
rect 15 30 19 31
rect 15 24 19 28
rect 33 35 39 36
rect 37 31 39 35
rect 33 30 39 31
rect 52 30 55 33
rect 33 24 39 28
rect 49 26 55 30
rect 15 21 19 22
rect 33 21 39 22
rect 49 21 55 24
<< ntransistor >>
rect -19 48 -15 50
rect -1 48 3 50
rect -19 42 -15 44
rect -1 42 3 44
rect -19 36 -15 38
rect -1 36 3 38
rect -33 28 -29 30
rect -19 28 -15 30
rect -1 28 3 30
rect -19 22 -15 24
rect -1 22 3 24
rect -19 16 -15 18
rect -1 16 3 18
<< ptransistor >>
rect 15 42 19 44
rect 33 42 39 44
rect 48 42 60 44
rect 15 36 19 38
rect 33 36 39 38
rect 15 28 19 30
rect 33 28 39 30
rect 49 24 55 26
rect 15 22 19 24
rect 33 22 39 24
<< polysilicon >>
rect -22 48 -19 50
rect -15 48 -1 50
rect 3 48 6 50
rect -22 42 -19 44
rect -15 42 -1 44
rect 3 42 15 44
rect 19 42 33 44
rect 39 42 42 44
rect 45 42 48 44
rect 60 42 63 44
rect -22 36 -19 38
rect -15 36 -12 38
rect -22 34 -21 36
rect -23 30 -21 34
rect -9 30 -7 42
rect -4 36 -1 38
rect 3 36 15 38
rect 19 36 27 38
rect 30 36 33 38
rect 39 36 43 38
rect -35 28 -33 30
rect -29 28 -26 30
rect -23 28 -19 30
rect -15 28 -12 30
rect -9 28 -1 30
rect 3 28 15 30
rect 19 28 22 30
rect 25 24 27 36
rect 41 34 43 36
rect 30 28 33 30
rect 39 28 43 30
rect 46 24 49 26
rect 55 24 57 26
rect -22 22 -19 24
rect -15 22 -1 24
rect 3 22 15 24
rect 19 22 33 24
rect 39 22 42 24
rect -22 16 -19 18
rect -15 16 -1 18
rect 3 16 6 18
<< ndcontact >>
rect -19 51 -15 55
rect -1 51 3 55
rect -33 35 -29 39
rect -19 31 -15 35
rect -1 31 3 35
rect -33 21 -29 25
rect -19 11 -15 15
rect -1 11 3 15
<< pdcontact >>
rect 15 45 19 49
rect 33 45 39 49
rect 48 45 60 49
rect 56 37 60 41
rect 15 31 19 35
rect 33 31 37 35
rect 48 30 52 34
rect 15 17 19 21
rect 33 17 39 21
rect 49 17 55 21
<< polycontact >>
rect -39 28 -35 32
rect -26 34 -22 38
rect 41 30 45 34
rect 57 24 61 28
<< metal1 >>
rect -19 51 3 55
rect 15 45 60 49
rect -33 38 -29 39
rect -25 38 44 41
rect -33 35 -22 38
rect -26 34 -22 35
rect -39 31 -35 32
rect -19 31 37 35
rect -39 28 -15 31
rect 33 27 37 31
rect 41 34 44 38
rect 56 37 60 41
rect 41 30 52 34
rect 57 28 60 37
rect 57 27 61 28
rect -33 15 -29 25
rect 33 24 61 27
rect 15 17 55 21
rect -33 11 3 15
<< labels >>
rlabel polysilicon 40 43 40 43 1 b
rlabel polysilicon 40 23 40 23 1 a
rlabel polysilicon -20 43 -20 43 3 b
rlabel polysilicon -20 23 -20 23 1 a
rlabel polysilicon -20 49 -20 49 1 _SReset!
rlabel polysilicon -20 17 -20 17 1 _SReset!
rlabel polysilicon 61 43 61 43 1 _PReset!
rlabel space 18 16 64 50 3 ^p
rlabel space -40 10 0 56 7 ^n
rlabel pdcontact 35 33 35 33 1 x
rlabel pdcontact 36 19 36 19 1 Vdd!
rlabel pdcontact 36 47 36 47 1 Vdd!
rlabel ndcontact 1 33 1 33 1 x
rlabel ndcontact 1 13 1 13 1 GND!
rlabel pdcontact 17 33 17 33 1 x
rlabel pdcontact 17 19 17 19 1 Vdd!
rlabel ndcontact 1 53 1 53 5 GND!
rlabel pdcontact 17 47 17 47 1 Vdd!
rlabel ndcontact -17 53 -17 53 5 GND!
rlabel ndcontact -17 13 -17 13 1 GND!
rlabel pdcontact 54 47 54 47 5 Vdd!
rlabel pdcontact 58 39 58 39 7 x
rlabel pdcontact 52 19 52 19 3 Vdd!
rlabel polycontact 59 26 59 26 7 x
rlabel ndcontact -17 33 -17 33 1 x
rlabel ndcontact -31 23 -31 23 1 GND!
rlabel polycontact -37 30 -37 30 3 x
<< end >>
