
/* ----------------------------------------------------------------------


   ----------------------------------------------------------------------
   file:    tlm_fuse_env.sv
   Date Created  :tlm_Fuse_Map_env.svh 25/7/2016
   Author        : dbenita
   Project       : TLM1 IP
   ----------------------------------------------------------------------
 
  TLM1 Soala FUSE ENV

  This file include the TLM1 IP configuration for fuses
 
 In this file the IP can add constraints on fuse and addd IP
 specific code for the IP fuses
 
 

*/

//Include tlm regs
import uvm_pkg::*;

`ifdef XVM
   import ovm_pkg::*;
   import xvm_pkg::*;
   `include "ovm_macros.svh"
   `include "sla_macros.svh"
`endif

import sla_pkg::*;
`include "uvm_macros.svh"
`include "slu_macros.svh"
  
class tlm_fuse_env extends toplevel_fuse_env;
   `uvm_component_utils(tlm_fuse_env);

`include "fusegen_api.vh"   // this file was generated by the SOCFUSEGEN tool
   
    // --------------------------
    function new( string n="tlm_fuse_env", uvm_component p = null);
        super.new( n, p);
    endfunction : new

  
    // --------------------------
    //virtual function void build_phase(uvm_phase phase);
    //  super.build_phase(phase);
    //endfunction : build_phase

  /*
   Function: connect()
   
   In this pahse the user can disbale the defualt constraints on the fuse
   */
   function void connect_phase(uvm_phase phase);
     super.connect_phase(phase);

     //Disable default fuse constraint
     tlm_fuse.tlm_fuse_tlm_fuse_fuse_1.set_default_constraint(0);
   endfunction // void

  
  /*
   constraint: tlm_fuse_1_c
   */
   constraint tlm_fuse_1_c {
			    tlm_fuse.tlm_fuse_tlm_fuse_fuse_1.cfg_val inside {8'h10,8'h15,8'h34,8'h67,8'hFF};
			    }
 
endclass : tlm_fuse_env
