magic
tech scmos
timestamp 965071231
<< ndiffusion >>
rect 26 120 34 121
rect 26 112 34 117
rect 26 104 34 109
rect 26 100 34 101
rect 15 92 19 97
rect 7 91 19 92
rect 26 91 34 92
rect 7 83 19 88
rect 26 83 34 88
rect 7 78 19 80
rect 7 70 11 78
rect 26 75 34 80
rect 7 69 19 70
rect 26 71 34 72
rect 7 65 19 66
rect 7 57 11 65
rect 7 56 19 57
rect 7 52 19 53
rect 7 44 9 52
rect 7 42 19 44
rect 7 38 19 39
<< pdiffusion >>
rect 57 130 88 131
rect 102 131 110 136
rect 94 130 110 131
rect 57 126 88 127
rect 57 118 65 126
rect 57 117 88 118
rect 94 126 110 127
rect 94 118 102 126
rect 94 117 110 118
rect 57 113 88 114
rect 80 105 88 113
rect 57 104 88 105
rect 94 113 110 114
rect 102 105 110 113
rect 94 104 110 105
rect 57 100 88 101
rect 94 100 110 101
rect 102 92 110 100
rect 94 91 110 92
rect 94 87 110 88
rect 57 78 73 79
rect 108 79 110 87
rect 94 78 110 79
rect 57 74 73 75
rect 57 66 65 74
rect 94 74 110 75
rect 94 69 102 74
rect 57 65 73 66
rect 57 61 73 62
rect 57 52 73 53
rect 57 48 73 49
<< ntransistor >>
rect 26 117 34 120
rect 26 109 34 112
rect 26 101 34 104
rect 7 88 19 91
rect 26 88 34 91
rect 7 80 19 83
rect 26 80 34 83
rect 26 72 34 75
rect 7 66 19 69
rect 7 53 19 56
rect 7 39 19 42
<< ptransistor >>
rect 57 127 88 130
rect 94 127 110 130
rect 57 114 88 117
rect 94 114 110 117
rect 57 101 88 104
rect 94 101 110 104
rect 94 88 110 91
rect 57 75 73 78
rect 94 75 110 78
rect 57 62 73 65
rect 57 49 73 52
<< polysilicon >>
rect 44 127 57 130
rect 88 127 94 130
rect 110 127 114 130
rect 44 120 47 127
rect 22 117 26 120
rect 34 117 47 120
rect 52 114 57 117
rect 88 114 94 117
rect 110 114 114 117
rect 52 112 55 114
rect 22 109 26 112
rect 34 109 55 112
rect 22 101 26 104
rect 34 101 57 104
rect 88 101 94 104
rect 110 101 114 104
rect 3 88 7 91
rect 19 88 26 91
rect 34 88 55 91
rect 90 88 94 91
rect 110 88 112 91
rect 3 80 7 83
rect 19 80 26 83
rect 34 80 47 83
rect 21 72 26 75
rect 34 72 39 75
rect 21 69 24 72
rect 3 66 7 69
rect 19 66 24 69
rect 36 57 39 72
rect 44 65 47 80
rect 52 78 55 88
rect 52 75 57 78
rect 73 75 77 78
rect 90 75 94 78
rect 110 75 114 78
rect 44 62 57 65
rect 73 62 77 65
rect 5 53 7 56
rect 19 53 23 56
rect 36 54 55 57
rect 52 52 55 54
rect 52 49 57 52
rect 73 49 77 52
rect 3 39 7 42
rect 19 39 39 42
<< ndcontact >>
rect 26 121 34 129
rect 7 92 15 100
rect 26 92 34 100
rect 11 70 19 78
rect 11 57 19 65
rect 26 63 34 71
rect 9 44 19 52
rect 7 30 19 38
<< pdcontact >>
rect 57 131 88 139
rect 94 131 102 139
rect 65 118 88 126
rect 102 118 110 126
rect 57 105 80 113
rect 94 105 102 113
rect 57 92 88 100
rect 94 92 102 100
rect 57 79 73 87
rect 94 79 108 87
rect 65 66 73 74
rect 102 66 110 74
rect 57 53 73 61
rect 57 40 73 48
<< polycontact >>
rect 112 83 120 91
rect 82 70 90 78
rect -3 48 5 56
rect 39 39 47 47
<< metal1 >>
rect 57 131 88 139
rect 94 131 102 139
rect 26 121 34 129
rect 57 113 61 131
rect 65 118 88 126
rect 94 113 98 131
rect 102 118 110 126
rect 57 105 80 113
rect 94 109 102 113
rect 84 105 102 109
rect 84 100 90 105
rect 106 100 110 118
rect 7 96 15 100
rect 26 96 90 100
rect 3 92 15 96
rect 22 92 90 96
rect 94 96 110 100
rect 94 92 102 96
rect 3 65 7 92
rect 22 82 26 92
rect 14 78 26 82
rect 11 70 19 78
rect 3 61 19 65
rect 11 57 19 61
rect -3 48 5 56
rect 26 52 34 71
rect 0 38 5 48
rect 9 44 34 52
rect 39 47 43 92
rect 57 79 73 87
rect 57 61 61 79
rect 82 74 90 92
rect 65 66 90 74
rect 94 79 108 87
rect 112 83 120 91
rect 57 53 73 61
rect 94 48 98 79
rect 112 74 117 83
rect 39 39 47 47
rect 57 40 98 48
rect 102 69 117 74
rect 102 66 110 69
rect 0 35 19 38
rect 102 35 107 66
rect 0 33 107 35
rect 7 30 107 33
<< labels >>
rlabel polysilicon 111 102 111 102 1 a
rlabel metal1 98 109 98 109 1 x
rlabel metal1 98 135 98 135 5 x
rlabel metal1 102 83 102 83 1 Vdd!
rlabel polysilicon 74 50 74 50 1 a
rlabel polysilicon 6 89 6 89 1 _b1
rlabel polysilicon 6 81 6 81 1 _b0
rlabel metal1 30 96 30 96 5 x
rlabel metal1 15 74 15 74 1 x
rlabel metal1 69 96 69 96 1 x
rlabel metal1 69 70 69 70 1 x
rlabel polysilicon 25 118 25 118 1 _b1
rlabel polysilicon 25 110 25 110 1 _b0
rlabel metal1 30 125 30 125 5 GND!
rlabel metal1 30 67 30 67 1 GND!
rlabel metal1 69 122 69 122 1 Vdd!
rlabel metal1 65 44 65 44 1 Vdd!
rlabel metal1 14 48 14 48 1 GND!
rlabel space 2 70 27 130 7 ^n
rlabel space -4 29 25 69 7 ^n
rlabel space 72 29 121 140 3 ^p
<< end >>
