`define pargpio 		 `soc.pargpio
`define pmu_wrapper1 		 `pargpio.pmu_wrapper1

