///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cm_usage_map_pkg.vh                                
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_CM_USAGE_MAP_PKG_VH
`define MBY_PPE_CM_USAGE_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_cm_usage_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_cm_usage_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_cm_usage_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_cm_usage_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic [14:0] WATERMARK;  // RW
} CM_TX_TC_PRIVATE_WM_t;

localparam CM_TX_TC_PRIVATE_WM_REG_STRIDE = 48'h8;
localparam CM_TX_TC_PRIVATE_WM_REG_ENTRIES = 8;
localparam CM_TX_TC_PRIVATE_WM_REGFILE_STRIDE = 48'h40;
localparam CM_TX_TC_PRIVATE_WM_REGFILE_ENTRIES = 64;
localparam CM_TX_TC_PRIVATE_WM_CR_ADDR = 48'h0;
localparam CM_TX_TC_PRIVATE_WM_SIZE = 64;
localparam CM_TX_TC_PRIVATE_WM_WATERMARK_LO = 0;
localparam CM_TX_TC_PRIVATE_WM_WATERMARK_HI = 14;
localparam CM_TX_TC_PRIVATE_WM_WATERMARK_RESET = 15'h7fff;
localparam CM_TX_TC_PRIVATE_WM_USEMASK = 64'h7FFF;
localparam CM_TX_TC_PRIVATE_WM_RO_MASK = 64'h0;
localparam CM_TX_TC_PRIVATE_WM_WO_MASK = 64'h0;
localparam CM_TX_TC_PRIVATE_WM_RESET = 64'h7FFF;

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic [14:0] WATERMARK;  // RW
} CM_TX_TC_HOG_WM_t;

localparam CM_TX_TC_HOG_WM_REG_STRIDE = 48'h8;
localparam CM_TX_TC_HOG_WM_REG_ENTRIES = 8;
localparam CM_TX_TC_HOG_WM_REGFILE_STRIDE = 48'h40;
localparam CM_TX_TC_HOG_WM_REGFILE_ENTRIES = 64;
localparam CM_TX_TC_HOG_WM_CR_ADDR = 48'h1000;
localparam CM_TX_TC_HOG_WM_SIZE = 64;
localparam CM_TX_TC_HOG_WM_WATERMARK_LO = 0;
localparam CM_TX_TC_HOG_WM_WATERMARK_HI = 14;
localparam CM_TX_TC_HOG_WM_WATERMARK_RESET = 15'h7fff;
localparam CM_TX_TC_HOG_WM_USEMASK = 64'h7FFF;
localparam CM_TX_TC_HOG_WM_RO_MASK = 64'h0;
localparam CM_TX_TC_HOG_WM_WO_MASK = 64'h0;
localparam CM_TX_TC_HOG_WM_RESET = 64'h7FFF;

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic [14:0] WATERMARK;  // RW
} CM_RX_SMP_PRIVATE_WM_t;

localparam CM_RX_SMP_PRIVATE_WM_REG_STRIDE = 48'h8;
localparam CM_RX_SMP_PRIVATE_WM_REG_ENTRIES = 2;
localparam CM_RX_SMP_PRIVATE_WM_REGFILE_STRIDE = 48'h10;
localparam CM_RX_SMP_PRIVATE_WM_REGFILE_ENTRIES = 32;
localparam CM_RX_SMP_PRIVATE_WM_CR_ADDR = 48'h2000;
localparam CM_RX_SMP_PRIVATE_WM_SIZE = 64;
localparam CM_RX_SMP_PRIVATE_WM_WATERMARK_LO = 0;
localparam CM_RX_SMP_PRIVATE_WM_WATERMARK_HI = 14;
localparam CM_RX_SMP_PRIVATE_WM_WATERMARK_RESET = 15'h7fff;
localparam CM_RX_SMP_PRIVATE_WM_USEMASK = 64'h7FFF;
localparam CM_RX_SMP_PRIVATE_WM_RO_MASK = 64'h0;
localparam CM_RX_SMP_PRIVATE_WM_WO_MASK = 64'h0;
localparam CM_RX_SMP_PRIVATE_WM_RESET = 64'h7FFF;

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic [14:0] WATERMARK;  // RW
} CM_RX_SMP_HOG_WM_t;

localparam CM_RX_SMP_HOG_WM_REG_STRIDE = 48'h8;
localparam CM_RX_SMP_HOG_WM_REG_ENTRIES = 2;
localparam CM_RX_SMP_HOG_WM_REGFILE_STRIDE = 48'h10;
localparam CM_RX_SMP_HOG_WM_REGFILE_ENTRIES = 32;
localparam CM_RX_SMP_HOG_WM_CR_ADDR = 48'h2200;
localparam CM_RX_SMP_HOG_WM_SIZE = 64;
localparam CM_RX_SMP_HOG_WM_WATERMARK_LO = 0;
localparam CM_RX_SMP_HOG_WM_WATERMARK_HI = 14;
localparam CM_RX_SMP_HOG_WM_WATERMARK_RESET = 15'h7fff;
localparam CM_RX_SMP_HOG_WM_USEMASK = 64'h7FFF;
localparam CM_RX_SMP_HOG_WM_RO_MASK = 64'h0;
localparam CM_RX_SMP_HOG_WM_WO_MASK = 64'h0;
localparam CM_RX_SMP_HOG_WM_RESET = 64'h7FFF;

typedef struct packed {
    logic [33:0] reserved0;  // RSVD
    logic [14:0] PAUSE_OFF;  // RW
    logic [14:0] PAUSE_ON;  // RW
} CM_RX_SMP_PAUSE_WM_t;

localparam CM_RX_SMP_PAUSE_WM_REG_STRIDE = 48'h8;
localparam CM_RX_SMP_PAUSE_WM_REG_ENTRIES = 2;
localparam CM_RX_SMP_PAUSE_WM_REGFILE_STRIDE = 48'h10;
localparam CM_RX_SMP_PAUSE_WM_REGFILE_ENTRIES = 32;
localparam CM_RX_SMP_PAUSE_WM_CR_ADDR = 48'h2400;
localparam CM_RX_SMP_PAUSE_WM_SIZE = 64;
localparam CM_RX_SMP_PAUSE_WM_PAUSE_OFF_LO = 15;
localparam CM_RX_SMP_PAUSE_WM_PAUSE_OFF_HI = 29;
localparam CM_RX_SMP_PAUSE_WM_PAUSE_OFF_RESET = 15'h7fff;
localparam CM_RX_SMP_PAUSE_WM_PAUSE_ON_LO = 0;
localparam CM_RX_SMP_PAUSE_WM_PAUSE_ON_HI = 14;
localparam CM_RX_SMP_PAUSE_WM_PAUSE_ON_RESET = 15'h7fff;
localparam CM_RX_SMP_PAUSE_WM_USEMASK = 64'h3FFFFFFF;
localparam CM_RX_SMP_PAUSE_WM_RO_MASK = 64'h0;
localparam CM_RX_SMP_PAUSE_WM_WO_MASK = 64'h0;
localparam CM_RX_SMP_PAUSE_WM_RESET = 64'h3FFFFFFF;

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic [14:0] WATERMARK;  // RW
} CM_SHARED_WM_t;

localparam CM_SHARED_WM_REG_STRIDE = 48'h8;
localparam CM_SHARED_WM_REG_ENTRIES = 8;
localparam CM_SHARED_WM_CR_ADDR = 48'h2600;
localparam CM_SHARED_WM_SIZE = 64;
localparam CM_SHARED_WM_WATERMARK_LO = 0;
localparam CM_SHARED_WM_WATERMARK_HI = 14;
localparam CM_SHARED_WM_WATERMARK_RESET = 15'h21c;
localparam CM_SHARED_WM_USEMASK = 64'h7FFF;
localparam CM_SHARED_WM_RO_MASK = 64'h0;
localparam CM_SHARED_WM_WO_MASK = 64'h0;
localparam CM_SHARED_WM_RESET = 64'h21C;

typedef struct packed {
    logic [33:0] reserved0;  // RSVD
    logic [14:0] HOG_SEGMENT_LIMIT;  // RW
    logic [14:0] SOFT_DROP_SEGMENT_LIMIT;  // RW
} CM_SOFTDROP_WM_t;

localparam CM_SOFTDROP_WM_REG_STRIDE = 48'h8;
localparam CM_SOFTDROP_WM_REG_ENTRIES = 8;
localparam CM_SOFTDROP_WM_CR_ADDR = 48'h2640;
localparam CM_SOFTDROP_WM_SIZE = 64;
localparam CM_SOFTDROP_WM_HOG_SEGMENT_LIMIT_LO = 15;
localparam CM_SOFTDROP_WM_HOG_SEGMENT_LIMIT_HI = 29;
localparam CM_SOFTDROP_WM_HOG_SEGMENT_LIMIT_RESET = 15'h7fff;
localparam CM_SOFTDROP_WM_SOFT_DROP_SEGMENT_LIMIT_LO = 0;
localparam CM_SOFTDROP_WM_SOFT_DROP_SEGMENT_LIMIT_HI = 14;
localparam CM_SOFTDROP_WM_SOFT_DROP_SEGMENT_LIMIT_RESET = 15'h7fff;
localparam CM_SOFTDROP_WM_USEMASK = 64'h3FFFFFFF;
localparam CM_SOFTDROP_WM_RO_MASK = 64'h0;
localparam CM_SOFTDROP_WM_WO_MASK = 64'h0;
localparam CM_SOFTDROP_WM_RESET = 64'h3FFFFFFF;

typedef struct packed {
    logic [33:0] reserved0;  // RSVD
    logic [14:0] PAUSE_OFF;  // RW
    logic [14:0] PAUSE_ON;  // RW
} CM_SHARED_SMP_PAUSE_WM_t;

localparam CM_SHARED_SMP_PAUSE_WM_REG_STRIDE = 48'h8;
localparam CM_SHARED_SMP_PAUSE_WM_REG_ENTRIES = 2;
localparam CM_SHARED_SMP_PAUSE_WM_CR_ADDR = 48'h2680;
localparam CM_SHARED_SMP_PAUSE_WM_SIZE = 64;
localparam CM_SHARED_SMP_PAUSE_WM_PAUSE_OFF_LO = 15;
localparam CM_SHARED_SMP_PAUSE_WM_PAUSE_OFF_HI = 29;
localparam CM_SHARED_SMP_PAUSE_WM_PAUSE_OFF_RESET = 15'h7fff;
localparam CM_SHARED_SMP_PAUSE_WM_PAUSE_ON_LO = 0;
localparam CM_SHARED_SMP_PAUSE_WM_PAUSE_ON_HI = 14;
localparam CM_SHARED_SMP_PAUSE_WM_PAUSE_ON_RESET = 15'h7fff;
localparam CM_SHARED_SMP_PAUSE_WM_USEMASK = 64'h3FFFFFFF;
localparam CM_SHARED_SMP_PAUSE_WM_RO_MASK = 64'h0;
localparam CM_SHARED_SMP_PAUSE_WM_WO_MASK = 64'h0;
localparam CM_SHARED_SMP_PAUSE_WM_RESET = 64'h3FFFFFFF;

typedef struct packed {
    logic [48:0] reserved0;  // RSVD
    logic [14:0] WATERMARK;  // RW
} CM_GLOBAL_WM_t;

localparam CM_GLOBAL_WM_REG_STRIDE = 48'h8;
localparam CM_GLOBAL_WM_REG_ENTRIES = 1;
localparam [47:0] CM_GLOBAL_WM_CR_ADDR = 48'h2690;
localparam CM_GLOBAL_WM_SIZE = 64;
localparam CM_GLOBAL_WM_WATERMARK_LO = 0;
localparam CM_GLOBAL_WM_WATERMARK_HI = 14;
localparam CM_GLOBAL_WM_WATERMARK_RESET = 15'h5e20;
localparam CM_GLOBAL_WM_USEMASK = 64'h7FFF;
localparam CM_GLOBAL_WM_RO_MASK = 64'h0;
localparam CM_GLOBAL_WM_WO_MASK = 64'h0;
localparam CM_GLOBAL_WM_RESET = 64'h5E20;

typedef struct packed {
    logic [58:0] reserved0;  // RSVD
    logic  [4:0] PHYS_PORT;  // RW
} CM_PAUSE_PHYS_PORT_CFG_t;

localparam CM_PAUSE_PHYS_PORT_CFG_REG_STRIDE = 48'h8;
localparam CM_PAUSE_PHYS_PORT_CFG_REG_ENTRIES = 32;
localparam CM_PAUSE_PHYS_PORT_CFG_CR_ADDR = 48'h2700;
localparam CM_PAUSE_PHYS_PORT_CFG_SIZE = 64;
localparam CM_PAUSE_PHYS_PORT_CFG_PHYS_PORT_LO = 0;
localparam CM_PAUSE_PHYS_PORT_CFG_PHYS_PORT_HI = 4;
localparam CM_PAUSE_PHYS_PORT_CFG_PHYS_PORT_RESET = 5'h0;
localparam CM_PAUSE_PHYS_PORT_CFG_USEMASK = 64'h1F;
localparam CM_PAUSE_PHYS_PORT_CFG_RO_MASK = 64'h0;
localparam CM_PAUSE_PHYS_PORT_CFG_WO_MASK = 64'h0;
localparam CM_PAUSE_PHYS_PORT_CFG_RESET = 64'h0;

typedef struct packed {
    logic [59:0] reserved0;  // RSVD
    logic  [1:0] FORCE_OFF;  // RW
    logic  [1:0] FORCE_ON;  // RW
} CM_FORCE_PAUSE_CFG_t;

localparam CM_FORCE_PAUSE_CFG_REG_STRIDE = 48'h8;
localparam CM_FORCE_PAUSE_CFG_REG_ENTRIES = 1;
localparam CM_FORCE_PAUSE_CFG_CR_ADDR = 48'h2800;
localparam CM_FORCE_PAUSE_CFG_SIZE = 64;
localparam CM_FORCE_PAUSE_CFG_FORCE_OFF_LO = 2;
localparam CM_FORCE_PAUSE_CFG_FORCE_OFF_HI = 3;
localparam CM_FORCE_PAUSE_CFG_FORCE_OFF_RESET = 2'h0;
localparam CM_FORCE_PAUSE_CFG_FORCE_ON_LO = 0;
localparam CM_FORCE_PAUSE_CFG_FORCE_ON_HI = 1;
localparam CM_FORCE_PAUSE_CFG_FORCE_ON_RESET = 2'h0;
localparam CM_FORCE_PAUSE_CFG_USEMASK = 64'hF;
localparam CM_FORCE_PAUSE_CFG_RO_MASK = 64'h0;
localparam CM_FORCE_PAUSE_CFG_WO_MASK = 64'h0;
localparam CM_FORCE_PAUSE_CFG_RESET = 64'h0;

typedef struct packed {
    logic [18:0] reserved0;  // RSVD
    logic  [7:0] UPDATE_INTERVAL;  // RW
    logic  [3:0] W;  // RW
    logic  [2:0] TC;  // RW
    logic [14:0] MIN_TH;  // RW
    logic [14:0] MAX_TH;  // RW
} CM_AQM_EWMA_CFG_t;

localparam CM_AQM_EWMA_CFG_REG_STRIDE = 48'h8;
localparam CM_AQM_EWMA_CFG_REG_ENTRIES = 2;
localparam CM_AQM_EWMA_CFG_REGFILE_STRIDE = 48'h10;
localparam CM_AQM_EWMA_CFG_REGFILE_ENTRIES = 64;
localparam CM_AQM_EWMA_CFG_CR_ADDR = 48'h2C00;
localparam CM_AQM_EWMA_CFG_SIZE = 64;
localparam CM_AQM_EWMA_CFG_UPDATE_INTERVAL_LO = 37;
localparam CM_AQM_EWMA_CFG_UPDATE_INTERVAL_HI = 44;
localparam CM_AQM_EWMA_CFG_UPDATE_INTERVAL_RESET = 8'h0;
localparam CM_AQM_EWMA_CFG_W_LO = 33;
localparam CM_AQM_EWMA_CFG_W_HI = 36;
localparam CM_AQM_EWMA_CFG_W_RESET = 4'h8;
localparam CM_AQM_EWMA_CFG_TC_LO = 30;
localparam CM_AQM_EWMA_CFG_TC_HI = 32;
localparam CM_AQM_EWMA_CFG_TC_RESET = 3'h0;
localparam CM_AQM_EWMA_CFG_MIN_TH_LO = 15;
localparam CM_AQM_EWMA_CFG_MIN_TH_HI = 29;
localparam CM_AQM_EWMA_CFG_MIN_TH_RESET = 15'h96;
localparam CM_AQM_EWMA_CFG_MAX_TH_LO = 0;
localparam CM_AQM_EWMA_CFG_MAX_TH_HI = 14;
localparam CM_AQM_EWMA_CFG_MAX_TH_RESET = 15'h384;
localparam CM_AQM_EWMA_CFG_USEMASK = 64'h1FFFFFFFFFFF;
localparam CM_AQM_EWMA_CFG_RO_MASK = 64'h0;
localparam CM_AQM_EWMA_CFG_WO_MASK = 64'h0;
localparam CM_AQM_EWMA_CFG_RESET = 64'h10004B0384;

typedef struct packed {
    logic [45:0] reserved0;  // RSVD
    logic  [2:0] TC;  // RW
    logic [14:0] THRESHOLD;  // RW
} CM_AQM_DCTCP_CFG_t;

localparam CM_AQM_DCTCP_CFG_REG_STRIDE = 48'h8;
localparam CM_AQM_DCTCP_CFG_REG_ENTRIES = 2;
localparam CM_AQM_DCTCP_CFG_REGFILE_STRIDE = 48'h10;
localparam CM_AQM_DCTCP_CFG_REGFILE_ENTRIES = 64;
localparam CM_AQM_DCTCP_CFG_CR_ADDR = 48'h3000;
localparam CM_AQM_DCTCP_CFG_SIZE = 64;
localparam CM_AQM_DCTCP_CFG_TC_LO = 15;
localparam CM_AQM_DCTCP_CFG_TC_HI = 17;
localparam CM_AQM_DCTCP_CFG_TC_RESET = 3'h0;
localparam CM_AQM_DCTCP_CFG_THRESHOLD_LO = 0;
localparam CM_AQM_DCTCP_CFG_THRESHOLD_HI = 14;
localparam CM_AQM_DCTCP_CFG_THRESHOLD_RESET = 15'h7FFF;
localparam CM_AQM_DCTCP_CFG_USEMASK = 64'h3FFFF;
localparam CM_AQM_DCTCP_CFG_RO_MASK = 64'h0;
localparam CM_AQM_DCTCP_CFG_WO_MASK = 64'h0;
localparam CM_AQM_DCTCP_CFG_RESET = 64'h7FFF;

typedef struct packed {
    logic [57:0] reserved0;  // RSVD
    logic  [0:0] SWEEPER_EN;  // RW
    logic  [4:0] NUM_SWEEPER_PORTS;  // RW
} CM_GLOBAL_CFG_t;

localparam CM_GLOBAL_CFG_REG_STRIDE = 48'h8;
localparam CM_GLOBAL_CFG_REG_ENTRIES = 1;
localparam [47:0] CM_GLOBAL_CFG_CR_ADDR = 48'h3400;
localparam CM_GLOBAL_CFG_SIZE = 64;
localparam CM_GLOBAL_CFG_SWEEPER_EN_LO = 5;
localparam CM_GLOBAL_CFG_SWEEPER_EN_HI = 5;
localparam CM_GLOBAL_CFG_SWEEPER_EN_RESET = 1'h0;
localparam CM_GLOBAL_CFG_NUM_SWEEPER_PORTS_LO = 0;
localparam CM_GLOBAL_CFG_NUM_SWEEPER_PORTS_HI = 4;
localparam CM_GLOBAL_CFG_NUM_SWEEPER_PORTS_RESET = 5'h0;
localparam CM_GLOBAL_CFG_USEMASK = 64'h3F;
localparam CM_GLOBAL_CFG_RO_MASK = 64'h0;
localparam CM_GLOBAL_CFG_WO_MASK = 64'h0;
localparam CM_GLOBAL_CFG_RESET = 64'h0;

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic [23:0] ENABLE_MASK;  // RW
} CM_SHARED_SMP_PAUSE_CFG_t;

localparam CM_SHARED_SMP_PAUSE_CFG_REG_STRIDE = 48'h8;
localparam CM_SHARED_SMP_PAUSE_CFG_REG_ENTRIES = 2;
localparam CM_SHARED_SMP_PAUSE_CFG_CR_ADDR = 48'h3410;
localparam CM_SHARED_SMP_PAUSE_CFG_SIZE = 64;
localparam CM_SHARED_SMP_PAUSE_CFG_ENABLE_MASK_LO = 0;
localparam CM_SHARED_SMP_PAUSE_CFG_ENABLE_MASK_HI = 23;
localparam CM_SHARED_SMP_PAUSE_CFG_ENABLE_MASK_RESET = 24'h0;
localparam CM_SHARED_SMP_PAUSE_CFG_USEMASK = 64'hFFFFFF;
localparam CM_SHARED_SMP_PAUSE_CFG_RO_MASK = 64'h0;
localparam CM_SHARED_SMP_PAUSE_CFG_WO_MASK = 64'h0;
localparam CM_SHARED_SMP_PAUSE_CFG_RESET = 64'h0;

typedef struct packed {
    logic [55:0] reserved0;  // RSVD
    logic  [0:0] SMP_7;  // RW
    logic  [0:0] SMP_6;  // RW
    logic  [0:0] SMP_5;  // RW
    logic  [0:0] SMP_4;  // RW
    logic  [0:0] SMP_3;  // RW
    logic  [0:0] SMP_2;  // RW
    logic  [0:0] SMP_1;  // RW
    logic  [0:0] SMP_0;  // RW
} CM_SWEEPER_TC_TO_SMP_t;

localparam CM_SWEEPER_TC_TO_SMP_REG_STRIDE = 48'h8;
localparam CM_SWEEPER_TC_TO_SMP_REG_ENTRIES = 1;
localparam [47:0] CM_SWEEPER_TC_TO_SMP_CR_ADDR = 48'h3420;
localparam CM_SWEEPER_TC_TO_SMP_SIZE = 64;
localparam CM_SWEEPER_TC_TO_SMP_SMP_7_LO = 7;
localparam CM_SWEEPER_TC_TO_SMP_SMP_7_HI = 7;
localparam CM_SWEEPER_TC_TO_SMP_SMP_7_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_6_LO = 6;
localparam CM_SWEEPER_TC_TO_SMP_SMP_6_HI = 6;
localparam CM_SWEEPER_TC_TO_SMP_SMP_6_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_5_LO = 5;
localparam CM_SWEEPER_TC_TO_SMP_SMP_5_HI = 5;
localparam CM_SWEEPER_TC_TO_SMP_SMP_5_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_4_LO = 4;
localparam CM_SWEEPER_TC_TO_SMP_SMP_4_HI = 4;
localparam CM_SWEEPER_TC_TO_SMP_SMP_4_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_3_LO = 3;
localparam CM_SWEEPER_TC_TO_SMP_SMP_3_HI = 3;
localparam CM_SWEEPER_TC_TO_SMP_SMP_3_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_2_LO = 2;
localparam CM_SWEEPER_TC_TO_SMP_SMP_2_HI = 2;
localparam CM_SWEEPER_TC_TO_SMP_SMP_2_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_1_LO = 1;
localparam CM_SWEEPER_TC_TO_SMP_SMP_1_HI = 1;
localparam CM_SWEEPER_TC_TO_SMP_SMP_1_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_0_LO = 0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_0_HI = 0;
localparam CM_SWEEPER_TC_TO_SMP_SMP_0_RESET = 1'h0;
localparam CM_SWEEPER_TC_TO_SMP_USEMASK = 64'hFF;
localparam CM_SWEEPER_TC_TO_SMP_RO_MASK = 64'h0;
localparam CM_SWEEPER_TC_TO_SMP_WO_MASK = 64'h0;
localparam CM_SWEEPER_TC_TO_SMP_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RO/V
} CM_GLOBAL_USAGE_t;

localparam CM_GLOBAL_USAGE_REG_STRIDE = 48'h8;
localparam CM_GLOBAL_USAGE_REG_ENTRIES = 1;
localparam [47:0] CM_GLOBAL_USAGE_CR_ADDR = 48'h3428;
localparam CM_GLOBAL_USAGE_SIZE = 64;
localparam CM_GLOBAL_USAGE_COUNT_LO = 0;
localparam CM_GLOBAL_USAGE_COUNT_HI = 15;
localparam CM_GLOBAL_USAGE_COUNT_RESET = 16'h0;
localparam CM_GLOBAL_USAGE_USEMASK = 64'hFFFF;
localparam CM_GLOBAL_USAGE_RO_MASK = 64'hFFFF;
localparam CM_GLOBAL_USAGE_WO_MASK = 64'h0;
localparam CM_GLOBAL_USAGE_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RW/V
} CM_GLOBAL_USAGE_MAX_t;

localparam CM_GLOBAL_USAGE_MAX_REG_STRIDE = 48'h8;
localparam CM_GLOBAL_USAGE_MAX_REG_ENTRIES = 1;
localparam [47:0] CM_GLOBAL_USAGE_MAX_CR_ADDR = 48'h3430;
localparam CM_GLOBAL_USAGE_MAX_SIZE = 64;
localparam CM_GLOBAL_USAGE_MAX_COUNT_LO = 0;
localparam CM_GLOBAL_USAGE_MAX_COUNT_HI = 15;
localparam CM_GLOBAL_USAGE_MAX_COUNT_RESET = 16'h0;
localparam CM_GLOBAL_USAGE_MAX_USEMASK = 64'hFFFF;
localparam CM_GLOBAL_USAGE_MAX_RO_MASK = 64'h0;
localparam CM_GLOBAL_USAGE_MAX_WO_MASK = 64'h0;
localparam CM_GLOBAL_USAGE_MAX_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RO/V
} CM_MCAST_EPOCH_USAGE_t;

localparam CM_MCAST_EPOCH_USAGE_REG_STRIDE = 48'h8;
localparam CM_MCAST_EPOCH_USAGE_REG_ENTRIES = 2;
localparam CM_MCAST_EPOCH_USAGE_CR_ADDR = 48'h3440;
localparam CM_MCAST_EPOCH_USAGE_SIZE = 64;
localparam CM_MCAST_EPOCH_USAGE_COUNT_LO = 0;
localparam CM_MCAST_EPOCH_USAGE_COUNT_HI = 15;
localparam CM_MCAST_EPOCH_USAGE_COUNT_RESET = 16'h0;
localparam CM_MCAST_EPOCH_USAGE_USEMASK = 64'hFFFF;
localparam CM_MCAST_EPOCH_USAGE_RO_MASK = 64'hFFFF;
localparam CM_MCAST_EPOCH_USAGE_WO_MASK = 64'h0;
localparam CM_MCAST_EPOCH_USAGE_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RO/V
} CM_SHARED_SMP_USAGE_t;

localparam CM_SHARED_SMP_USAGE_REG_STRIDE = 48'h8;
localparam CM_SHARED_SMP_USAGE_REG_ENTRIES = 2;
localparam CM_SHARED_SMP_USAGE_CR_ADDR = 48'h3450;
localparam CM_SHARED_SMP_USAGE_SIZE = 64;
localparam CM_SHARED_SMP_USAGE_COUNT_LO = 0;
localparam CM_SHARED_SMP_USAGE_COUNT_HI = 15;
localparam CM_SHARED_SMP_USAGE_COUNT_RESET = 16'h0;
localparam CM_SHARED_SMP_USAGE_USEMASK = 64'hFFFF;
localparam CM_SHARED_SMP_USAGE_RO_MASK = 64'hFFFF;
localparam CM_SHARED_SMP_USAGE_WO_MASK = 64'h0;
localparam CM_SHARED_SMP_USAGE_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RO/V
} CM_SMP_USAGE_t;

localparam CM_SMP_USAGE_REG_STRIDE = 48'h8;
localparam CM_SMP_USAGE_REG_ENTRIES = 2;
localparam CM_SMP_USAGE_CR_ADDR = 48'h3460;
localparam CM_SMP_USAGE_SIZE = 64;
localparam CM_SMP_USAGE_COUNT_LO = 0;
localparam CM_SMP_USAGE_COUNT_HI = 15;
localparam CM_SMP_USAGE_COUNT_RESET = 16'h0;
localparam CM_SMP_USAGE_USEMASK = 64'hFFFF;
localparam CM_SMP_USAGE_RO_MASK = 64'hFFFF;
localparam CM_SMP_USAGE_WO_MASK = 64'h0;
localparam CM_SMP_USAGE_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RO/V
} CM_RX_SMP_USAGE_t;

localparam CM_RX_SMP_USAGE_REG_STRIDE = 48'h8;
localparam CM_RX_SMP_USAGE_REG_ENTRIES = 2;
localparam CM_RX_SMP_USAGE_REGFILE_STRIDE = 48'h10;
localparam CM_RX_SMP_USAGE_REGFILE_ENTRIES = 32;
localparam CM_RX_SMP_USAGE_CR_ADDR = 48'h3600;
localparam CM_RX_SMP_USAGE_SIZE = 64;
localparam CM_RX_SMP_USAGE_COUNT_LO = 0;
localparam CM_RX_SMP_USAGE_COUNT_HI = 15;
localparam CM_RX_SMP_USAGE_COUNT_RESET = 16'h0;
localparam CM_RX_SMP_USAGE_USEMASK = 64'hFFFF;
localparam CM_RX_SMP_USAGE_RO_MASK = 64'hFFFF;
localparam CM_RX_SMP_USAGE_WO_MASK = 64'h0;
localparam CM_RX_SMP_USAGE_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RW/V
} CM_RX_SMP_USAGE_MAX_t;

localparam CM_RX_SMP_USAGE_MAX_REG_STRIDE = 48'h8;
localparam CM_RX_SMP_USAGE_MAX_REG_ENTRIES = 2;
localparam CM_RX_SMP_USAGE_MAX_REGFILE_STRIDE = 48'h10;
localparam CM_RX_SMP_USAGE_MAX_REGFILE_ENTRIES = 4;
localparam CM_RX_SMP_USAGE_MAX_CR_ADDR = 48'h3800;
localparam CM_RX_SMP_USAGE_MAX_SIZE = 64;
localparam CM_RX_SMP_USAGE_MAX_COUNT_LO = 0;
localparam CM_RX_SMP_USAGE_MAX_COUNT_HI = 15;
localparam CM_RX_SMP_USAGE_MAX_COUNT_RESET = 16'h0;
localparam CM_RX_SMP_USAGE_MAX_USEMASK = 64'hFFFF;
localparam CM_RX_SMP_USAGE_MAX_RO_MASK = 64'h0;
localparam CM_RX_SMP_USAGE_MAX_WO_MASK = 64'h0;
localparam CM_RX_SMP_USAGE_MAX_RESET = 64'h0;

typedef struct packed {
    logic [43:0] reserved0;  // RSVD
    logic  [4:0] PORT3;  // RW
    logic  [4:0] PORT2;  // RW
    logic  [4:0] PORT1;  // RW
    logic  [4:0] PORT0;  // RW
} CM_RX_SMP_USAGE_MAX_CTRL_t;

localparam CM_RX_SMP_USAGE_MAX_CTRL_REG_STRIDE = 48'h8;
localparam CM_RX_SMP_USAGE_MAX_CTRL_REG_ENTRIES = 1;
localparam CM_RX_SMP_USAGE_MAX_CTRL_CR_ADDR = 48'h3840;
localparam CM_RX_SMP_USAGE_MAX_CTRL_SIZE = 64;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT3_LO = 15;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT3_HI = 19;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT3_RESET = 5'h0;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT2_LO = 10;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT2_HI = 14;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT2_RESET = 5'h0;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT1_LO = 5;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT1_HI = 9;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT1_RESET = 5'h0;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT0_LO = 0;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT0_HI = 4;
localparam CM_RX_SMP_USAGE_MAX_CTRL_PORT0_RESET = 5'h0;
localparam CM_RX_SMP_USAGE_MAX_CTRL_USEMASK = 64'hFFFFF;
localparam CM_RX_SMP_USAGE_MAX_CTRL_RO_MASK = 64'h0;
localparam CM_RX_SMP_USAGE_MAX_CTRL_WO_MASK = 64'h0;
localparam CM_RX_SMP_USAGE_MAX_CTRL_RESET = 64'h0;

typedef struct packed {
    logic [61:0] reserved0;  // RSVD
    logic  [0:0] SMP1;  // RO/V
    logic  [0:0] SMP0;  // RO/V
} CM_PAUSE_GEN_STATE_t;

localparam CM_PAUSE_GEN_STATE_REG_STRIDE = 48'h8;
localparam CM_PAUSE_GEN_STATE_REG_ENTRIES = 32;
localparam CM_PAUSE_GEN_STATE_CR_ADDR = 48'h3900;
localparam CM_PAUSE_GEN_STATE_SIZE = 64;
localparam CM_PAUSE_GEN_STATE_SMP1_LO = 1;
localparam CM_PAUSE_GEN_STATE_SMP1_HI = 1;
localparam CM_PAUSE_GEN_STATE_SMP1_RESET = 1'h0;
localparam CM_PAUSE_GEN_STATE_SMP0_LO = 0;
localparam CM_PAUSE_GEN_STATE_SMP0_HI = 0;
localparam CM_PAUSE_GEN_STATE_SMP0_RESET = 1'h0;
localparam CM_PAUSE_GEN_STATE_USEMASK = 64'h3;
localparam CM_PAUSE_GEN_STATE_RO_MASK = 64'h3;
localparam CM_PAUSE_GEN_STATE_WO_MASK = 64'h0;
localparam CM_PAUSE_GEN_STATE_RESET = 64'h0;

typedef struct packed {
    logic [47:0] reserved0;  // RSVD
    logic [15:0] COUNT;  // RO/V
} CM_TX_TC_USAGE_t;

localparam CM_TX_TC_USAGE_REG_STRIDE = 48'h8;
localparam CM_TX_TC_USAGE_REG_ENTRIES = 8;
localparam CM_TX_TC_USAGE_REGFILE_STRIDE = 48'h40;
localparam CM_TX_TC_USAGE_REGFILE_ENTRIES = 64;
localparam CM_TX_TC_USAGE_CR_ADDR = 48'h4000;
localparam CM_TX_TC_USAGE_SIZE = 64;
localparam CM_TX_TC_USAGE_COUNT_LO = 0;
localparam CM_TX_TC_USAGE_COUNT_HI = 15;
localparam CM_TX_TC_USAGE_COUNT_RESET = 16'h0;
localparam CM_TX_TC_USAGE_USEMASK = 64'hFFFF;
localparam CM_TX_TC_USAGE_RO_MASK = 64'hFFFF;
localparam CM_TX_TC_USAGE_WO_MASK = 64'h0;
localparam CM_TX_TC_USAGE_RESET = 64'h0;

typedef struct packed {
    logic [31:0] reserved0;  // RSVD
    logic  [7:0] INTERVAL;  // RO/V
    logic [15:0] EWMA_WHOLE;  // RO/V
    logic  [7:0] EWMA_FRAC;  // RO/V
} CM_TX_EWMA_t;

localparam CM_TX_EWMA_REG_STRIDE = 48'h8;
localparam CM_TX_EWMA_REG_ENTRIES = 2;
localparam CM_TX_EWMA_REGFILE_STRIDE = 48'h10;
localparam CM_TX_EWMA_REGFILE_ENTRIES = 64;
localparam CM_TX_EWMA_CR_ADDR = 48'h5000;
localparam CM_TX_EWMA_SIZE = 64;
localparam CM_TX_EWMA_INTERVAL_LO = 24;
localparam CM_TX_EWMA_INTERVAL_HI = 31;
localparam CM_TX_EWMA_INTERVAL_RESET = 8'h0;
localparam CM_TX_EWMA_EWMA_WHOLE_LO = 8;
localparam CM_TX_EWMA_EWMA_WHOLE_HI = 23;
localparam CM_TX_EWMA_EWMA_WHOLE_RESET = 16'h0;
localparam CM_TX_EWMA_EWMA_FRAC_LO = 0;
localparam CM_TX_EWMA_EWMA_FRAC_HI = 7;
localparam CM_TX_EWMA_EWMA_FRAC_RESET = 8'h0;
localparam CM_TX_EWMA_USEMASK = 64'hFFFFFFFF;
localparam CM_TX_EWMA_RO_MASK = 64'hFFFFFFFF;
localparam CM_TX_EWMA_WO_MASK = 64'h0;
localparam CM_TX_EWMA_RESET = 64'h0;

typedef struct packed {
    CM_GLOBAL_WM_t  CM_GLOBAL_WM;
    CM_GLOBAL_CFG_t  CM_GLOBAL_CFG;
    CM_SWEEPER_TC_TO_SMP_t  CM_SWEEPER_TC_TO_SMP;
    CM_GLOBAL_USAGE_t  CM_GLOBAL_USAGE;
    CM_GLOBAL_USAGE_MAX_t  CM_GLOBAL_USAGE_MAX;
} mby_ppe_cm_usage_map_registers_t;

// ===================================================
// load

typedef struct packed {
    logic  [0:0] COUNT;  // RW/V
} load_CM_GLOBAL_USAGE_MAX_t;

typedef struct packed {
    load_CM_GLOBAL_USAGE_MAX_t  CM_GLOBAL_USAGE_MAX;
} mby_ppe_cm_usage_map_load_t;

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

typedef struct packed {
    logic [15:0] COUNT;  // RO/V
} new_CM_GLOBAL_USAGE_t;

typedef struct packed {
    logic [15:0] COUNT;  // RW/V
} new_CM_GLOBAL_USAGE_MAX_t;

typedef struct packed {
    new_CM_GLOBAL_USAGE_t  CM_GLOBAL_USAGE;
    new_CM_GLOBAL_USAGE_MAX_t  CM_GLOBAL_USAGE_MAX;
} mby_ppe_cm_usage_map_new_t;

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_CM_TX_TC_PRIVATE_WM_t;

typedef logic [7:0] we_CM_TX_TC_HOG_WM_t;

typedef logic [7:0] we_CM_RX_SMP_PRIVATE_WM_t;

typedef logic [7:0] we_CM_RX_SMP_HOG_WM_t;

typedef logic [7:0] we_CM_RX_SMP_PAUSE_WM_t;

typedef logic [7:0] we_CM_SHARED_WM_t;

typedef logic [7:0] we_CM_SOFTDROP_WM_t;

typedef logic [7:0] we_CM_SHARED_SMP_PAUSE_WM_t;

typedef logic [7:0] we_CM_PAUSE_PHYS_PORT_CFG_t;

typedef logic [7:0] we_CM_FORCE_PAUSE_CFG_t;

typedef logic [7:0] we_CM_AQM_EWMA_CFG_t;

typedef logic [7:0] we_CM_AQM_DCTCP_CFG_t;

typedef logic [7:0] we_CM_SHARED_SMP_PAUSE_CFG_t;

typedef logic [7:0] we_CM_MCAST_EPOCH_USAGE_t;

typedef logic [7:0] we_CM_SHARED_SMP_USAGE_t;

typedef logic [7:0] we_CM_SMP_USAGE_t;

typedef logic [7:0] we_CM_RX_SMP_USAGE_t;

typedef logic [7:0] we_CM_RX_SMP_USAGE_MAX_t;

typedef logic [7:0] we_CM_RX_SMP_USAGE_MAX_CTRL_t;

typedef logic [7:0] we_CM_PAUSE_GEN_STATE_t;

typedef logic [7:0] we_CM_TX_TC_USAGE_t;

typedef logic [7:0] we_CM_TX_EWMA_t;

typedef struct packed {
    we_CM_TX_TC_PRIVATE_WM_t CM_TX_TC_PRIVATE_WM;
    we_CM_TX_TC_HOG_WM_t CM_TX_TC_HOG_WM;
    we_CM_RX_SMP_PRIVATE_WM_t CM_RX_SMP_PRIVATE_WM;
    we_CM_RX_SMP_HOG_WM_t CM_RX_SMP_HOG_WM;
    we_CM_RX_SMP_PAUSE_WM_t CM_RX_SMP_PAUSE_WM;
    we_CM_SHARED_WM_t CM_SHARED_WM;
    we_CM_SOFTDROP_WM_t CM_SOFTDROP_WM;
    we_CM_SHARED_SMP_PAUSE_WM_t CM_SHARED_SMP_PAUSE_WM;
    we_CM_PAUSE_PHYS_PORT_CFG_t CM_PAUSE_PHYS_PORT_CFG;
    we_CM_FORCE_PAUSE_CFG_t CM_FORCE_PAUSE_CFG;
    we_CM_AQM_EWMA_CFG_t CM_AQM_EWMA_CFG;
    we_CM_AQM_DCTCP_CFG_t CM_AQM_DCTCP_CFG;
    we_CM_SHARED_SMP_PAUSE_CFG_t CM_SHARED_SMP_PAUSE_CFG;
    we_CM_MCAST_EPOCH_USAGE_t CM_MCAST_EPOCH_USAGE;
    we_CM_SHARED_SMP_USAGE_t CM_SHARED_SMP_USAGE;
    we_CM_SMP_USAGE_t CM_SMP_USAGE;
    we_CM_RX_SMP_USAGE_t CM_RX_SMP_USAGE;
    we_CM_RX_SMP_USAGE_MAX_t CM_RX_SMP_USAGE_MAX;
    we_CM_RX_SMP_USAGE_MAX_CTRL_t CM_RX_SMP_USAGE_MAX_CTRL;
    we_CM_PAUSE_GEN_STATE_t CM_PAUSE_GEN_STATE;
    we_CM_TX_TC_USAGE_t CM_TX_TC_USAGE;
    we_CM_TX_EWMA_t CM_TX_EWMA;
} mby_ppe_cm_usage_map_handcoded_t;

typedef logic [7:0] re_CM_TX_TC_PRIVATE_WM_t;

typedef logic [7:0] re_CM_TX_TC_HOG_WM_t;

typedef logic [7:0] re_CM_RX_SMP_PRIVATE_WM_t;

typedef logic [7:0] re_CM_RX_SMP_HOG_WM_t;

typedef logic [7:0] re_CM_RX_SMP_PAUSE_WM_t;

typedef logic [7:0] re_CM_SHARED_WM_t;

typedef logic [7:0] re_CM_SOFTDROP_WM_t;

typedef logic [7:0] re_CM_SHARED_SMP_PAUSE_WM_t;

typedef logic [7:0] re_CM_PAUSE_PHYS_PORT_CFG_t;

typedef logic [7:0] re_CM_FORCE_PAUSE_CFG_t;

typedef logic [7:0] re_CM_AQM_EWMA_CFG_t;

typedef logic [7:0] re_CM_AQM_DCTCP_CFG_t;

typedef logic [7:0] re_CM_SHARED_SMP_PAUSE_CFG_t;

typedef logic [7:0] re_CM_MCAST_EPOCH_USAGE_t;

typedef logic [7:0] re_CM_SHARED_SMP_USAGE_t;

typedef logic [7:0] re_CM_SMP_USAGE_t;

typedef logic [7:0] re_CM_RX_SMP_USAGE_t;

typedef logic [7:0] re_CM_RX_SMP_USAGE_MAX_t;

typedef logic [7:0] re_CM_RX_SMP_USAGE_MAX_CTRL_t;

typedef logic [7:0] re_CM_PAUSE_GEN_STATE_t;

typedef logic [7:0] re_CM_TX_TC_USAGE_t;

typedef logic [7:0] re_CM_TX_EWMA_t;

typedef struct packed {
    re_CM_TX_TC_PRIVATE_WM_t CM_TX_TC_PRIVATE_WM;
    re_CM_TX_TC_HOG_WM_t CM_TX_TC_HOG_WM;
    re_CM_RX_SMP_PRIVATE_WM_t CM_RX_SMP_PRIVATE_WM;
    re_CM_RX_SMP_HOG_WM_t CM_RX_SMP_HOG_WM;
    re_CM_RX_SMP_PAUSE_WM_t CM_RX_SMP_PAUSE_WM;
    re_CM_SHARED_WM_t CM_SHARED_WM;
    re_CM_SOFTDROP_WM_t CM_SOFTDROP_WM;
    re_CM_SHARED_SMP_PAUSE_WM_t CM_SHARED_SMP_PAUSE_WM;
    re_CM_PAUSE_PHYS_PORT_CFG_t CM_PAUSE_PHYS_PORT_CFG;
    re_CM_FORCE_PAUSE_CFG_t CM_FORCE_PAUSE_CFG;
    re_CM_AQM_EWMA_CFG_t CM_AQM_EWMA_CFG;
    re_CM_AQM_DCTCP_CFG_t CM_AQM_DCTCP_CFG;
    re_CM_SHARED_SMP_PAUSE_CFG_t CM_SHARED_SMP_PAUSE_CFG;
    re_CM_MCAST_EPOCH_USAGE_t CM_MCAST_EPOCH_USAGE;
    re_CM_SHARED_SMP_USAGE_t CM_SHARED_SMP_USAGE;
    re_CM_SMP_USAGE_t CM_SMP_USAGE;
    re_CM_RX_SMP_USAGE_t CM_RX_SMP_USAGE;
    re_CM_RX_SMP_USAGE_MAX_t CM_RX_SMP_USAGE_MAX;
    re_CM_RX_SMP_USAGE_MAX_CTRL_t CM_RX_SMP_USAGE_MAX_CTRL;
    re_CM_PAUSE_GEN_STATE_t CM_PAUSE_GEN_STATE;
    re_CM_TX_TC_USAGE_t CM_TX_TC_USAGE;
    re_CM_TX_EWMA_t CM_TX_EWMA;
} mby_ppe_cm_usage_map_hc_re_t;

typedef logic handcode_rvalid_CM_TX_TC_PRIVATE_WM_t;

typedef logic handcode_rvalid_CM_TX_TC_HOG_WM_t;

typedef logic handcode_rvalid_CM_RX_SMP_PRIVATE_WM_t;

typedef logic handcode_rvalid_CM_RX_SMP_HOG_WM_t;

typedef logic handcode_rvalid_CM_RX_SMP_PAUSE_WM_t;

typedef logic handcode_rvalid_CM_SHARED_WM_t;

typedef logic handcode_rvalid_CM_SOFTDROP_WM_t;

typedef logic handcode_rvalid_CM_SHARED_SMP_PAUSE_WM_t;

typedef logic handcode_rvalid_CM_PAUSE_PHYS_PORT_CFG_t;

typedef logic handcode_rvalid_CM_FORCE_PAUSE_CFG_t;

typedef logic handcode_rvalid_CM_AQM_EWMA_CFG_t;

typedef logic handcode_rvalid_CM_AQM_DCTCP_CFG_t;

typedef logic handcode_rvalid_CM_SHARED_SMP_PAUSE_CFG_t;

typedef logic handcode_rvalid_CM_MCAST_EPOCH_USAGE_t;

typedef logic handcode_rvalid_CM_SHARED_SMP_USAGE_t;

typedef logic handcode_rvalid_CM_SMP_USAGE_t;

typedef logic handcode_rvalid_CM_RX_SMP_USAGE_t;

typedef logic handcode_rvalid_CM_RX_SMP_USAGE_MAX_t;

typedef logic handcode_rvalid_CM_RX_SMP_USAGE_MAX_CTRL_t;

typedef logic handcode_rvalid_CM_PAUSE_GEN_STATE_t;

typedef logic handcode_rvalid_CM_TX_TC_USAGE_t;

typedef logic handcode_rvalid_CM_TX_EWMA_t;

typedef struct packed {
    handcode_rvalid_CM_TX_TC_PRIVATE_WM_t CM_TX_TC_PRIVATE_WM;
    handcode_rvalid_CM_TX_TC_HOG_WM_t CM_TX_TC_HOG_WM;
    handcode_rvalid_CM_RX_SMP_PRIVATE_WM_t CM_RX_SMP_PRIVATE_WM;
    handcode_rvalid_CM_RX_SMP_HOG_WM_t CM_RX_SMP_HOG_WM;
    handcode_rvalid_CM_RX_SMP_PAUSE_WM_t CM_RX_SMP_PAUSE_WM;
    handcode_rvalid_CM_SHARED_WM_t CM_SHARED_WM;
    handcode_rvalid_CM_SOFTDROP_WM_t CM_SOFTDROP_WM;
    handcode_rvalid_CM_SHARED_SMP_PAUSE_WM_t CM_SHARED_SMP_PAUSE_WM;
    handcode_rvalid_CM_PAUSE_PHYS_PORT_CFG_t CM_PAUSE_PHYS_PORT_CFG;
    handcode_rvalid_CM_FORCE_PAUSE_CFG_t CM_FORCE_PAUSE_CFG;
    handcode_rvalid_CM_AQM_EWMA_CFG_t CM_AQM_EWMA_CFG;
    handcode_rvalid_CM_AQM_DCTCP_CFG_t CM_AQM_DCTCP_CFG;
    handcode_rvalid_CM_SHARED_SMP_PAUSE_CFG_t CM_SHARED_SMP_PAUSE_CFG;
    handcode_rvalid_CM_MCAST_EPOCH_USAGE_t CM_MCAST_EPOCH_USAGE;
    handcode_rvalid_CM_SHARED_SMP_USAGE_t CM_SHARED_SMP_USAGE;
    handcode_rvalid_CM_SMP_USAGE_t CM_SMP_USAGE;
    handcode_rvalid_CM_RX_SMP_USAGE_t CM_RX_SMP_USAGE;
    handcode_rvalid_CM_RX_SMP_USAGE_MAX_t CM_RX_SMP_USAGE_MAX;
    handcode_rvalid_CM_RX_SMP_USAGE_MAX_CTRL_t CM_RX_SMP_USAGE_MAX_CTRL;
    handcode_rvalid_CM_PAUSE_GEN_STATE_t CM_PAUSE_GEN_STATE;
    handcode_rvalid_CM_TX_TC_USAGE_t CM_TX_TC_USAGE;
    handcode_rvalid_CM_TX_EWMA_t CM_TX_EWMA;
} mby_ppe_cm_usage_map_hc_rvalid_t;

typedef logic handcode_wvalid_CM_TX_TC_PRIVATE_WM_t;

typedef logic handcode_wvalid_CM_TX_TC_HOG_WM_t;

typedef logic handcode_wvalid_CM_RX_SMP_PRIVATE_WM_t;

typedef logic handcode_wvalid_CM_RX_SMP_HOG_WM_t;

typedef logic handcode_wvalid_CM_RX_SMP_PAUSE_WM_t;

typedef logic handcode_wvalid_CM_SHARED_WM_t;

typedef logic handcode_wvalid_CM_SOFTDROP_WM_t;

typedef logic handcode_wvalid_CM_SHARED_SMP_PAUSE_WM_t;

typedef logic handcode_wvalid_CM_PAUSE_PHYS_PORT_CFG_t;

typedef logic handcode_wvalid_CM_FORCE_PAUSE_CFG_t;

typedef logic handcode_wvalid_CM_AQM_EWMA_CFG_t;

typedef logic handcode_wvalid_CM_AQM_DCTCP_CFG_t;

typedef logic handcode_wvalid_CM_SHARED_SMP_PAUSE_CFG_t;

typedef logic handcode_wvalid_CM_MCAST_EPOCH_USAGE_t;

typedef logic handcode_wvalid_CM_SHARED_SMP_USAGE_t;

typedef logic handcode_wvalid_CM_SMP_USAGE_t;

typedef logic handcode_wvalid_CM_RX_SMP_USAGE_t;

typedef logic handcode_wvalid_CM_RX_SMP_USAGE_MAX_t;

typedef logic handcode_wvalid_CM_RX_SMP_USAGE_MAX_CTRL_t;

typedef logic handcode_wvalid_CM_PAUSE_GEN_STATE_t;

typedef logic handcode_wvalid_CM_TX_TC_USAGE_t;

typedef logic handcode_wvalid_CM_TX_EWMA_t;

typedef struct packed {
    handcode_wvalid_CM_TX_TC_PRIVATE_WM_t CM_TX_TC_PRIVATE_WM;
    handcode_wvalid_CM_TX_TC_HOG_WM_t CM_TX_TC_HOG_WM;
    handcode_wvalid_CM_RX_SMP_PRIVATE_WM_t CM_RX_SMP_PRIVATE_WM;
    handcode_wvalid_CM_RX_SMP_HOG_WM_t CM_RX_SMP_HOG_WM;
    handcode_wvalid_CM_RX_SMP_PAUSE_WM_t CM_RX_SMP_PAUSE_WM;
    handcode_wvalid_CM_SHARED_WM_t CM_SHARED_WM;
    handcode_wvalid_CM_SOFTDROP_WM_t CM_SOFTDROP_WM;
    handcode_wvalid_CM_SHARED_SMP_PAUSE_WM_t CM_SHARED_SMP_PAUSE_WM;
    handcode_wvalid_CM_PAUSE_PHYS_PORT_CFG_t CM_PAUSE_PHYS_PORT_CFG;
    handcode_wvalid_CM_FORCE_PAUSE_CFG_t CM_FORCE_PAUSE_CFG;
    handcode_wvalid_CM_AQM_EWMA_CFG_t CM_AQM_EWMA_CFG;
    handcode_wvalid_CM_AQM_DCTCP_CFG_t CM_AQM_DCTCP_CFG;
    handcode_wvalid_CM_SHARED_SMP_PAUSE_CFG_t CM_SHARED_SMP_PAUSE_CFG;
    handcode_wvalid_CM_MCAST_EPOCH_USAGE_t CM_MCAST_EPOCH_USAGE;
    handcode_wvalid_CM_SHARED_SMP_USAGE_t CM_SHARED_SMP_USAGE;
    handcode_wvalid_CM_SMP_USAGE_t CM_SMP_USAGE;
    handcode_wvalid_CM_RX_SMP_USAGE_t CM_RX_SMP_USAGE;
    handcode_wvalid_CM_RX_SMP_USAGE_MAX_t CM_RX_SMP_USAGE_MAX;
    handcode_wvalid_CM_RX_SMP_USAGE_MAX_CTRL_t CM_RX_SMP_USAGE_MAX_CTRL;
    handcode_wvalid_CM_PAUSE_GEN_STATE_t CM_PAUSE_GEN_STATE;
    handcode_wvalid_CM_TX_TC_USAGE_t CM_TX_TC_USAGE;
    handcode_wvalid_CM_TX_EWMA_t CM_TX_EWMA;
} mby_ppe_cm_usage_map_hc_wvalid_t;

typedef logic handcode_error_CM_TX_TC_PRIVATE_WM_t;

typedef logic handcode_error_CM_TX_TC_HOG_WM_t;

typedef logic handcode_error_CM_RX_SMP_PRIVATE_WM_t;

typedef logic handcode_error_CM_RX_SMP_HOG_WM_t;

typedef logic handcode_error_CM_RX_SMP_PAUSE_WM_t;

typedef logic handcode_error_CM_SHARED_WM_t;

typedef logic handcode_error_CM_SOFTDROP_WM_t;

typedef logic handcode_error_CM_SHARED_SMP_PAUSE_WM_t;

typedef logic handcode_error_CM_PAUSE_PHYS_PORT_CFG_t;

typedef logic handcode_error_CM_FORCE_PAUSE_CFG_t;

typedef logic handcode_error_CM_AQM_EWMA_CFG_t;

typedef logic handcode_error_CM_AQM_DCTCP_CFG_t;

typedef logic handcode_error_CM_SHARED_SMP_PAUSE_CFG_t;

typedef logic handcode_error_CM_MCAST_EPOCH_USAGE_t;

typedef logic handcode_error_CM_SHARED_SMP_USAGE_t;

typedef logic handcode_error_CM_SMP_USAGE_t;

typedef logic handcode_error_CM_RX_SMP_USAGE_t;

typedef logic handcode_error_CM_RX_SMP_USAGE_MAX_t;

typedef logic handcode_error_CM_RX_SMP_USAGE_MAX_CTRL_t;

typedef logic handcode_error_CM_PAUSE_GEN_STATE_t;

typedef logic handcode_error_CM_TX_TC_USAGE_t;

typedef logic handcode_error_CM_TX_EWMA_t;

typedef struct packed {
    handcode_error_CM_TX_TC_PRIVATE_WM_t CM_TX_TC_PRIVATE_WM;
    handcode_error_CM_TX_TC_HOG_WM_t CM_TX_TC_HOG_WM;
    handcode_error_CM_RX_SMP_PRIVATE_WM_t CM_RX_SMP_PRIVATE_WM;
    handcode_error_CM_RX_SMP_HOG_WM_t CM_RX_SMP_HOG_WM;
    handcode_error_CM_RX_SMP_PAUSE_WM_t CM_RX_SMP_PAUSE_WM;
    handcode_error_CM_SHARED_WM_t CM_SHARED_WM;
    handcode_error_CM_SOFTDROP_WM_t CM_SOFTDROP_WM;
    handcode_error_CM_SHARED_SMP_PAUSE_WM_t CM_SHARED_SMP_PAUSE_WM;
    handcode_error_CM_PAUSE_PHYS_PORT_CFG_t CM_PAUSE_PHYS_PORT_CFG;
    handcode_error_CM_FORCE_PAUSE_CFG_t CM_FORCE_PAUSE_CFG;
    handcode_error_CM_AQM_EWMA_CFG_t CM_AQM_EWMA_CFG;
    handcode_error_CM_AQM_DCTCP_CFG_t CM_AQM_DCTCP_CFG;
    handcode_error_CM_SHARED_SMP_PAUSE_CFG_t CM_SHARED_SMP_PAUSE_CFG;
    handcode_error_CM_MCAST_EPOCH_USAGE_t CM_MCAST_EPOCH_USAGE;
    handcode_error_CM_SHARED_SMP_USAGE_t CM_SHARED_SMP_USAGE;
    handcode_error_CM_SMP_USAGE_t CM_SMP_USAGE;
    handcode_error_CM_RX_SMP_USAGE_t CM_RX_SMP_USAGE;
    handcode_error_CM_RX_SMP_USAGE_MAX_t CM_RX_SMP_USAGE_MAX;
    handcode_error_CM_RX_SMP_USAGE_MAX_CTRL_t CM_RX_SMP_USAGE_MAX_CTRL;
    handcode_error_CM_PAUSE_GEN_STATE_t CM_PAUSE_GEN_STATE;
    handcode_error_CM_TX_TC_USAGE_t CM_TX_TC_USAGE;
    handcode_error_CM_TX_EWMA_t CM_TX_EWMA;
} mby_ppe_cm_usage_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    CM_TX_TC_PRIVATE_WM_t CM_TX_TC_PRIVATE_WM;
    CM_TX_TC_HOG_WM_t CM_TX_TC_HOG_WM;
    CM_RX_SMP_PRIVATE_WM_t CM_RX_SMP_PRIVATE_WM;
    CM_RX_SMP_HOG_WM_t CM_RX_SMP_HOG_WM;
    CM_RX_SMP_PAUSE_WM_t CM_RX_SMP_PAUSE_WM;
    CM_SHARED_WM_t CM_SHARED_WM;
    CM_SOFTDROP_WM_t CM_SOFTDROP_WM;
    CM_SHARED_SMP_PAUSE_WM_t CM_SHARED_SMP_PAUSE_WM;
    CM_PAUSE_PHYS_PORT_CFG_t CM_PAUSE_PHYS_PORT_CFG;
    CM_FORCE_PAUSE_CFG_t CM_FORCE_PAUSE_CFG;
    CM_AQM_EWMA_CFG_t CM_AQM_EWMA_CFG;
    CM_AQM_DCTCP_CFG_t CM_AQM_DCTCP_CFG;
    CM_SHARED_SMP_PAUSE_CFG_t CM_SHARED_SMP_PAUSE_CFG;
    CM_MCAST_EPOCH_USAGE_t CM_MCAST_EPOCH_USAGE;
    CM_SHARED_SMP_USAGE_t CM_SHARED_SMP_USAGE;
    CM_SMP_USAGE_t CM_SMP_USAGE;
    CM_RX_SMP_USAGE_t CM_RX_SMP_USAGE;
    CM_RX_SMP_USAGE_MAX_t CM_RX_SMP_USAGE_MAX;
    CM_RX_SMP_USAGE_MAX_CTRL_t CM_RX_SMP_USAGE_MAX_CTRL;
    CM_PAUSE_GEN_STATE_t CM_PAUSE_GEN_STATE;
    CM_TX_TC_USAGE_t CM_TX_TC_USAGE;
    CM_TX_EWMA_t CM_TX_EWMA;
} mby_ppe_cm_usage_map_hc_reg_read_t;

typedef struct packed {
    CM_TX_TC_PRIVATE_WM_t CM_TX_TC_PRIVATE_WM;
    CM_TX_TC_HOG_WM_t CM_TX_TC_HOG_WM;
    CM_RX_SMP_PRIVATE_WM_t CM_RX_SMP_PRIVATE_WM;
    CM_RX_SMP_HOG_WM_t CM_RX_SMP_HOG_WM;
    CM_RX_SMP_PAUSE_WM_t CM_RX_SMP_PAUSE_WM;
    CM_SHARED_WM_t CM_SHARED_WM;
    CM_SOFTDROP_WM_t CM_SOFTDROP_WM;
    CM_SHARED_SMP_PAUSE_WM_t CM_SHARED_SMP_PAUSE_WM;
    CM_PAUSE_PHYS_PORT_CFG_t CM_PAUSE_PHYS_PORT_CFG;
    CM_FORCE_PAUSE_CFG_t CM_FORCE_PAUSE_CFG;
    CM_AQM_EWMA_CFG_t CM_AQM_EWMA_CFG;
    CM_AQM_DCTCP_CFG_t CM_AQM_DCTCP_CFG;
    CM_SHARED_SMP_PAUSE_CFG_t CM_SHARED_SMP_PAUSE_CFG;
    CM_MCAST_EPOCH_USAGE_t CM_MCAST_EPOCH_USAGE;
    CM_SHARED_SMP_USAGE_t CM_SHARED_SMP_USAGE;
    CM_SMP_USAGE_t CM_SMP_USAGE;
    CM_RX_SMP_USAGE_t CM_RX_SMP_USAGE;
    CM_RX_SMP_USAGE_MAX_t CM_RX_SMP_USAGE_MAX;
    CM_RX_SMP_USAGE_MAX_CTRL_t CM_RX_SMP_USAGE_MAX_CTRL;
    CM_PAUSE_GEN_STATE_t CM_PAUSE_GEN_STATE;
    CM_TX_TC_USAGE_t CM_TX_TC_USAGE;
    CM_TX_EWMA_t CM_TX_EWMA;
} mby_ppe_cm_usage_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_cm_usage_map_pkg

`endif // MBY_PPE_CM_USAGE_MAP_PKG_VH
