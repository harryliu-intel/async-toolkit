//-----------------------------------------------------------------------------
// Title         : Madison Bay Base Package
// Project       : Madison Bay
//-----------------------------------------------------------------------------
// File          : mby_base_pkg.svh
// Author        : jose.j.godinez.carrillo  <jjgodine@ichips.intel.com>
// Created       : 29.10.2018
//-----------------------------------------------------------------------------
// Description :
// This is the base sequencer class for Madison Bay
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by Intel Corporation This model is the confidential and
// proprietary property of Intel Corporation and the possession or use of this
// file requires a written license from Intel Corporation.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors. The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
`ifndef __MBY_BASE_PKG__
`define __MBY_BASE_PKG__
//------------------------------------------------------------------------------
//
// PACKAGE: mby_base_pkg
// This is the Madison Bay base agent package, currently it depends on the uvm,
// and shdv_base_pkg verification packages. It defines a base agent, which
// is a parameterized class that can be used to create simple agents quickly.
// Image:
//    (see ./mby_base_pkg.png)
//
//------------------------------------------------------------------------------
package mby_base_pkg;

   import uvm_pkg::*;
   import shdv_base_pkg::*;

   `include "uvm_macros.svh"
   `include "mby_base_config.svh"
   `include "mby_base_sequence_item.svh"
   `include "mby_base_sequence_item_param.svh"
   `include "mby_base_flow_control.svh"
   `include "mby_base_io_policy.svh"
   `include "mby_base_io_policy_param.svh"
   `include "mby_base_sequencer.svh"
   `include "mby_base_monitor.svh"
   `include "mby_base_driver.svh"
   `include "mby_base_agent.svh"

endpackage

`endif
