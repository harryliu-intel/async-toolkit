///
///  INTEL CONFIDENTIAL
///
///  Copyright 2019 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_rx_pb.sv                                               
// Creator:         edwardro                                                   
// Time:            Wednesday Jan 23, 2019 [5:27:04 am]                        
//                                                                             
// Path:            /tmp/edwardro/nebulon_run/211708214340_2019-01-23.05:26:34 
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1130/edwardro/mby/work_root/mby.edr.pbb/tools/srdl
//                  -sv_no_sai_checks -sverilog -crif -expand_handcoded_arrays 
//                  -maximize_crif -input mby_rx_pb_map.rdl -timeout 60000     
//                  -out_dir /tmp/tmp.QONdsBBv97 -log_file                     
//                  /nfs/site/disks/slx_1130/edwardro/mby/work_root/mby.edr.pbb/target/GenRTL/regflow/mby/subblock/mby_rx_pb_map_crif.xml.log
//                                                                             
// MRE:             5.2018.3.p1                                                
// Machine:         sccj019434                                                 
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww52.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2019 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww52.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_rx_pb_map.vh"
`include "rtlgen_pkg_mby_rx_pb_map.vh"
`include "mby_rx_pb_pkg.vh"

//lintra push -68094

// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_RX_PB_FF
`define RTLGEN_MBY_RX_PB_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_RX_PB_FF

`ifndef RTLGEN_MBY_RX_PB_EN_FF
`define RTLGEN_MBY_RX_PB_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_RX_PB_EN_FF

`ifndef RTLGEN_MBY_RX_PB_FF_RSTD
`define RTLGEN_MBY_RX_PB_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_RX_PB_FF_RSTD


module rtlgen_mby_rx_pb_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_RX_PB_EN_FF_RSTD
`define RTLGEN_MBY_RX_PB_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_rx_pb_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_RX_PB_EN_FF_RSTD


`ifndef RTLGEN_MBY_RX_PB_FF_SYNCRST
`define RTLGEN_MBY_RX_PB_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_RX_PB_FF_SYNCRST

`ifndef RTLGEN_MBY_RX_PB_EN_FF_SYNCRST
`define RTLGEN_MBY_RX_PB_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_RX_PB_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_RX_PB_FF_BOTHRST
// `define RTLGEN_MBY_RX_PB_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_RX_PB_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_RX_PB_EN_FF_BOTHRST
// `define RTLGEN_MBY_RX_PB_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_RX_PB_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_RX_PB_LATCH_LOW
`define RTLGEN_MBY_RX_PB_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_RX_PB_LATCH_LOW

`ifndef RTLGEN_MBY_RX_PB_PH2_FF
`define RTLGEN_MBY_RX_PB_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) \
     q <= d;
`endif // RTLGEN_MBY_RX_PB_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_RX_PB_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_RX_PB_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_RX_PB_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_RX_PB_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_RX_PB_PH2_FF_ASSIGN
`define RTLGEN_MBY_RX_PB_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_RX_PB_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_RX_PB_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_RX_PB_LATCH
`define RTLGEN_MBY_RX_PB_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_RX_PB_LATCH

`ifndef RTLGEN_MBY_RX_PB_EN_LATCH
`define RTLGEN_MBY_RX_PB_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_RX_PB_EN_LATCH

`ifndef RTLGEN_MBY_RX_PB_EN_LATCH_LOW
`define RTLGEN_MBY_RX_PB_EN_LATCH_LOW(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_RX_PB_EN_LATCH_LOW

`ifndef RTLGEN_MBY_RX_PB_LATCH_SYNCRST
`define RTLGEN_MBY_RX_PB_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_RX_PB_LATCH_SYNCRST

`ifndef RTLGEN_MBY_RX_PB_EN_LATCH_SYNCRST
`define RTLGEN_MBY_RX_PB_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_RX_PB_EN_LATCH_SYNCRST

`ifndef RTLGEN_MBY_RX_PB_EN_LATCH_LOW_SYNCRST
`define RTLGEN_MBY_RX_PB_EN_LATCH_LOW_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_RX_PB_EN_LATCH_LOW_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_RX_PB_LATCH_BOTHRST
// `define RTLGEN_MBY_RX_PB_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_RX_PB_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_RX_PB_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_RX_PB_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_RX_PB_EN_LATCH_BOTHRST


// ===================================================================
// LCB macros 
// ===================================================================

`ifndef RTLGEN_MBY_RX_PB_LCB_HOLD_REQ_2CYCLES
`define RTLGEN_MBY_RX_PB_LCB_HOLD_REQ_2CYCLES(clock, enable, lcb_clk) \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & enable;
`endif // RTLGEN_MBY_RX_PB_LCB_HOLD_REQ_2CYCLES

`ifndef RTLGEN_MBY_RX_PB_LCB_HOLD_REQ_2CYCLES_SYNCRST
`define RTLGEN_MBY_RX_PB_LCB_HOLD_REQ_2CYCLES_SYNCRST(clock, enable, lcb_clk, sync_rst) \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & (enable | {$bits(lcb_clk){!sync_rst}});
`endif // RTLGEN_MBY_RX_PB_LCB_HOLD_REQ_2CYCLES_SYNCRST

`ifndef RTLGEN_MBY_RX_PB_LCB_DELAY
`define RTLGEN_MBY_RX_PB_LCB_DELAY(clock, delay_rst_n, enable, lcb_clk, seq_type, nxt_expr) \
   logic [$bits(lcb_clk)-1:0] ``enable``_up;  \
   logic [$bits(lcb_clk)-1:0] ``enable``_nxt; \
   logic [$bits(lcb_clk)-1:0] ``enable``_dly; \
   always_comb ``enable``_nxt = ``nxt_expr``; \
   always_comb ``enable``_up = ``enable``_nxt | ``enable``_dly; \
   genvar ``enable``_gen_var ; \
   generate \
      if (1) begin : rtlgen_lcb_``enable``_dly \
         for ( ``enable``_gen_var = 0 ; ``enable``_gen_var < $bits(lcb_clk); ``enable``_gen_var = ``enable``_gen_var + 1) \
  `RTLGEN_MBY_RX_PB_``seq_type``(clock,delay_rst_n,1'b0,``enable``_up[ ``enable``_gen_var ],``enable``_nxt[ ``enable``_gen_var ],``enable``_dly[ ``enable``_gen_var ]) \
      end      \
   endgenerate \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & ``enable``_dly;
`endif // RTLGEN_MBY_RX_PB_LCB_DELAY

`ifndef RTLGEN_MBY_RX_PB_LCB_LATCH_LOW_PHASE
`define RTLGEN_MBY_RX_PB_LCB_LATCH_LOW_PHASE(clock, delay_rst_n, enable, lcb_clk) \
   `RTLGEN_MBY_RX_PB_LCB_DELAY(clock,delay_rst_n,enable,lcb_clk,EN_LATCH_LOW,enable)
`endif // RTLGEN_MBY_RX_PB_LCB_LATCH_LOW_PHASE

`ifndef RTLGEN_MBY_RX_PB_LCB_LATCH_LOW_PHASE_SYNCRST
`define RTLGEN_MBY_RX_PB_LCB_LATCH_LOW_PHASE_SYNCRST(clock, delay_rst_n, enable, lcb_clk, sync_rst) \
   `RTLGEN_MBY_RX_PB_LCB_DELAY(clock,1'b1,enable,lcb_clk,EN_LATCH_LOW_SYNCRST,enable|{$bits(lcb_clk){!sync_rst}})
`endif // RTLGEN_MBY_RX_PB_LCB_LATCH_LOW_PHASE_SYNCRST

`ifndef RTLGEN_MBY_RX_PB_LCB_FF_POSEDGE
`define RTLGEN_MBY_RX_PB_LCB_FF_POSEDGE(clock, delay_rst_n, enable, lcb_clk)  \
   `RTLGEN_MBY_RX_PB_LCB_DELAY(clock,delay_rst_n,enable,lcb_clk,EN_FF,enable)
`endif // RTLGEN_MBY_RX_PB_LCB_FF_POSEDGE

`ifndef RTLGEN_MBY_RX_PB_LCB_FF_POSEDGE_SYNCRST
`define RTLGEN_MBY_RX_PB_LCB_FF_POSEDGE_SYNCRST(clock, delay_rst_n, enable, lcb_clk, sync_rst) \
   `RTLGEN_MBY_RX_PB_LCB_DELAY(clock,1'b1,enable,lcb_clk,EN_FF_SYNCRST,enable|{$bits(lcb_clk){!sync_rst}})
`endif // RTLGEN_MBY_RX_PB_LCB_FF_POSEDGE_SYNCRST



//lintra pop

module mby_rx_pb ( //lintra s-2096
    // Clocks
    gated_clk,

    // Resets
    rst_n,


    // Register Inputs


    // Register Outputs
    RX_PB_PORT_CFG,
    RX_PB_WM,


    // Register signals for HandCoded registers



    // Config Access
    req,
    ack
    

);

import mby_rx_pb_pkg::*;
import rtlgen_pkg_mby_rx_pb_map::*;

parameter  MBY_RX_PB_MEM_ADDR_MSB = 47;
parameter [MBY_RX_PB_MEM_ADDR_MSB:0] MBY_RX_PB_MAP_OFFSET = {MBY_RX_PB_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] MBY_RX_PB_MAP_SB_BAR = 3'b0;
parameter [7:0] MBY_RX_PB_MAP_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
`define RX_PB_WM_CR_ADDR_def(INDEX) RX_PB_WM_CR_ADDR``INDEX``[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_RX_PB_MAP_OFFSET[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
localparam [MBY_RX_PB_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] RX_PB_PORT_CFG_DECODE_ADDR = RX_PB_PORT_CFG_CR_ADDR[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_RX_PB_MAP_OFFSET[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [16:0][7:0][MBY_RX_PB_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] RX_PB_WM_DECODE_ADDR = {{`RX_PB_WM_CR_ADDR_def([16][7]),`RX_PB_WM_CR_ADDR_def([16][6]),`RX_PB_WM_CR_ADDR_def([16][5]),`RX_PB_WM_CR_ADDR_def([16][4]),`RX_PB_WM_CR_ADDR_def([16][3]),`RX_PB_WM_CR_ADDR_def([16][2]),`RX_PB_WM_CR_ADDR_def([16][1]),`RX_PB_WM_CR_ADDR_def([16][0])},{`RX_PB_WM_CR_ADDR_def([15][7]),`RX_PB_WM_CR_ADDR_def([15][6]),`RX_PB_WM_CR_ADDR_def([15][5]),`RX_PB_WM_CR_ADDR_def([15][4]),`RX_PB_WM_CR_ADDR_def([15][3]),`RX_PB_WM_CR_ADDR_def([15][2]),`RX_PB_WM_CR_ADDR_def([15][1]),`RX_PB_WM_CR_ADDR_def([15][0])},{`RX_PB_WM_CR_ADDR_def([14][7]),`RX_PB_WM_CR_ADDR_def([14][6]),`RX_PB_WM_CR_ADDR_def([14][5]),`RX_PB_WM_CR_ADDR_def([14][4]),`RX_PB_WM_CR_ADDR_def([14][3]),`RX_PB_WM_CR_ADDR_def([14][2]),`RX_PB_WM_CR_ADDR_def([14][1]),`RX_PB_WM_CR_ADDR_def([14][0])},{`RX_PB_WM_CR_ADDR_def([13][7]),`RX_PB_WM_CR_ADDR_def([13][6]),`RX_PB_WM_CR_ADDR_def([13][5]),`RX_PB_WM_CR_ADDR_def([13][4]),`RX_PB_WM_CR_ADDR_def([13][3]),`RX_PB_WM_CR_ADDR_def([13][2]),`RX_PB_WM_CR_ADDR_def([13][1]),`RX_PB_WM_CR_ADDR_def([13][0])},{`RX_PB_WM_CR_ADDR_def([12][7]),`RX_PB_WM_CR_ADDR_def([12][6]),`RX_PB_WM_CR_ADDR_def([12][5]),`RX_PB_WM_CR_ADDR_def([12][4]),`RX_PB_WM_CR_ADDR_def([12][3]),`RX_PB_WM_CR_ADDR_def([12][2]),`RX_PB_WM_CR_ADDR_def([12][1]),`RX_PB_WM_CR_ADDR_def([12][0])},{`RX_PB_WM_CR_ADDR_def([11][7]),`RX_PB_WM_CR_ADDR_def([11][6]),`RX_PB_WM_CR_ADDR_def([11][5]),`RX_PB_WM_CR_ADDR_def([11][4]),`RX_PB_WM_CR_ADDR_def([11][3]),`RX_PB_WM_CR_ADDR_def([11][2]),`RX_PB_WM_CR_ADDR_def([11][1]),`RX_PB_WM_CR_ADDR_def([11][0])},{`RX_PB_WM_CR_ADDR_def([10][7]),`RX_PB_WM_CR_ADDR_def([10][6]),`RX_PB_WM_CR_ADDR_def([10][5]),`RX_PB_WM_CR_ADDR_def([10][4]),`RX_PB_WM_CR_ADDR_def([10][3]),`RX_PB_WM_CR_ADDR_def([10][2]),`RX_PB_WM_CR_ADDR_def([10][1]),`RX_PB_WM_CR_ADDR_def([10][0])},{`RX_PB_WM_CR_ADDR_def([9][7]),`RX_PB_WM_CR_ADDR_def([9][6]),`RX_PB_WM_CR_ADDR_def([9][5]),`RX_PB_WM_CR_ADDR_def([9][4]),`RX_PB_WM_CR_ADDR_def([9][3]),`RX_PB_WM_CR_ADDR_def([9][2]),`RX_PB_WM_CR_ADDR_def([9][1]),`RX_PB_WM_CR_ADDR_def([9][0])},{`RX_PB_WM_CR_ADDR_def([8][7]),`RX_PB_WM_CR_ADDR_def([8][6]),`RX_PB_WM_CR_ADDR_def([8][5]),`RX_PB_WM_CR_ADDR_def([8][4]),`RX_PB_WM_CR_ADDR_def([8][3]),`RX_PB_WM_CR_ADDR_def([8][2]),`RX_PB_WM_CR_ADDR_def([8][1]),`RX_PB_WM_CR_ADDR_def([8][0])},{`RX_PB_WM_CR_ADDR_def([7][7]),`RX_PB_WM_CR_ADDR_def([7][6]),`RX_PB_WM_CR_ADDR_def([7][5]),`RX_PB_WM_CR_ADDR_def([7][4]),`RX_PB_WM_CR_ADDR_def([7][3]),`RX_PB_WM_CR_ADDR_def([7][2]),`RX_PB_WM_CR_ADDR_def([7][1]),`RX_PB_WM_CR_ADDR_def([7][0])},{`RX_PB_WM_CR_ADDR_def([6][7]),`RX_PB_WM_CR_ADDR_def([6][6]),`RX_PB_WM_CR_ADDR_def([6][5]),`RX_PB_WM_CR_ADDR_def([6][4]),`RX_PB_WM_CR_ADDR_def([6][3]),`RX_PB_WM_CR_ADDR_def([6][2]),`RX_PB_WM_CR_ADDR_def([6][1]),`RX_PB_WM_CR_ADDR_def([6][0])},{`RX_PB_WM_CR_ADDR_def([5][7]),`RX_PB_WM_CR_ADDR_def([5][6]),`RX_PB_WM_CR_ADDR_def([5][5]),`RX_PB_WM_CR_ADDR_def([5][4]),`RX_PB_WM_CR_ADDR_def([5][3]),`RX_PB_WM_CR_ADDR_def([5][2]),`RX_PB_WM_CR_ADDR_def([5][1]),`RX_PB_WM_CR_ADDR_def([5][0])},{`RX_PB_WM_CR_ADDR_def([4][7]),`RX_PB_WM_CR_ADDR_def([4][6]),`RX_PB_WM_CR_ADDR_def([4][5]),`RX_PB_WM_CR_ADDR_def([4][4]),`RX_PB_WM_CR_ADDR_def([4][3]),`RX_PB_WM_CR_ADDR_def([4][2]),`RX_PB_WM_CR_ADDR_def([4][1]),`RX_PB_WM_CR_ADDR_def([4][0])},{`RX_PB_WM_CR_ADDR_def([3][7]),`RX_PB_WM_CR_ADDR_def([3][6]),`RX_PB_WM_CR_ADDR_def([3][5]),`RX_PB_WM_CR_ADDR_def([3][4]),`RX_PB_WM_CR_ADDR_def([3][3]),`RX_PB_WM_CR_ADDR_def([3][2]),`RX_PB_WM_CR_ADDR_def([3][1]),`RX_PB_WM_CR_ADDR_def([3][0])},{`RX_PB_WM_CR_ADDR_def([2][7]),`RX_PB_WM_CR_ADDR_def([2][6]),`RX_PB_WM_CR_ADDR_def([2][5]),`RX_PB_WM_CR_ADDR_def([2][4]),`RX_PB_WM_CR_ADDR_def([2][3]),`RX_PB_WM_CR_ADDR_def([2][2]),`RX_PB_WM_CR_ADDR_def([2][1]),`RX_PB_WM_CR_ADDR_def([2][0])},{`RX_PB_WM_CR_ADDR_def([1][7]),`RX_PB_WM_CR_ADDR_def([1][6]),`RX_PB_WM_CR_ADDR_def([1][5]),`RX_PB_WM_CR_ADDR_def([1][4]),`RX_PB_WM_CR_ADDR_def([1][3]),`RX_PB_WM_CR_ADDR_def([1][2]),`RX_PB_WM_CR_ADDR_def([1][1]),`RX_PB_WM_CR_ADDR_def([1][0])},{`RX_PB_WM_CR_ADDR_def([0][7]),`RX_PB_WM_CR_ADDR_def([0][6]),`RX_PB_WM_CR_ADDR_def([0][5]),`RX_PB_WM_CR_ADDR_def([0][4]),`RX_PB_WM_CR_ADDR_def([0][3]),`RX_PB_WM_CR_ADDR_def([0][2]),`RX_PB_WM_CR_ADDR_def([0][1]),`RX_PB_WM_CR_ADDR_def([0][0])}};

    // Clocks
input logic  gated_clk;

    // Resets
input logic  rst_n;


    // Register Inputs


    // Register Outputs
output RX_PB_PORT_CFG_t  RX_PB_PORT_CFG;
output RX_PB_WM_t [16:0][7:0] RX_PB_WM;


    // Register signals for HandCoded registers



    // Config Access
input mby_rx_pb_cr_req_t  req;
output mby_rx_pb_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_rx_pb_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode

// Shared registers definitions





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_RX_PB_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_RX_PB_MEM;
assign case_req_addr_MBY_RX_PB_MEM = req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_mby_rx_pb_map;
always_comb begin : sb_fid_cond_mby_rx_pb_map_BLOCK
    unique casez (req_fid) 
		MBY_RX_PB_MAP_SB_FID: sb_fid_cond_mby_rx_pb_map = 1;
		default: sb_fid_cond_mby_rx_pb_map = 0;
    endcase 
end


logic sb_bar_cond_mby_rx_pb_map;
always_comb begin : sb_bar_cond_mby_rx_pb_map_BLOCK
    unique casez (req_bar) 
		MBY_RX_PB_MAP_SB_BAR: sb_bar_cond_mby_rx_pb_map = 1;
		default: sb_bar_cond_mby_rx_pb_map = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

//---------------------------------------------------------------------
// RX_PB_PORT_CFG Address Decode
logic  addr_decode_RX_PB_PORT_CFG;
logic  write_req_RX_PB_PORT_CFG;
always_comb begin
   addr_decode_RX_PB_PORT_CFG = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_PORT_CFG_DECODE_ADDR) && req.valid ;
   write_req_RX_PB_PORT_CFG = IsMEMWr && addr_decode_RX_PB_PORT_CFG && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
end

// ----------------------------------------------------------------------
// RX_PB_PORT_CFG.PORT x8 RW, using RW template.
logic [3:0] up_RX_PB_PORT_CFG_PORT;
always_comb begin
 up_RX_PB_PORT_CFG_PORT =
    ({4{write_req_RX_PB_PORT_CFG }} &
    be[3:0]);
end

logic [31:0] nxt_RX_PB_PORT_CFG_PORT;
always_comb begin
 nxt_RX_PB_PORT_CFG_PORT = write_data[31:0];

end


`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_PORT_CFG_PORT[0], nxt_RX_PB_PORT_CFG_PORT[7:0], RX_PB_PORT_CFG.PORT[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_PORT_CFG_PORT[1], nxt_RX_PB_PORT_CFG_PORT[15:8], RX_PB_PORT_CFG.PORT[15:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_PORT_CFG_PORT[2], nxt_RX_PB_PORT_CFG_PORT[23:16], RX_PB_PORT_CFG.PORT[23:16])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_PORT_CFG_PORT[3], nxt_RX_PB_PORT_CFG_PORT[31:24], RX_PB_PORT_CFG.PORT[31:24])

//---------------------------------------------------------------------
// RX_PB_WM Address Decode
logic [16:0][7:0] addr_decode_RX_PB_WM;
logic [16:0][7:0] write_req_RX_PB_WM;
always_comb begin
   addr_decode_RX_PB_WM[0][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][0]) && req.valid ;
   addr_decode_RX_PB_WM[0][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][1]) && req.valid ;
   addr_decode_RX_PB_WM[0][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][2]) && req.valid ;
   addr_decode_RX_PB_WM[0][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][3]) && req.valid ;
   addr_decode_RX_PB_WM[0][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][4]) && req.valid ;
   addr_decode_RX_PB_WM[0][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][5]) && req.valid ;
   addr_decode_RX_PB_WM[0][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][6]) && req.valid ;
   addr_decode_RX_PB_WM[0][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[0][7]) && req.valid ;
   addr_decode_RX_PB_WM[1][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][0]) && req.valid ;
   addr_decode_RX_PB_WM[1][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][1]) && req.valid ;
   addr_decode_RX_PB_WM[1][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][2]) && req.valid ;
   addr_decode_RX_PB_WM[1][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][3]) && req.valid ;
   addr_decode_RX_PB_WM[1][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][4]) && req.valid ;
   addr_decode_RX_PB_WM[1][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][5]) && req.valid ;
   addr_decode_RX_PB_WM[1][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][6]) && req.valid ;
   addr_decode_RX_PB_WM[1][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[1][7]) && req.valid ;
   addr_decode_RX_PB_WM[2][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][0]) && req.valid ;
   addr_decode_RX_PB_WM[2][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][1]) && req.valid ;
   addr_decode_RX_PB_WM[2][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][2]) && req.valid ;
   addr_decode_RX_PB_WM[2][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][3]) && req.valid ;
   addr_decode_RX_PB_WM[2][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][4]) && req.valid ;
   addr_decode_RX_PB_WM[2][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][5]) && req.valid ;
   addr_decode_RX_PB_WM[2][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][6]) && req.valid ;
   addr_decode_RX_PB_WM[2][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[2][7]) && req.valid ;
   addr_decode_RX_PB_WM[3][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][0]) && req.valid ;
   addr_decode_RX_PB_WM[3][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][1]) && req.valid ;
   addr_decode_RX_PB_WM[3][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][2]) && req.valid ;
   addr_decode_RX_PB_WM[3][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][3]) && req.valid ;
   addr_decode_RX_PB_WM[3][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][4]) && req.valid ;
   addr_decode_RX_PB_WM[3][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][5]) && req.valid ;
   addr_decode_RX_PB_WM[3][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][6]) && req.valid ;
   addr_decode_RX_PB_WM[3][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[3][7]) && req.valid ;
   addr_decode_RX_PB_WM[4][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][0]) && req.valid ;
   addr_decode_RX_PB_WM[4][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][1]) && req.valid ;
   addr_decode_RX_PB_WM[4][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][2]) && req.valid ;
   addr_decode_RX_PB_WM[4][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][3]) && req.valid ;
   addr_decode_RX_PB_WM[4][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][4]) && req.valid ;
   addr_decode_RX_PB_WM[4][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][5]) && req.valid ;
   addr_decode_RX_PB_WM[4][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][6]) && req.valid ;
   addr_decode_RX_PB_WM[4][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[4][7]) && req.valid ;
   addr_decode_RX_PB_WM[5][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][0]) && req.valid ;
   addr_decode_RX_PB_WM[5][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][1]) && req.valid ;
   addr_decode_RX_PB_WM[5][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][2]) && req.valid ;
   addr_decode_RX_PB_WM[5][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][3]) && req.valid ;
   addr_decode_RX_PB_WM[5][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][4]) && req.valid ;
   addr_decode_RX_PB_WM[5][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][5]) && req.valid ;
   addr_decode_RX_PB_WM[5][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][6]) && req.valid ;
   addr_decode_RX_PB_WM[5][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[5][7]) && req.valid ;
   addr_decode_RX_PB_WM[6][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][0]) && req.valid ;
   addr_decode_RX_PB_WM[6][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][1]) && req.valid ;
   addr_decode_RX_PB_WM[6][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][2]) && req.valid ;
   addr_decode_RX_PB_WM[6][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][3]) && req.valid ;
   addr_decode_RX_PB_WM[6][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][4]) && req.valid ;
   addr_decode_RX_PB_WM[6][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][5]) && req.valid ;
   addr_decode_RX_PB_WM[6][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][6]) && req.valid ;
   addr_decode_RX_PB_WM[6][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[6][7]) && req.valid ;
   addr_decode_RX_PB_WM[7][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][0]) && req.valid ;
   addr_decode_RX_PB_WM[7][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][1]) && req.valid ;
   addr_decode_RX_PB_WM[7][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][2]) && req.valid ;
   addr_decode_RX_PB_WM[7][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][3]) && req.valid ;
   addr_decode_RX_PB_WM[7][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][4]) && req.valid ;
   addr_decode_RX_PB_WM[7][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][5]) && req.valid ;
   addr_decode_RX_PB_WM[7][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][6]) && req.valid ;
   addr_decode_RX_PB_WM[7][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[7][7]) && req.valid ;
   addr_decode_RX_PB_WM[8][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][0]) && req.valid ;
   addr_decode_RX_PB_WM[8][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][1]) && req.valid ;
   addr_decode_RX_PB_WM[8][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][2]) && req.valid ;
   addr_decode_RX_PB_WM[8][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][3]) && req.valid ;
   addr_decode_RX_PB_WM[8][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][4]) && req.valid ;
   addr_decode_RX_PB_WM[8][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][5]) && req.valid ;
   addr_decode_RX_PB_WM[8][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][6]) && req.valid ;
   addr_decode_RX_PB_WM[8][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[8][7]) && req.valid ;
   addr_decode_RX_PB_WM[9][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][0]) && req.valid ;
   addr_decode_RX_PB_WM[9][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][1]) && req.valid ;
   addr_decode_RX_PB_WM[9][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][2]) && req.valid ;
   addr_decode_RX_PB_WM[9][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][3]) && req.valid ;
   addr_decode_RX_PB_WM[9][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][4]) && req.valid ;
   addr_decode_RX_PB_WM[9][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][5]) && req.valid ;
   addr_decode_RX_PB_WM[9][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][6]) && req.valid ;
   addr_decode_RX_PB_WM[9][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[9][7]) && req.valid ;
   addr_decode_RX_PB_WM[10][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][0]) && req.valid ;
   addr_decode_RX_PB_WM[10][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][1]) && req.valid ;
   addr_decode_RX_PB_WM[10][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][2]) && req.valid ;
   addr_decode_RX_PB_WM[10][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][3]) && req.valid ;
   addr_decode_RX_PB_WM[10][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][4]) && req.valid ;
   addr_decode_RX_PB_WM[10][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][5]) && req.valid ;
   addr_decode_RX_PB_WM[10][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][6]) && req.valid ;
   addr_decode_RX_PB_WM[10][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[10][7]) && req.valid ;
   addr_decode_RX_PB_WM[11][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][0]) && req.valid ;
   addr_decode_RX_PB_WM[11][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][1]) && req.valid ;
   addr_decode_RX_PB_WM[11][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][2]) && req.valid ;
   addr_decode_RX_PB_WM[11][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][3]) && req.valid ;
   addr_decode_RX_PB_WM[11][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][4]) && req.valid ;
   addr_decode_RX_PB_WM[11][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][5]) && req.valid ;
   addr_decode_RX_PB_WM[11][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][6]) && req.valid ;
   addr_decode_RX_PB_WM[11][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[11][7]) && req.valid ;
   addr_decode_RX_PB_WM[12][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][0]) && req.valid ;
   addr_decode_RX_PB_WM[12][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][1]) && req.valid ;
   addr_decode_RX_PB_WM[12][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][2]) && req.valid ;
   addr_decode_RX_PB_WM[12][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][3]) && req.valid ;
   addr_decode_RX_PB_WM[12][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][4]) && req.valid ;
   addr_decode_RX_PB_WM[12][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][5]) && req.valid ;
   addr_decode_RX_PB_WM[12][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][6]) && req.valid ;
   addr_decode_RX_PB_WM[12][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[12][7]) && req.valid ;
   addr_decode_RX_PB_WM[13][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][0]) && req.valid ;
   addr_decode_RX_PB_WM[13][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][1]) && req.valid ;
   addr_decode_RX_PB_WM[13][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][2]) && req.valid ;
   addr_decode_RX_PB_WM[13][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][3]) && req.valid ;
   addr_decode_RX_PB_WM[13][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][4]) && req.valid ;
   addr_decode_RX_PB_WM[13][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][5]) && req.valid ;
   addr_decode_RX_PB_WM[13][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][6]) && req.valid ;
   addr_decode_RX_PB_WM[13][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[13][7]) && req.valid ;
   addr_decode_RX_PB_WM[14][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][0]) && req.valid ;
   addr_decode_RX_PB_WM[14][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][1]) && req.valid ;
   addr_decode_RX_PB_WM[14][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][2]) && req.valid ;
   addr_decode_RX_PB_WM[14][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][3]) && req.valid ;
   addr_decode_RX_PB_WM[14][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][4]) && req.valid ;
   addr_decode_RX_PB_WM[14][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][5]) && req.valid ;
   addr_decode_RX_PB_WM[14][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][6]) && req.valid ;
   addr_decode_RX_PB_WM[14][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[14][7]) && req.valid ;
   addr_decode_RX_PB_WM[15][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][0]) && req.valid ;
   addr_decode_RX_PB_WM[15][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][1]) && req.valid ;
   addr_decode_RX_PB_WM[15][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][2]) && req.valid ;
   addr_decode_RX_PB_WM[15][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][3]) && req.valid ;
   addr_decode_RX_PB_WM[15][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][4]) && req.valid ;
   addr_decode_RX_PB_WM[15][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][5]) && req.valid ;
   addr_decode_RX_PB_WM[15][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][6]) && req.valid ;
   addr_decode_RX_PB_WM[15][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[15][7]) && req.valid ;
   addr_decode_RX_PB_WM[16][0] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][0]) && req.valid ;
   addr_decode_RX_PB_WM[16][1] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][1]) && req.valid ;
   addr_decode_RX_PB_WM[16][2] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][2]) && req.valid ;
   addr_decode_RX_PB_WM[16][3] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][3]) && req.valid ;
   addr_decode_RX_PB_WM[16][4] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][4]) && req.valid ;
   addr_decode_RX_PB_WM[16][5] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][5]) && req.valid ;
   addr_decode_RX_PB_WM[16][6] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][6]) && req.valid ;
   addr_decode_RX_PB_WM[16][7] = (req_addr[MBY_RX_PB_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == RX_PB_WM_DECODE_ADDR[16][7]) && req.valid ;
   write_req_RX_PB_WM[0][0] = IsMEMWr && addr_decode_RX_PB_WM[0][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[0][1] = IsMEMWr && addr_decode_RX_PB_WM[0][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[0][2] = IsMEMWr && addr_decode_RX_PB_WM[0][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[0][3] = IsMEMWr && addr_decode_RX_PB_WM[0][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[0][4] = IsMEMWr && addr_decode_RX_PB_WM[0][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[0][5] = IsMEMWr && addr_decode_RX_PB_WM[0][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[0][6] = IsMEMWr && addr_decode_RX_PB_WM[0][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[0][7] = IsMEMWr && addr_decode_RX_PB_WM[0][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][0] = IsMEMWr && addr_decode_RX_PB_WM[1][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][1] = IsMEMWr && addr_decode_RX_PB_WM[1][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][2] = IsMEMWr && addr_decode_RX_PB_WM[1][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][3] = IsMEMWr && addr_decode_RX_PB_WM[1][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][4] = IsMEMWr && addr_decode_RX_PB_WM[1][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][5] = IsMEMWr && addr_decode_RX_PB_WM[1][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][6] = IsMEMWr && addr_decode_RX_PB_WM[1][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[1][7] = IsMEMWr && addr_decode_RX_PB_WM[1][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][0] = IsMEMWr && addr_decode_RX_PB_WM[2][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][1] = IsMEMWr && addr_decode_RX_PB_WM[2][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][2] = IsMEMWr && addr_decode_RX_PB_WM[2][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][3] = IsMEMWr && addr_decode_RX_PB_WM[2][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][4] = IsMEMWr && addr_decode_RX_PB_WM[2][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][5] = IsMEMWr && addr_decode_RX_PB_WM[2][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][6] = IsMEMWr && addr_decode_RX_PB_WM[2][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[2][7] = IsMEMWr && addr_decode_RX_PB_WM[2][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][0] = IsMEMWr && addr_decode_RX_PB_WM[3][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][1] = IsMEMWr && addr_decode_RX_PB_WM[3][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][2] = IsMEMWr && addr_decode_RX_PB_WM[3][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][3] = IsMEMWr && addr_decode_RX_PB_WM[3][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][4] = IsMEMWr && addr_decode_RX_PB_WM[3][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][5] = IsMEMWr && addr_decode_RX_PB_WM[3][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][6] = IsMEMWr && addr_decode_RX_PB_WM[3][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[3][7] = IsMEMWr && addr_decode_RX_PB_WM[3][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][0] = IsMEMWr && addr_decode_RX_PB_WM[4][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][1] = IsMEMWr && addr_decode_RX_PB_WM[4][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][2] = IsMEMWr && addr_decode_RX_PB_WM[4][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][3] = IsMEMWr && addr_decode_RX_PB_WM[4][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][4] = IsMEMWr && addr_decode_RX_PB_WM[4][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][5] = IsMEMWr && addr_decode_RX_PB_WM[4][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][6] = IsMEMWr && addr_decode_RX_PB_WM[4][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[4][7] = IsMEMWr && addr_decode_RX_PB_WM[4][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][0] = IsMEMWr && addr_decode_RX_PB_WM[5][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][1] = IsMEMWr && addr_decode_RX_PB_WM[5][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][2] = IsMEMWr && addr_decode_RX_PB_WM[5][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][3] = IsMEMWr && addr_decode_RX_PB_WM[5][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][4] = IsMEMWr && addr_decode_RX_PB_WM[5][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][5] = IsMEMWr && addr_decode_RX_PB_WM[5][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][6] = IsMEMWr && addr_decode_RX_PB_WM[5][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[5][7] = IsMEMWr && addr_decode_RX_PB_WM[5][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][0] = IsMEMWr && addr_decode_RX_PB_WM[6][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][1] = IsMEMWr && addr_decode_RX_PB_WM[6][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][2] = IsMEMWr && addr_decode_RX_PB_WM[6][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][3] = IsMEMWr && addr_decode_RX_PB_WM[6][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][4] = IsMEMWr && addr_decode_RX_PB_WM[6][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][5] = IsMEMWr && addr_decode_RX_PB_WM[6][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][6] = IsMEMWr && addr_decode_RX_PB_WM[6][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[6][7] = IsMEMWr && addr_decode_RX_PB_WM[6][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][0] = IsMEMWr && addr_decode_RX_PB_WM[7][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][1] = IsMEMWr && addr_decode_RX_PB_WM[7][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][2] = IsMEMWr && addr_decode_RX_PB_WM[7][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][3] = IsMEMWr && addr_decode_RX_PB_WM[7][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][4] = IsMEMWr && addr_decode_RX_PB_WM[7][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][5] = IsMEMWr && addr_decode_RX_PB_WM[7][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][6] = IsMEMWr && addr_decode_RX_PB_WM[7][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[7][7] = IsMEMWr && addr_decode_RX_PB_WM[7][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][0] = IsMEMWr && addr_decode_RX_PB_WM[8][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][1] = IsMEMWr && addr_decode_RX_PB_WM[8][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][2] = IsMEMWr && addr_decode_RX_PB_WM[8][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][3] = IsMEMWr && addr_decode_RX_PB_WM[8][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][4] = IsMEMWr && addr_decode_RX_PB_WM[8][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][5] = IsMEMWr && addr_decode_RX_PB_WM[8][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][6] = IsMEMWr && addr_decode_RX_PB_WM[8][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[8][7] = IsMEMWr && addr_decode_RX_PB_WM[8][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][0] = IsMEMWr && addr_decode_RX_PB_WM[9][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][1] = IsMEMWr && addr_decode_RX_PB_WM[9][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][2] = IsMEMWr && addr_decode_RX_PB_WM[9][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][3] = IsMEMWr && addr_decode_RX_PB_WM[9][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][4] = IsMEMWr && addr_decode_RX_PB_WM[9][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][5] = IsMEMWr && addr_decode_RX_PB_WM[9][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][6] = IsMEMWr && addr_decode_RX_PB_WM[9][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[9][7] = IsMEMWr && addr_decode_RX_PB_WM[9][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][0] = IsMEMWr && addr_decode_RX_PB_WM[10][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][1] = IsMEMWr && addr_decode_RX_PB_WM[10][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][2] = IsMEMWr && addr_decode_RX_PB_WM[10][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][3] = IsMEMWr && addr_decode_RX_PB_WM[10][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][4] = IsMEMWr && addr_decode_RX_PB_WM[10][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][5] = IsMEMWr && addr_decode_RX_PB_WM[10][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][6] = IsMEMWr && addr_decode_RX_PB_WM[10][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[10][7] = IsMEMWr && addr_decode_RX_PB_WM[10][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][0] = IsMEMWr && addr_decode_RX_PB_WM[11][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][1] = IsMEMWr && addr_decode_RX_PB_WM[11][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][2] = IsMEMWr && addr_decode_RX_PB_WM[11][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][3] = IsMEMWr && addr_decode_RX_PB_WM[11][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][4] = IsMEMWr && addr_decode_RX_PB_WM[11][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][5] = IsMEMWr && addr_decode_RX_PB_WM[11][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][6] = IsMEMWr && addr_decode_RX_PB_WM[11][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[11][7] = IsMEMWr && addr_decode_RX_PB_WM[11][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][0] = IsMEMWr && addr_decode_RX_PB_WM[12][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][1] = IsMEMWr && addr_decode_RX_PB_WM[12][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][2] = IsMEMWr && addr_decode_RX_PB_WM[12][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][3] = IsMEMWr && addr_decode_RX_PB_WM[12][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][4] = IsMEMWr && addr_decode_RX_PB_WM[12][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][5] = IsMEMWr && addr_decode_RX_PB_WM[12][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][6] = IsMEMWr && addr_decode_RX_PB_WM[12][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[12][7] = IsMEMWr && addr_decode_RX_PB_WM[12][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][0] = IsMEMWr && addr_decode_RX_PB_WM[13][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][1] = IsMEMWr && addr_decode_RX_PB_WM[13][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][2] = IsMEMWr && addr_decode_RX_PB_WM[13][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][3] = IsMEMWr && addr_decode_RX_PB_WM[13][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][4] = IsMEMWr && addr_decode_RX_PB_WM[13][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][5] = IsMEMWr && addr_decode_RX_PB_WM[13][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][6] = IsMEMWr && addr_decode_RX_PB_WM[13][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[13][7] = IsMEMWr && addr_decode_RX_PB_WM[13][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][0] = IsMEMWr && addr_decode_RX_PB_WM[14][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][1] = IsMEMWr && addr_decode_RX_PB_WM[14][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][2] = IsMEMWr && addr_decode_RX_PB_WM[14][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][3] = IsMEMWr && addr_decode_RX_PB_WM[14][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][4] = IsMEMWr && addr_decode_RX_PB_WM[14][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][5] = IsMEMWr && addr_decode_RX_PB_WM[14][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][6] = IsMEMWr && addr_decode_RX_PB_WM[14][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[14][7] = IsMEMWr && addr_decode_RX_PB_WM[14][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][0] = IsMEMWr && addr_decode_RX_PB_WM[15][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][1] = IsMEMWr && addr_decode_RX_PB_WM[15][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][2] = IsMEMWr && addr_decode_RX_PB_WM[15][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][3] = IsMEMWr && addr_decode_RX_PB_WM[15][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][4] = IsMEMWr && addr_decode_RX_PB_WM[15][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][5] = IsMEMWr && addr_decode_RX_PB_WM[15][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][6] = IsMEMWr && addr_decode_RX_PB_WM[15][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[15][7] = IsMEMWr && addr_decode_RX_PB_WM[15][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][0] = IsMEMWr && addr_decode_RX_PB_WM[16][0] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][1] = IsMEMWr && addr_decode_RX_PB_WM[16][1] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][2] = IsMEMWr && addr_decode_RX_PB_WM[16][2] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][3] = IsMEMWr && addr_decode_RX_PB_WM[16][3] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][4] = IsMEMWr && addr_decode_RX_PB_WM[16][4] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][5] = IsMEMWr && addr_decode_RX_PB_WM[16][5] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][6] = IsMEMWr && addr_decode_RX_PB_WM[16][6] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
   write_req_RX_PB_WM[16][7] = IsMEMWr && addr_decode_RX_PB_WM[16][7] && sb_fid_cond_mby_rx_pb_map && sb_bar_cond_mby_rx_pb_map;
end

// ----------------------------------------------------------------------
// RX_PB_WM.XOFF_OR_DROP x2 RW, using RW template.
logic [16:0][7:0][1:0] up_RX_PB_WM_XOFF_OR_DROP;
always_comb begin
 up_RX_PB_WM_XOFF_OR_DROP[0][0] =
    ({2{write_req_RX_PB_WM[0][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[0][1] =
    ({2{write_req_RX_PB_WM[0][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[0][2] =
    ({2{write_req_RX_PB_WM[0][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[0][3] =
    ({2{write_req_RX_PB_WM[0][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[0][4] =
    ({2{write_req_RX_PB_WM[0][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[0][5] =
    ({2{write_req_RX_PB_WM[0][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[0][6] =
    ({2{write_req_RX_PB_WM[0][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[0][7] =
    ({2{write_req_RX_PB_WM[0][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][0] =
    ({2{write_req_RX_PB_WM[1][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][1] =
    ({2{write_req_RX_PB_WM[1][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][2] =
    ({2{write_req_RX_PB_WM[1][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][3] =
    ({2{write_req_RX_PB_WM[1][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][4] =
    ({2{write_req_RX_PB_WM[1][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][5] =
    ({2{write_req_RX_PB_WM[1][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][6] =
    ({2{write_req_RX_PB_WM[1][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[1][7] =
    ({2{write_req_RX_PB_WM[1][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][0] =
    ({2{write_req_RX_PB_WM[2][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][1] =
    ({2{write_req_RX_PB_WM[2][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][2] =
    ({2{write_req_RX_PB_WM[2][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][3] =
    ({2{write_req_RX_PB_WM[2][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][4] =
    ({2{write_req_RX_PB_WM[2][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][5] =
    ({2{write_req_RX_PB_WM[2][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][6] =
    ({2{write_req_RX_PB_WM[2][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[2][7] =
    ({2{write_req_RX_PB_WM[2][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][0] =
    ({2{write_req_RX_PB_WM[3][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][1] =
    ({2{write_req_RX_PB_WM[3][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][2] =
    ({2{write_req_RX_PB_WM[3][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][3] =
    ({2{write_req_RX_PB_WM[3][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][4] =
    ({2{write_req_RX_PB_WM[3][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][5] =
    ({2{write_req_RX_PB_WM[3][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][6] =
    ({2{write_req_RX_PB_WM[3][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[3][7] =
    ({2{write_req_RX_PB_WM[3][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][0] =
    ({2{write_req_RX_PB_WM[4][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][1] =
    ({2{write_req_RX_PB_WM[4][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][2] =
    ({2{write_req_RX_PB_WM[4][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][3] =
    ({2{write_req_RX_PB_WM[4][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][4] =
    ({2{write_req_RX_PB_WM[4][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][5] =
    ({2{write_req_RX_PB_WM[4][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][6] =
    ({2{write_req_RX_PB_WM[4][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[4][7] =
    ({2{write_req_RX_PB_WM[4][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][0] =
    ({2{write_req_RX_PB_WM[5][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][1] =
    ({2{write_req_RX_PB_WM[5][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][2] =
    ({2{write_req_RX_PB_WM[5][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][3] =
    ({2{write_req_RX_PB_WM[5][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][4] =
    ({2{write_req_RX_PB_WM[5][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][5] =
    ({2{write_req_RX_PB_WM[5][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][6] =
    ({2{write_req_RX_PB_WM[5][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[5][7] =
    ({2{write_req_RX_PB_WM[5][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][0] =
    ({2{write_req_RX_PB_WM[6][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][1] =
    ({2{write_req_RX_PB_WM[6][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][2] =
    ({2{write_req_RX_PB_WM[6][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][3] =
    ({2{write_req_RX_PB_WM[6][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][4] =
    ({2{write_req_RX_PB_WM[6][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][5] =
    ({2{write_req_RX_PB_WM[6][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][6] =
    ({2{write_req_RX_PB_WM[6][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[6][7] =
    ({2{write_req_RX_PB_WM[6][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][0] =
    ({2{write_req_RX_PB_WM[7][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][1] =
    ({2{write_req_RX_PB_WM[7][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][2] =
    ({2{write_req_RX_PB_WM[7][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][3] =
    ({2{write_req_RX_PB_WM[7][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][4] =
    ({2{write_req_RX_PB_WM[7][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][5] =
    ({2{write_req_RX_PB_WM[7][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][6] =
    ({2{write_req_RX_PB_WM[7][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[7][7] =
    ({2{write_req_RX_PB_WM[7][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][0] =
    ({2{write_req_RX_PB_WM[8][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][1] =
    ({2{write_req_RX_PB_WM[8][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][2] =
    ({2{write_req_RX_PB_WM[8][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][3] =
    ({2{write_req_RX_PB_WM[8][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][4] =
    ({2{write_req_RX_PB_WM[8][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][5] =
    ({2{write_req_RX_PB_WM[8][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][6] =
    ({2{write_req_RX_PB_WM[8][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[8][7] =
    ({2{write_req_RX_PB_WM[8][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][0] =
    ({2{write_req_RX_PB_WM[9][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][1] =
    ({2{write_req_RX_PB_WM[9][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][2] =
    ({2{write_req_RX_PB_WM[9][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][3] =
    ({2{write_req_RX_PB_WM[9][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][4] =
    ({2{write_req_RX_PB_WM[9][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][5] =
    ({2{write_req_RX_PB_WM[9][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][6] =
    ({2{write_req_RX_PB_WM[9][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[9][7] =
    ({2{write_req_RX_PB_WM[9][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][0] =
    ({2{write_req_RX_PB_WM[10][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][1] =
    ({2{write_req_RX_PB_WM[10][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][2] =
    ({2{write_req_RX_PB_WM[10][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][3] =
    ({2{write_req_RX_PB_WM[10][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][4] =
    ({2{write_req_RX_PB_WM[10][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][5] =
    ({2{write_req_RX_PB_WM[10][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][6] =
    ({2{write_req_RX_PB_WM[10][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[10][7] =
    ({2{write_req_RX_PB_WM[10][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][0] =
    ({2{write_req_RX_PB_WM[11][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][1] =
    ({2{write_req_RX_PB_WM[11][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][2] =
    ({2{write_req_RX_PB_WM[11][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][3] =
    ({2{write_req_RX_PB_WM[11][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][4] =
    ({2{write_req_RX_PB_WM[11][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][5] =
    ({2{write_req_RX_PB_WM[11][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][6] =
    ({2{write_req_RX_PB_WM[11][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[11][7] =
    ({2{write_req_RX_PB_WM[11][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][0] =
    ({2{write_req_RX_PB_WM[12][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][1] =
    ({2{write_req_RX_PB_WM[12][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][2] =
    ({2{write_req_RX_PB_WM[12][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][3] =
    ({2{write_req_RX_PB_WM[12][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][4] =
    ({2{write_req_RX_PB_WM[12][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][5] =
    ({2{write_req_RX_PB_WM[12][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][6] =
    ({2{write_req_RX_PB_WM[12][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[12][7] =
    ({2{write_req_RX_PB_WM[12][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][0] =
    ({2{write_req_RX_PB_WM[13][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][1] =
    ({2{write_req_RX_PB_WM[13][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][2] =
    ({2{write_req_RX_PB_WM[13][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][3] =
    ({2{write_req_RX_PB_WM[13][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][4] =
    ({2{write_req_RX_PB_WM[13][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][5] =
    ({2{write_req_RX_PB_WM[13][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][6] =
    ({2{write_req_RX_PB_WM[13][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[13][7] =
    ({2{write_req_RX_PB_WM[13][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][0] =
    ({2{write_req_RX_PB_WM[14][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][1] =
    ({2{write_req_RX_PB_WM[14][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][2] =
    ({2{write_req_RX_PB_WM[14][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][3] =
    ({2{write_req_RX_PB_WM[14][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][4] =
    ({2{write_req_RX_PB_WM[14][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][5] =
    ({2{write_req_RX_PB_WM[14][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][6] =
    ({2{write_req_RX_PB_WM[14][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[14][7] =
    ({2{write_req_RX_PB_WM[14][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][0] =
    ({2{write_req_RX_PB_WM[15][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][1] =
    ({2{write_req_RX_PB_WM[15][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][2] =
    ({2{write_req_RX_PB_WM[15][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][3] =
    ({2{write_req_RX_PB_WM[15][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][4] =
    ({2{write_req_RX_PB_WM[15][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][5] =
    ({2{write_req_RX_PB_WM[15][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][6] =
    ({2{write_req_RX_PB_WM[15][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[15][7] =
    ({2{write_req_RX_PB_WM[15][7] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][0] =
    ({2{write_req_RX_PB_WM[16][0] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][1] =
    ({2{write_req_RX_PB_WM[16][1] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][2] =
    ({2{write_req_RX_PB_WM[16][2] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][3] =
    ({2{write_req_RX_PB_WM[16][3] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][4] =
    ({2{write_req_RX_PB_WM[16][4] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][5] =
    ({2{write_req_RX_PB_WM[16][5] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][6] =
    ({2{write_req_RX_PB_WM[16][6] }} &
    be[1:0]);
 up_RX_PB_WM_XOFF_OR_DROP[16][7] =
    ({2{write_req_RX_PB_WM[16][7] }} &
    be[1:0]);
end

logic [16:0][7:0][9:0] nxt_RX_PB_WM_XOFF_OR_DROP;
always_comb begin
 nxt_RX_PB_WM_XOFF_OR_DROP[0][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[0][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[0][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[0][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[0][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[0][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[0][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[0][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[1][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[2][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[3][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[4][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[5][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[6][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[7][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[8][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[9][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[10][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[11][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[12][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[13][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[14][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[15][7] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][0] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][1] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][2] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][3] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][4] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][5] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][6] = write_data[9:0];

 nxt_RX_PB_WM_XOFF_OR_DROP[16][7] = write_data[9:0];

end


`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][0][7:0], RX_PB_WM[0][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][0][9:8], RX_PB_WM[0][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][1][7:0], RX_PB_WM[0][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][1][9:8], RX_PB_WM[0][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][2][7:0], RX_PB_WM[0][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][2][9:8], RX_PB_WM[0][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][3][7:0], RX_PB_WM[0][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][3][9:8], RX_PB_WM[0][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][4][7:0], RX_PB_WM[0][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][4][9:8], RX_PB_WM[0][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][5][7:0], RX_PB_WM[0][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][5][9:8], RX_PB_WM[0][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][6][7:0], RX_PB_WM[0][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][6][9:8], RX_PB_WM[0][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[0][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[0][7][7:0], RX_PB_WM[0][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[0][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[0][7][9:8], RX_PB_WM[0][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][0][7:0], RX_PB_WM[1][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][0][9:8], RX_PB_WM[1][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][1][7:0], RX_PB_WM[1][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][1][9:8], RX_PB_WM[1][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][2][7:0], RX_PB_WM[1][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][2][9:8], RX_PB_WM[1][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][3][7:0], RX_PB_WM[1][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][3][9:8], RX_PB_WM[1][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][4][7:0], RX_PB_WM[1][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][4][9:8], RX_PB_WM[1][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][5][7:0], RX_PB_WM[1][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][5][9:8], RX_PB_WM[1][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][6][7:0], RX_PB_WM[1][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][6][9:8], RX_PB_WM[1][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[1][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[1][7][7:0], RX_PB_WM[1][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[1][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[1][7][9:8], RX_PB_WM[1][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][0][7:0], RX_PB_WM[2][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][0][9:8], RX_PB_WM[2][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][1][7:0], RX_PB_WM[2][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][1][9:8], RX_PB_WM[2][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][2][7:0], RX_PB_WM[2][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][2][9:8], RX_PB_WM[2][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][3][7:0], RX_PB_WM[2][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][3][9:8], RX_PB_WM[2][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][4][7:0], RX_PB_WM[2][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][4][9:8], RX_PB_WM[2][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][5][7:0], RX_PB_WM[2][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][5][9:8], RX_PB_WM[2][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][6][7:0], RX_PB_WM[2][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][6][9:8], RX_PB_WM[2][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[2][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[2][7][7:0], RX_PB_WM[2][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[2][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[2][7][9:8], RX_PB_WM[2][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][0][7:0], RX_PB_WM[3][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][0][9:8], RX_PB_WM[3][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][1][7:0], RX_PB_WM[3][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][1][9:8], RX_PB_WM[3][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][2][7:0], RX_PB_WM[3][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][2][9:8], RX_PB_WM[3][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][3][7:0], RX_PB_WM[3][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][3][9:8], RX_PB_WM[3][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][4][7:0], RX_PB_WM[3][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][4][9:8], RX_PB_WM[3][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][5][7:0], RX_PB_WM[3][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][5][9:8], RX_PB_WM[3][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][6][7:0], RX_PB_WM[3][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][6][9:8], RX_PB_WM[3][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[3][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[3][7][7:0], RX_PB_WM[3][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[3][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[3][7][9:8], RX_PB_WM[3][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][0][7:0], RX_PB_WM[4][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][0][9:8], RX_PB_WM[4][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][1][7:0], RX_PB_WM[4][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][1][9:8], RX_PB_WM[4][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][2][7:0], RX_PB_WM[4][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][2][9:8], RX_PB_WM[4][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][3][7:0], RX_PB_WM[4][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][3][9:8], RX_PB_WM[4][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][4][7:0], RX_PB_WM[4][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][4][9:8], RX_PB_WM[4][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][5][7:0], RX_PB_WM[4][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][5][9:8], RX_PB_WM[4][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][6][7:0], RX_PB_WM[4][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][6][9:8], RX_PB_WM[4][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[4][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[4][7][7:0], RX_PB_WM[4][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[4][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[4][7][9:8], RX_PB_WM[4][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][0][7:0], RX_PB_WM[5][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][0][9:8], RX_PB_WM[5][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][1][7:0], RX_PB_WM[5][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][1][9:8], RX_PB_WM[5][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][2][7:0], RX_PB_WM[5][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][2][9:8], RX_PB_WM[5][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][3][7:0], RX_PB_WM[5][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][3][9:8], RX_PB_WM[5][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][4][7:0], RX_PB_WM[5][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][4][9:8], RX_PB_WM[5][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][5][7:0], RX_PB_WM[5][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][5][9:8], RX_PB_WM[5][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][6][7:0], RX_PB_WM[5][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][6][9:8], RX_PB_WM[5][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[5][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[5][7][7:0], RX_PB_WM[5][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[5][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[5][7][9:8], RX_PB_WM[5][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][0][7:0], RX_PB_WM[6][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][0][9:8], RX_PB_WM[6][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][1][7:0], RX_PB_WM[6][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][1][9:8], RX_PB_WM[6][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][2][7:0], RX_PB_WM[6][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][2][9:8], RX_PB_WM[6][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][3][7:0], RX_PB_WM[6][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][3][9:8], RX_PB_WM[6][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][4][7:0], RX_PB_WM[6][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][4][9:8], RX_PB_WM[6][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][5][7:0], RX_PB_WM[6][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][5][9:8], RX_PB_WM[6][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][6][7:0], RX_PB_WM[6][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][6][9:8], RX_PB_WM[6][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[6][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[6][7][7:0], RX_PB_WM[6][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[6][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[6][7][9:8], RX_PB_WM[6][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][0][7:0], RX_PB_WM[7][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][0][9:8], RX_PB_WM[7][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][1][7:0], RX_PB_WM[7][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][1][9:8], RX_PB_WM[7][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][2][7:0], RX_PB_WM[7][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][2][9:8], RX_PB_WM[7][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][3][7:0], RX_PB_WM[7][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][3][9:8], RX_PB_WM[7][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][4][7:0], RX_PB_WM[7][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][4][9:8], RX_PB_WM[7][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][5][7:0], RX_PB_WM[7][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][5][9:8], RX_PB_WM[7][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][6][7:0], RX_PB_WM[7][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][6][9:8], RX_PB_WM[7][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[7][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[7][7][7:0], RX_PB_WM[7][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[7][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[7][7][9:8], RX_PB_WM[7][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][0][7:0], RX_PB_WM[8][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][0][9:8], RX_PB_WM[8][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][1][7:0], RX_PB_WM[8][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][1][9:8], RX_PB_WM[8][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][2][7:0], RX_PB_WM[8][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][2][9:8], RX_PB_WM[8][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][3][7:0], RX_PB_WM[8][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][3][9:8], RX_PB_WM[8][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][4][7:0], RX_PB_WM[8][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][4][9:8], RX_PB_WM[8][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][5][7:0], RX_PB_WM[8][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][5][9:8], RX_PB_WM[8][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][6][7:0], RX_PB_WM[8][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][6][9:8], RX_PB_WM[8][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[8][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[8][7][7:0], RX_PB_WM[8][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[8][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[8][7][9:8], RX_PB_WM[8][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][0][7:0], RX_PB_WM[9][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][0][9:8], RX_PB_WM[9][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][1][7:0], RX_PB_WM[9][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][1][9:8], RX_PB_WM[9][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][2][7:0], RX_PB_WM[9][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][2][9:8], RX_PB_WM[9][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][3][7:0], RX_PB_WM[9][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][3][9:8], RX_PB_WM[9][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][4][7:0], RX_PB_WM[9][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][4][9:8], RX_PB_WM[9][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][5][7:0], RX_PB_WM[9][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][5][9:8], RX_PB_WM[9][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][6][7:0], RX_PB_WM[9][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][6][9:8], RX_PB_WM[9][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[9][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[9][7][7:0], RX_PB_WM[9][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[9][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[9][7][9:8], RX_PB_WM[9][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][0][7:0], RX_PB_WM[10][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][0][9:8], RX_PB_WM[10][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][1][7:0], RX_PB_WM[10][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][1][9:8], RX_PB_WM[10][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][2][7:0], RX_PB_WM[10][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][2][9:8], RX_PB_WM[10][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][3][7:0], RX_PB_WM[10][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][3][9:8], RX_PB_WM[10][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][4][7:0], RX_PB_WM[10][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][4][9:8], RX_PB_WM[10][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][5][7:0], RX_PB_WM[10][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][5][9:8], RX_PB_WM[10][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][6][7:0], RX_PB_WM[10][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][6][9:8], RX_PB_WM[10][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[10][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[10][7][7:0], RX_PB_WM[10][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[10][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[10][7][9:8], RX_PB_WM[10][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][0][7:0], RX_PB_WM[11][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][0][9:8], RX_PB_WM[11][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][1][7:0], RX_PB_WM[11][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][1][9:8], RX_PB_WM[11][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][2][7:0], RX_PB_WM[11][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][2][9:8], RX_PB_WM[11][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][3][7:0], RX_PB_WM[11][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][3][9:8], RX_PB_WM[11][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][4][7:0], RX_PB_WM[11][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][4][9:8], RX_PB_WM[11][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][5][7:0], RX_PB_WM[11][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][5][9:8], RX_PB_WM[11][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][6][7:0], RX_PB_WM[11][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][6][9:8], RX_PB_WM[11][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[11][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[11][7][7:0], RX_PB_WM[11][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[11][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[11][7][9:8], RX_PB_WM[11][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][0][7:0], RX_PB_WM[12][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][0][9:8], RX_PB_WM[12][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][1][7:0], RX_PB_WM[12][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][1][9:8], RX_PB_WM[12][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][2][7:0], RX_PB_WM[12][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][2][9:8], RX_PB_WM[12][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][3][7:0], RX_PB_WM[12][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][3][9:8], RX_PB_WM[12][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][4][7:0], RX_PB_WM[12][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][4][9:8], RX_PB_WM[12][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][5][7:0], RX_PB_WM[12][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][5][9:8], RX_PB_WM[12][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][6][7:0], RX_PB_WM[12][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][6][9:8], RX_PB_WM[12][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[12][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[12][7][7:0], RX_PB_WM[12][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[12][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[12][7][9:8], RX_PB_WM[12][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][0][7:0], RX_PB_WM[13][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][0][9:8], RX_PB_WM[13][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][1][7:0], RX_PB_WM[13][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][1][9:8], RX_PB_WM[13][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][2][7:0], RX_PB_WM[13][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][2][9:8], RX_PB_WM[13][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][3][7:0], RX_PB_WM[13][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][3][9:8], RX_PB_WM[13][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][4][7:0], RX_PB_WM[13][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][4][9:8], RX_PB_WM[13][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][5][7:0], RX_PB_WM[13][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][5][9:8], RX_PB_WM[13][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][6][7:0], RX_PB_WM[13][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][6][9:8], RX_PB_WM[13][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[13][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[13][7][7:0], RX_PB_WM[13][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[13][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[13][7][9:8], RX_PB_WM[13][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][0][7:0], RX_PB_WM[14][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][0][9:8], RX_PB_WM[14][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][1][7:0], RX_PB_WM[14][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][1][9:8], RX_PB_WM[14][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][2][7:0], RX_PB_WM[14][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][2][9:8], RX_PB_WM[14][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][3][7:0], RX_PB_WM[14][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][3][9:8], RX_PB_WM[14][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][4][7:0], RX_PB_WM[14][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][4][9:8], RX_PB_WM[14][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][5][7:0], RX_PB_WM[14][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][5][9:8], RX_PB_WM[14][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][6][7:0], RX_PB_WM[14][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][6][9:8], RX_PB_WM[14][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[14][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[14][7][7:0], RX_PB_WM[14][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[14][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[14][7][9:8], RX_PB_WM[14][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][0][7:0], RX_PB_WM[15][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][0][9:8], RX_PB_WM[15][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][1][7:0], RX_PB_WM[15][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][1][9:8], RX_PB_WM[15][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][2][7:0], RX_PB_WM[15][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][2][9:8], RX_PB_WM[15][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][3][7:0], RX_PB_WM[15][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][3][9:8], RX_PB_WM[15][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][4][7:0], RX_PB_WM[15][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][4][9:8], RX_PB_WM[15][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][5][7:0], RX_PB_WM[15][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][5][9:8], RX_PB_WM[15][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][6][7:0], RX_PB_WM[15][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][6][9:8], RX_PB_WM[15][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[15][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[15][7][7:0], RX_PB_WM[15][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[15][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[15][7][9:8], RX_PB_WM[15][7].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][0][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][0][7:0], RX_PB_WM[16][0].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][0][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][0][9:8], RX_PB_WM[16][0].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][1][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][1][7:0], RX_PB_WM[16][1].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][1][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][1][9:8], RX_PB_WM[16][1].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][2][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][2][7:0], RX_PB_WM[16][2].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][2][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][2][9:8], RX_PB_WM[16][2].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][3][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][3][7:0], RX_PB_WM[16][3].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][3][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][3][9:8], RX_PB_WM[16][3].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][4][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][4][7:0], RX_PB_WM[16][4].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][4][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][4][9:8], RX_PB_WM[16][4].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][5][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][5][7:0], RX_PB_WM[16][5].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][5][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][5][9:8], RX_PB_WM[16][5].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][6][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][6][7:0], RX_PB_WM[16][6].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][6][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][6][9:8], RX_PB_WM[16][6].XOFF_OR_DROP[9:8])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 8'h0, up_RX_PB_WM_XOFF_OR_DROP[16][7][0], nxt_RX_PB_WM_XOFF_OR_DROP[16][7][7:0], RX_PB_WM[16][7].XOFF_OR_DROP[7:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 2'h2, up_RX_PB_WM_XOFF_OR_DROP[16][7][1], nxt_RX_PB_WM_XOFF_OR_DROP[16][7][9:8], RX_PB_WM[16][7].XOFF_OR_DROP[9:8])

// ----------------------------------------------------------------------
// RX_PB_WM.XON x4 RW, using RW template.
logic [16:0][7:0][1:0] up_RX_PB_WM_XON;
always_comb begin
 up_RX_PB_WM_XON[0][0] =
    ({2{write_req_RX_PB_WM[0][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[0][1] =
    ({2{write_req_RX_PB_WM[0][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[0][2] =
    ({2{write_req_RX_PB_WM[0][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[0][3] =
    ({2{write_req_RX_PB_WM[0][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[0][4] =
    ({2{write_req_RX_PB_WM[0][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[0][5] =
    ({2{write_req_RX_PB_WM[0][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[0][6] =
    ({2{write_req_RX_PB_WM[0][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[0][7] =
    ({2{write_req_RX_PB_WM[0][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][0] =
    ({2{write_req_RX_PB_WM[1][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][1] =
    ({2{write_req_RX_PB_WM[1][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][2] =
    ({2{write_req_RX_PB_WM[1][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][3] =
    ({2{write_req_RX_PB_WM[1][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][4] =
    ({2{write_req_RX_PB_WM[1][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][5] =
    ({2{write_req_RX_PB_WM[1][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][6] =
    ({2{write_req_RX_PB_WM[1][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[1][7] =
    ({2{write_req_RX_PB_WM[1][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][0] =
    ({2{write_req_RX_PB_WM[2][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][1] =
    ({2{write_req_RX_PB_WM[2][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][2] =
    ({2{write_req_RX_PB_WM[2][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][3] =
    ({2{write_req_RX_PB_WM[2][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][4] =
    ({2{write_req_RX_PB_WM[2][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][5] =
    ({2{write_req_RX_PB_WM[2][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][6] =
    ({2{write_req_RX_PB_WM[2][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[2][7] =
    ({2{write_req_RX_PB_WM[2][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][0] =
    ({2{write_req_RX_PB_WM[3][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][1] =
    ({2{write_req_RX_PB_WM[3][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][2] =
    ({2{write_req_RX_PB_WM[3][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][3] =
    ({2{write_req_RX_PB_WM[3][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][4] =
    ({2{write_req_RX_PB_WM[3][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][5] =
    ({2{write_req_RX_PB_WM[3][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][6] =
    ({2{write_req_RX_PB_WM[3][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[3][7] =
    ({2{write_req_RX_PB_WM[3][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][0] =
    ({2{write_req_RX_PB_WM[4][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][1] =
    ({2{write_req_RX_PB_WM[4][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][2] =
    ({2{write_req_RX_PB_WM[4][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][3] =
    ({2{write_req_RX_PB_WM[4][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][4] =
    ({2{write_req_RX_PB_WM[4][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][5] =
    ({2{write_req_RX_PB_WM[4][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][6] =
    ({2{write_req_RX_PB_WM[4][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[4][7] =
    ({2{write_req_RX_PB_WM[4][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][0] =
    ({2{write_req_RX_PB_WM[5][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][1] =
    ({2{write_req_RX_PB_WM[5][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][2] =
    ({2{write_req_RX_PB_WM[5][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][3] =
    ({2{write_req_RX_PB_WM[5][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][4] =
    ({2{write_req_RX_PB_WM[5][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][5] =
    ({2{write_req_RX_PB_WM[5][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][6] =
    ({2{write_req_RX_PB_WM[5][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[5][7] =
    ({2{write_req_RX_PB_WM[5][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][0] =
    ({2{write_req_RX_PB_WM[6][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][1] =
    ({2{write_req_RX_PB_WM[6][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][2] =
    ({2{write_req_RX_PB_WM[6][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][3] =
    ({2{write_req_RX_PB_WM[6][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][4] =
    ({2{write_req_RX_PB_WM[6][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][5] =
    ({2{write_req_RX_PB_WM[6][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][6] =
    ({2{write_req_RX_PB_WM[6][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[6][7] =
    ({2{write_req_RX_PB_WM[6][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][0] =
    ({2{write_req_RX_PB_WM[7][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][1] =
    ({2{write_req_RX_PB_WM[7][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][2] =
    ({2{write_req_RX_PB_WM[7][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][3] =
    ({2{write_req_RX_PB_WM[7][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][4] =
    ({2{write_req_RX_PB_WM[7][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][5] =
    ({2{write_req_RX_PB_WM[7][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][6] =
    ({2{write_req_RX_PB_WM[7][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[7][7] =
    ({2{write_req_RX_PB_WM[7][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][0] =
    ({2{write_req_RX_PB_WM[8][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][1] =
    ({2{write_req_RX_PB_WM[8][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][2] =
    ({2{write_req_RX_PB_WM[8][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][3] =
    ({2{write_req_RX_PB_WM[8][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][4] =
    ({2{write_req_RX_PB_WM[8][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][5] =
    ({2{write_req_RX_PB_WM[8][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][6] =
    ({2{write_req_RX_PB_WM[8][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[8][7] =
    ({2{write_req_RX_PB_WM[8][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][0] =
    ({2{write_req_RX_PB_WM[9][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][1] =
    ({2{write_req_RX_PB_WM[9][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][2] =
    ({2{write_req_RX_PB_WM[9][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][3] =
    ({2{write_req_RX_PB_WM[9][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][4] =
    ({2{write_req_RX_PB_WM[9][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][5] =
    ({2{write_req_RX_PB_WM[9][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][6] =
    ({2{write_req_RX_PB_WM[9][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[9][7] =
    ({2{write_req_RX_PB_WM[9][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][0] =
    ({2{write_req_RX_PB_WM[10][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][1] =
    ({2{write_req_RX_PB_WM[10][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][2] =
    ({2{write_req_RX_PB_WM[10][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][3] =
    ({2{write_req_RX_PB_WM[10][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][4] =
    ({2{write_req_RX_PB_WM[10][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][5] =
    ({2{write_req_RX_PB_WM[10][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][6] =
    ({2{write_req_RX_PB_WM[10][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[10][7] =
    ({2{write_req_RX_PB_WM[10][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][0] =
    ({2{write_req_RX_PB_WM[11][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][1] =
    ({2{write_req_RX_PB_WM[11][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][2] =
    ({2{write_req_RX_PB_WM[11][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][3] =
    ({2{write_req_RX_PB_WM[11][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][4] =
    ({2{write_req_RX_PB_WM[11][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][5] =
    ({2{write_req_RX_PB_WM[11][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][6] =
    ({2{write_req_RX_PB_WM[11][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[11][7] =
    ({2{write_req_RX_PB_WM[11][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][0] =
    ({2{write_req_RX_PB_WM[12][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][1] =
    ({2{write_req_RX_PB_WM[12][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][2] =
    ({2{write_req_RX_PB_WM[12][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][3] =
    ({2{write_req_RX_PB_WM[12][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][4] =
    ({2{write_req_RX_PB_WM[12][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][5] =
    ({2{write_req_RX_PB_WM[12][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][6] =
    ({2{write_req_RX_PB_WM[12][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[12][7] =
    ({2{write_req_RX_PB_WM[12][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][0] =
    ({2{write_req_RX_PB_WM[13][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][1] =
    ({2{write_req_RX_PB_WM[13][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][2] =
    ({2{write_req_RX_PB_WM[13][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][3] =
    ({2{write_req_RX_PB_WM[13][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][4] =
    ({2{write_req_RX_PB_WM[13][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][5] =
    ({2{write_req_RX_PB_WM[13][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][6] =
    ({2{write_req_RX_PB_WM[13][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[13][7] =
    ({2{write_req_RX_PB_WM[13][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][0] =
    ({2{write_req_RX_PB_WM[14][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][1] =
    ({2{write_req_RX_PB_WM[14][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][2] =
    ({2{write_req_RX_PB_WM[14][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][3] =
    ({2{write_req_RX_PB_WM[14][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][4] =
    ({2{write_req_RX_PB_WM[14][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][5] =
    ({2{write_req_RX_PB_WM[14][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][6] =
    ({2{write_req_RX_PB_WM[14][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[14][7] =
    ({2{write_req_RX_PB_WM[14][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][0] =
    ({2{write_req_RX_PB_WM[15][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][1] =
    ({2{write_req_RX_PB_WM[15][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][2] =
    ({2{write_req_RX_PB_WM[15][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][3] =
    ({2{write_req_RX_PB_WM[15][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][4] =
    ({2{write_req_RX_PB_WM[15][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][5] =
    ({2{write_req_RX_PB_WM[15][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][6] =
    ({2{write_req_RX_PB_WM[15][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[15][7] =
    ({2{write_req_RX_PB_WM[15][7] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][0] =
    ({2{write_req_RX_PB_WM[16][0] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][1] =
    ({2{write_req_RX_PB_WM[16][1] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][2] =
    ({2{write_req_RX_PB_WM[16][2] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][3] =
    ({2{write_req_RX_PB_WM[16][3] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][4] =
    ({2{write_req_RX_PB_WM[16][4] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][5] =
    ({2{write_req_RX_PB_WM[16][5] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][6] =
    ({2{write_req_RX_PB_WM[16][6] }} &
    be[2:1]);
 up_RX_PB_WM_XON[16][7] =
    ({2{write_req_RX_PB_WM[16][7] }} &
    be[2:1]);
end

logic [16:0][7:0][9:0] nxt_RX_PB_WM_XON;
always_comb begin
 nxt_RX_PB_WM_XON[0][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[0][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[0][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[0][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[0][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[0][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[0][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[0][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[1][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[2][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[3][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[4][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[5][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[6][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[7][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[8][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[9][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[10][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[11][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[12][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[13][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[14][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[15][7] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][0] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][1] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][2] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][3] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][4] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][5] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][6] = write_data[19:10];

 nxt_RX_PB_WM_XON[16][7] = write_data[19:10];

end


`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][0][0], nxt_RX_PB_WM_XON[0][0][5:0], RX_PB_WM[0][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][0][1], nxt_RX_PB_WM_XON[0][0][9:6], RX_PB_WM[0][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][1][0], nxt_RX_PB_WM_XON[0][1][5:0], RX_PB_WM[0][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][1][1], nxt_RX_PB_WM_XON[0][1][9:6], RX_PB_WM[0][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][2][0], nxt_RX_PB_WM_XON[0][2][5:0], RX_PB_WM[0][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][2][1], nxt_RX_PB_WM_XON[0][2][9:6], RX_PB_WM[0][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][3][0], nxt_RX_PB_WM_XON[0][3][5:0], RX_PB_WM[0][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][3][1], nxt_RX_PB_WM_XON[0][3][9:6], RX_PB_WM[0][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][4][0], nxt_RX_PB_WM_XON[0][4][5:0], RX_PB_WM[0][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][4][1], nxt_RX_PB_WM_XON[0][4][9:6], RX_PB_WM[0][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][5][0], nxt_RX_PB_WM_XON[0][5][5:0], RX_PB_WM[0][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][5][1], nxt_RX_PB_WM_XON[0][5][9:6], RX_PB_WM[0][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][6][0], nxt_RX_PB_WM_XON[0][6][5:0], RX_PB_WM[0][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][6][1], nxt_RX_PB_WM_XON[0][6][9:6], RX_PB_WM[0][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[0][7][0], nxt_RX_PB_WM_XON[0][7][5:0], RX_PB_WM[0][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[0][7][1], nxt_RX_PB_WM_XON[0][7][9:6], RX_PB_WM[0][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][0][0], nxt_RX_PB_WM_XON[1][0][5:0], RX_PB_WM[1][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][0][1], nxt_RX_PB_WM_XON[1][0][9:6], RX_PB_WM[1][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][1][0], nxt_RX_PB_WM_XON[1][1][5:0], RX_PB_WM[1][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][1][1], nxt_RX_PB_WM_XON[1][1][9:6], RX_PB_WM[1][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][2][0], nxt_RX_PB_WM_XON[1][2][5:0], RX_PB_WM[1][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][2][1], nxt_RX_PB_WM_XON[1][2][9:6], RX_PB_WM[1][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][3][0], nxt_RX_PB_WM_XON[1][3][5:0], RX_PB_WM[1][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][3][1], nxt_RX_PB_WM_XON[1][3][9:6], RX_PB_WM[1][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][4][0], nxt_RX_PB_WM_XON[1][4][5:0], RX_PB_WM[1][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][4][1], nxt_RX_PB_WM_XON[1][4][9:6], RX_PB_WM[1][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][5][0], nxt_RX_PB_WM_XON[1][5][5:0], RX_PB_WM[1][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][5][1], nxt_RX_PB_WM_XON[1][5][9:6], RX_PB_WM[1][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][6][0], nxt_RX_PB_WM_XON[1][6][5:0], RX_PB_WM[1][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][6][1], nxt_RX_PB_WM_XON[1][6][9:6], RX_PB_WM[1][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[1][7][0], nxt_RX_PB_WM_XON[1][7][5:0], RX_PB_WM[1][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[1][7][1], nxt_RX_PB_WM_XON[1][7][9:6], RX_PB_WM[1][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][0][0], nxt_RX_PB_WM_XON[2][0][5:0], RX_PB_WM[2][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][0][1], nxt_RX_PB_WM_XON[2][0][9:6], RX_PB_WM[2][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][1][0], nxt_RX_PB_WM_XON[2][1][5:0], RX_PB_WM[2][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][1][1], nxt_RX_PB_WM_XON[2][1][9:6], RX_PB_WM[2][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][2][0], nxt_RX_PB_WM_XON[2][2][5:0], RX_PB_WM[2][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][2][1], nxt_RX_PB_WM_XON[2][2][9:6], RX_PB_WM[2][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][3][0], nxt_RX_PB_WM_XON[2][3][5:0], RX_PB_WM[2][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][3][1], nxt_RX_PB_WM_XON[2][3][9:6], RX_PB_WM[2][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][4][0], nxt_RX_PB_WM_XON[2][4][5:0], RX_PB_WM[2][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][4][1], nxt_RX_PB_WM_XON[2][4][9:6], RX_PB_WM[2][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][5][0], nxt_RX_PB_WM_XON[2][5][5:0], RX_PB_WM[2][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][5][1], nxt_RX_PB_WM_XON[2][5][9:6], RX_PB_WM[2][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][6][0], nxt_RX_PB_WM_XON[2][6][5:0], RX_PB_WM[2][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][6][1], nxt_RX_PB_WM_XON[2][6][9:6], RX_PB_WM[2][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[2][7][0], nxt_RX_PB_WM_XON[2][7][5:0], RX_PB_WM[2][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[2][7][1], nxt_RX_PB_WM_XON[2][7][9:6], RX_PB_WM[2][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][0][0], nxt_RX_PB_WM_XON[3][0][5:0], RX_PB_WM[3][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][0][1], nxt_RX_PB_WM_XON[3][0][9:6], RX_PB_WM[3][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][1][0], nxt_RX_PB_WM_XON[3][1][5:0], RX_PB_WM[3][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][1][1], nxt_RX_PB_WM_XON[3][1][9:6], RX_PB_WM[3][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][2][0], nxt_RX_PB_WM_XON[3][2][5:0], RX_PB_WM[3][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][2][1], nxt_RX_PB_WM_XON[3][2][9:6], RX_PB_WM[3][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][3][0], nxt_RX_PB_WM_XON[3][3][5:0], RX_PB_WM[3][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][3][1], nxt_RX_PB_WM_XON[3][3][9:6], RX_PB_WM[3][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][4][0], nxt_RX_PB_WM_XON[3][4][5:0], RX_PB_WM[3][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][4][1], nxt_RX_PB_WM_XON[3][4][9:6], RX_PB_WM[3][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][5][0], nxt_RX_PB_WM_XON[3][5][5:0], RX_PB_WM[3][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][5][1], nxt_RX_PB_WM_XON[3][5][9:6], RX_PB_WM[3][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][6][0], nxt_RX_PB_WM_XON[3][6][5:0], RX_PB_WM[3][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][6][1], nxt_RX_PB_WM_XON[3][6][9:6], RX_PB_WM[3][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[3][7][0], nxt_RX_PB_WM_XON[3][7][5:0], RX_PB_WM[3][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[3][7][1], nxt_RX_PB_WM_XON[3][7][9:6], RX_PB_WM[3][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][0][0], nxt_RX_PB_WM_XON[4][0][5:0], RX_PB_WM[4][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][0][1], nxt_RX_PB_WM_XON[4][0][9:6], RX_PB_WM[4][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][1][0], nxt_RX_PB_WM_XON[4][1][5:0], RX_PB_WM[4][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][1][1], nxt_RX_PB_WM_XON[4][1][9:6], RX_PB_WM[4][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][2][0], nxt_RX_PB_WM_XON[4][2][5:0], RX_PB_WM[4][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][2][1], nxt_RX_PB_WM_XON[4][2][9:6], RX_PB_WM[4][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][3][0], nxt_RX_PB_WM_XON[4][3][5:0], RX_PB_WM[4][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][3][1], nxt_RX_PB_WM_XON[4][3][9:6], RX_PB_WM[4][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][4][0], nxt_RX_PB_WM_XON[4][4][5:0], RX_PB_WM[4][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][4][1], nxt_RX_PB_WM_XON[4][4][9:6], RX_PB_WM[4][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][5][0], nxt_RX_PB_WM_XON[4][5][5:0], RX_PB_WM[4][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][5][1], nxt_RX_PB_WM_XON[4][5][9:6], RX_PB_WM[4][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][6][0], nxt_RX_PB_WM_XON[4][6][5:0], RX_PB_WM[4][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][6][1], nxt_RX_PB_WM_XON[4][6][9:6], RX_PB_WM[4][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[4][7][0], nxt_RX_PB_WM_XON[4][7][5:0], RX_PB_WM[4][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[4][7][1], nxt_RX_PB_WM_XON[4][7][9:6], RX_PB_WM[4][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][0][0], nxt_RX_PB_WM_XON[5][0][5:0], RX_PB_WM[5][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][0][1], nxt_RX_PB_WM_XON[5][0][9:6], RX_PB_WM[5][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][1][0], nxt_RX_PB_WM_XON[5][1][5:0], RX_PB_WM[5][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][1][1], nxt_RX_PB_WM_XON[5][1][9:6], RX_PB_WM[5][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][2][0], nxt_RX_PB_WM_XON[5][2][5:0], RX_PB_WM[5][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][2][1], nxt_RX_PB_WM_XON[5][2][9:6], RX_PB_WM[5][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][3][0], nxt_RX_PB_WM_XON[5][3][5:0], RX_PB_WM[5][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][3][1], nxt_RX_PB_WM_XON[5][3][9:6], RX_PB_WM[5][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][4][0], nxt_RX_PB_WM_XON[5][4][5:0], RX_PB_WM[5][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][4][1], nxt_RX_PB_WM_XON[5][4][9:6], RX_PB_WM[5][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][5][0], nxt_RX_PB_WM_XON[5][5][5:0], RX_PB_WM[5][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][5][1], nxt_RX_PB_WM_XON[5][5][9:6], RX_PB_WM[5][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][6][0], nxt_RX_PB_WM_XON[5][6][5:0], RX_PB_WM[5][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][6][1], nxt_RX_PB_WM_XON[5][6][9:6], RX_PB_WM[5][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[5][7][0], nxt_RX_PB_WM_XON[5][7][5:0], RX_PB_WM[5][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[5][7][1], nxt_RX_PB_WM_XON[5][7][9:6], RX_PB_WM[5][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][0][0], nxt_RX_PB_WM_XON[6][0][5:0], RX_PB_WM[6][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][0][1], nxt_RX_PB_WM_XON[6][0][9:6], RX_PB_WM[6][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][1][0], nxt_RX_PB_WM_XON[6][1][5:0], RX_PB_WM[6][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][1][1], nxt_RX_PB_WM_XON[6][1][9:6], RX_PB_WM[6][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][2][0], nxt_RX_PB_WM_XON[6][2][5:0], RX_PB_WM[6][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][2][1], nxt_RX_PB_WM_XON[6][2][9:6], RX_PB_WM[6][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][3][0], nxt_RX_PB_WM_XON[6][3][5:0], RX_PB_WM[6][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][3][1], nxt_RX_PB_WM_XON[6][3][9:6], RX_PB_WM[6][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][4][0], nxt_RX_PB_WM_XON[6][4][5:0], RX_PB_WM[6][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][4][1], nxt_RX_PB_WM_XON[6][4][9:6], RX_PB_WM[6][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][5][0], nxt_RX_PB_WM_XON[6][5][5:0], RX_PB_WM[6][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][5][1], nxt_RX_PB_WM_XON[6][5][9:6], RX_PB_WM[6][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][6][0], nxt_RX_PB_WM_XON[6][6][5:0], RX_PB_WM[6][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][6][1], nxt_RX_PB_WM_XON[6][6][9:6], RX_PB_WM[6][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[6][7][0], nxt_RX_PB_WM_XON[6][7][5:0], RX_PB_WM[6][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[6][7][1], nxt_RX_PB_WM_XON[6][7][9:6], RX_PB_WM[6][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][0][0], nxt_RX_PB_WM_XON[7][0][5:0], RX_PB_WM[7][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][0][1], nxt_RX_PB_WM_XON[7][0][9:6], RX_PB_WM[7][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][1][0], nxt_RX_PB_WM_XON[7][1][5:0], RX_PB_WM[7][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][1][1], nxt_RX_PB_WM_XON[7][1][9:6], RX_PB_WM[7][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][2][0], nxt_RX_PB_WM_XON[7][2][5:0], RX_PB_WM[7][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][2][1], nxt_RX_PB_WM_XON[7][2][9:6], RX_PB_WM[7][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][3][0], nxt_RX_PB_WM_XON[7][3][5:0], RX_PB_WM[7][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][3][1], nxt_RX_PB_WM_XON[7][3][9:6], RX_PB_WM[7][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][4][0], nxt_RX_PB_WM_XON[7][4][5:0], RX_PB_WM[7][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][4][1], nxt_RX_PB_WM_XON[7][4][9:6], RX_PB_WM[7][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][5][0], nxt_RX_PB_WM_XON[7][5][5:0], RX_PB_WM[7][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][5][1], nxt_RX_PB_WM_XON[7][5][9:6], RX_PB_WM[7][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][6][0], nxt_RX_PB_WM_XON[7][6][5:0], RX_PB_WM[7][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][6][1], nxt_RX_PB_WM_XON[7][6][9:6], RX_PB_WM[7][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[7][7][0], nxt_RX_PB_WM_XON[7][7][5:0], RX_PB_WM[7][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[7][7][1], nxt_RX_PB_WM_XON[7][7][9:6], RX_PB_WM[7][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][0][0], nxt_RX_PB_WM_XON[8][0][5:0], RX_PB_WM[8][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][0][1], nxt_RX_PB_WM_XON[8][0][9:6], RX_PB_WM[8][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][1][0], nxt_RX_PB_WM_XON[8][1][5:0], RX_PB_WM[8][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][1][1], nxt_RX_PB_WM_XON[8][1][9:6], RX_PB_WM[8][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][2][0], nxt_RX_PB_WM_XON[8][2][5:0], RX_PB_WM[8][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][2][1], nxt_RX_PB_WM_XON[8][2][9:6], RX_PB_WM[8][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][3][0], nxt_RX_PB_WM_XON[8][3][5:0], RX_PB_WM[8][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][3][1], nxt_RX_PB_WM_XON[8][3][9:6], RX_PB_WM[8][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][4][0], nxt_RX_PB_WM_XON[8][4][5:0], RX_PB_WM[8][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][4][1], nxt_RX_PB_WM_XON[8][4][9:6], RX_PB_WM[8][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][5][0], nxt_RX_PB_WM_XON[8][5][5:0], RX_PB_WM[8][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][5][1], nxt_RX_PB_WM_XON[8][5][9:6], RX_PB_WM[8][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][6][0], nxt_RX_PB_WM_XON[8][6][5:0], RX_PB_WM[8][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][6][1], nxt_RX_PB_WM_XON[8][6][9:6], RX_PB_WM[8][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[8][7][0], nxt_RX_PB_WM_XON[8][7][5:0], RX_PB_WM[8][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[8][7][1], nxt_RX_PB_WM_XON[8][7][9:6], RX_PB_WM[8][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][0][0], nxt_RX_PB_WM_XON[9][0][5:0], RX_PB_WM[9][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][0][1], nxt_RX_PB_WM_XON[9][0][9:6], RX_PB_WM[9][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][1][0], nxt_RX_PB_WM_XON[9][1][5:0], RX_PB_WM[9][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][1][1], nxt_RX_PB_WM_XON[9][1][9:6], RX_PB_WM[9][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][2][0], nxt_RX_PB_WM_XON[9][2][5:0], RX_PB_WM[9][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][2][1], nxt_RX_PB_WM_XON[9][2][9:6], RX_PB_WM[9][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][3][0], nxt_RX_PB_WM_XON[9][3][5:0], RX_PB_WM[9][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][3][1], nxt_RX_PB_WM_XON[9][3][9:6], RX_PB_WM[9][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][4][0], nxt_RX_PB_WM_XON[9][4][5:0], RX_PB_WM[9][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][4][1], nxt_RX_PB_WM_XON[9][4][9:6], RX_PB_WM[9][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][5][0], nxt_RX_PB_WM_XON[9][5][5:0], RX_PB_WM[9][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][5][1], nxt_RX_PB_WM_XON[9][5][9:6], RX_PB_WM[9][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][6][0], nxt_RX_PB_WM_XON[9][6][5:0], RX_PB_WM[9][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][6][1], nxt_RX_PB_WM_XON[9][6][9:6], RX_PB_WM[9][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[9][7][0], nxt_RX_PB_WM_XON[9][7][5:0], RX_PB_WM[9][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[9][7][1], nxt_RX_PB_WM_XON[9][7][9:6], RX_PB_WM[9][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][0][0], nxt_RX_PB_WM_XON[10][0][5:0], RX_PB_WM[10][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][0][1], nxt_RX_PB_WM_XON[10][0][9:6], RX_PB_WM[10][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][1][0], nxt_RX_PB_WM_XON[10][1][5:0], RX_PB_WM[10][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][1][1], nxt_RX_PB_WM_XON[10][1][9:6], RX_PB_WM[10][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][2][0], nxt_RX_PB_WM_XON[10][2][5:0], RX_PB_WM[10][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][2][1], nxt_RX_PB_WM_XON[10][2][9:6], RX_PB_WM[10][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][3][0], nxt_RX_PB_WM_XON[10][3][5:0], RX_PB_WM[10][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][3][1], nxt_RX_PB_WM_XON[10][3][9:6], RX_PB_WM[10][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][4][0], nxt_RX_PB_WM_XON[10][4][5:0], RX_PB_WM[10][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][4][1], nxt_RX_PB_WM_XON[10][4][9:6], RX_PB_WM[10][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][5][0], nxt_RX_PB_WM_XON[10][5][5:0], RX_PB_WM[10][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][5][1], nxt_RX_PB_WM_XON[10][5][9:6], RX_PB_WM[10][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][6][0], nxt_RX_PB_WM_XON[10][6][5:0], RX_PB_WM[10][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][6][1], nxt_RX_PB_WM_XON[10][6][9:6], RX_PB_WM[10][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[10][7][0], nxt_RX_PB_WM_XON[10][7][5:0], RX_PB_WM[10][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[10][7][1], nxt_RX_PB_WM_XON[10][7][9:6], RX_PB_WM[10][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][0][0], nxt_RX_PB_WM_XON[11][0][5:0], RX_PB_WM[11][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][0][1], nxt_RX_PB_WM_XON[11][0][9:6], RX_PB_WM[11][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][1][0], nxt_RX_PB_WM_XON[11][1][5:0], RX_PB_WM[11][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][1][1], nxt_RX_PB_WM_XON[11][1][9:6], RX_PB_WM[11][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][2][0], nxt_RX_PB_WM_XON[11][2][5:0], RX_PB_WM[11][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][2][1], nxt_RX_PB_WM_XON[11][2][9:6], RX_PB_WM[11][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][3][0], nxt_RX_PB_WM_XON[11][3][5:0], RX_PB_WM[11][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][3][1], nxt_RX_PB_WM_XON[11][3][9:6], RX_PB_WM[11][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][4][0], nxt_RX_PB_WM_XON[11][4][5:0], RX_PB_WM[11][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][4][1], nxt_RX_PB_WM_XON[11][4][9:6], RX_PB_WM[11][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][5][0], nxt_RX_PB_WM_XON[11][5][5:0], RX_PB_WM[11][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][5][1], nxt_RX_PB_WM_XON[11][5][9:6], RX_PB_WM[11][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][6][0], nxt_RX_PB_WM_XON[11][6][5:0], RX_PB_WM[11][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][6][1], nxt_RX_PB_WM_XON[11][6][9:6], RX_PB_WM[11][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[11][7][0], nxt_RX_PB_WM_XON[11][7][5:0], RX_PB_WM[11][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[11][7][1], nxt_RX_PB_WM_XON[11][7][9:6], RX_PB_WM[11][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][0][0], nxt_RX_PB_WM_XON[12][0][5:0], RX_PB_WM[12][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][0][1], nxt_RX_PB_WM_XON[12][0][9:6], RX_PB_WM[12][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][1][0], nxt_RX_PB_WM_XON[12][1][5:0], RX_PB_WM[12][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][1][1], nxt_RX_PB_WM_XON[12][1][9:6], RX_PB_WM[12][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][2][0], nxt_RX_PB_WM_XON[12][2][5:0], RX_PB_WM[12][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][2][1], nxt_RX_PB_WM_XON[12][2][9:6], RX_PB_WM[12][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][3][0], nxt_RX_PB_WM_XON[12][3][5:0], RX_PB_WM[12][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][3][1], nxt_RX_PB_WM_XON[12][3][9:6], RX_PB_WM[12][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][4][0], nxt_RX_PB_WM_XON[12][4][5:0], RX_PB_WM[12][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][4][1], nxt_RX_PB_WM_XON[12][4][9:6], RX_PB_WM[12][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][5][0], nxt_RX_PB_WM_XON[12][5][5:0], RX_PB_WM[12][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][5][1], nxt_RX_PB_WM_XON[12][5][9:6], RX_PB_WM[12][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][6][0], nxt_RX_PB_WM_XON[12][6][5:0], RX_PB_WM[12][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][6][1], nxt_RX_PB_WM_XON[12][6][9:6], RX_PB_WM[12][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[12][7][0], nxt_RX_PB_WM_XON[12][7][5:0], RX_PB_WM[12][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[12][7][1], nxt_RX_PB_WM_XON[12][7][9:6], RX_PB_WM[12][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][0][0], nxt_RX_PB_WM_XON[13][0][5:0], RX_PB_WM[13][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][0][1], nxt_RX_PB_WM_XON[13][0][9:6], RX_PB_WM[13][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][1][0], nxt_RX_PB_WM_XON[13][1][5:0], RX_PB_WM[13][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][1][1], nxt_RX_PB_WM_XON[13][1][9:6], RX_PB_WM[13][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][2][0], nxt_RX_PB_WM_XON[13][2][5:0], RX_PB_WM[13][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][2][1], nxt_RX_PB_WM_XON[13][2][9:6], RX_PB_WM[13][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][3][0], nxt_RX_PB_WM_XON[13][3][5:0], RX_PB_WM[13][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][3][1], nxt_RX_PB_WM_XON[13][3][9:6], RX_PB_WM[13][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][4][0], nxt_RX_PB_WM_XON[13][4][5:0], RX_PB_WM[13][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][4][1], nxt_RX_PB_WM_XON[13][4][9:6], RX_PB_WM[13][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][5][0], nxt_RX_PB_WM_XON[13][5][5:0], RX_PB_WM[13][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][5][1], nxt_RX_PB_WM_XON[13][5][9:6], RX_PB_WM[13][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][6][0], nxt_RX_PB_WM_XON[13][6][5:0], RX_PB_WM[13][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][6][1], nxt_RX_PB_WM_XON[13][6][9:6], RX_PB_WM[13][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[13][7][0], nxt_RX_PB_WM_XON[13][7][5:0], RX_PB_WM[13][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[13][7][1], nxt_RX_PB_WM_XON[13][7][9:6], RX_PB_WM[13][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][0][0], nxt_RX_PB_WM_XON[14][0][5:0], RX_PB_WM[14][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][0][1], nxt_RX_PB_WM_XON[14][0][9:6], RX_PB_WM[14][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][1][0], nxt_RX_PB_WM_XON[14][1][5:0], RX_PB_WM[14][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][1][1], nxt_RX_PB_WM_XON[14][1][9:6], RX_PB_WM[14][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][2][0], nxt_RX_PB_WM_XON[14][2][5:0], RX_PB_WM[14][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][2][1], nxt_RX_PB_WM_XON[14][2][9:6], RX_PB_WM[14][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][3][0], nxt_RX_PB_WM_XON[14][3][5:0], RX_PB_WM[14][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][3][1], nxt_RX_PB_WM_XON[14][3][9:6], RX_PB_WM[14][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][4][0], nxt_RX_PB_WM_XON[14][4][5:0], RX_PB_WM[14][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][4][1], nxt_RX_PB_WM_XON[14][4][9:6], RX_PB_WM[14][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][5][0], nxt_RX_PB_WM_XON[14][5][5:0], RX_PB_WM[14][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][5][1], nxt_RX_PB_WM_XON[14][5][9:6], RX_PB_WM[14][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][6][0], nxt_RX_PB_WM_XON[14][6][5:0], RX_PB_WM[14][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][6][1], nxt_RX_PB_WM_XON[14][6][9:6], RX_PB_WM[14][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[14][7][0], nxt_RX_PB_WM_XON[14][7][5:0], RX_PB_WM[14][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[14][7][1], nxt_RX_PB_WM_XON[14][7][9:6], RX_PB_WM[14][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][0][0], nxt_RX_PB_WM_XON[15][0][5:0], RX_PB_WM[15][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][0][1], nxt_RX_PB_WM_XON[15][0][9:6], RX_PB_WM[15][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][1][0], nxt_RX_PB_WM_XON[15][1][5:0], RX_PB_WM[15][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][1][1], nxt_RX_PB_WM_XON[15][1][9:6], RX_PB_WM[15][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][2][0], nxt_RX_PB_WM_XON[15][2][5:0], RX_PB_WM[15][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][2][1], nxt_RX_PB_WM_XON[15][2][9:6], RX_PB_WM[15][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][3][0], nxt_RX_PB_WM_XON[15][3][5:0], RX_PB_WM[15][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][3][1], nxt_RX_PB_WM_XON[15][3][9:6], RX_PB_WM[15][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][4][0], nxt_RX_PB_WM_XON[15][4][5:0], RX_PB_WM[15][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][4][1], nxt_RX_PB_WM_XON[15][4][9:6], RX_PB_WM[15][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][5][0], nxt_RX_PB_WM_XON[15][5][5:0], RX_PB_WM[15][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][5][1], nxt_RX_PB_WM_XON[15][5][9:6], RX_PB_WM[15][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][6][0], nxt_RX_PB_WM_XON[15][6][5:0], RX_PB_WM[15][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][6][1], nxt_RX_PB_WM_XON[15][6][9:6], RX_PB_WM[15][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[15][7][0], nxt_RX_PB_WM_XON[15][7][5:0], RX_PB_WM[15][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[15][7][1], nxt_RX_PB_WM_XON[15][7][9:6], RX_PB_WM[15][7].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][0][0], nxt_RX_PB_WM_XON[16][0][5:0], RX_PB_WM[16][0].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][0][1], nxt_RX_PB_WM_XON[16][0][9:6], RX_PB_WM[16][0].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][1][0], nxt_RX_PB_WM_XON[16][1][5:0], RX_PB_WM[16][1].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][1][1], nxt_RX_PB_WM_XON[16][1][9:6], RX_PB_WM[16][1].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][2][0], nxt_RX_PB_WM_XON[16][2][5:0], RX_PB_WM[16][2].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][2][1], nxt_RX_PB_WM_XON[16][2][9:6], RX_PB_WM[16][2].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][3][0], nxt_RX_PB_WM_XON[16][3][5:0], RX_PB_WM[16][3].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][3][1], nxt_RX_PB_WM_XON[16][3][9:6], RX_PB_WM[16][3].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][4][0], nxt_RX_PB_WM_XON[16][4][5:0], RX_PB_WM[16][4].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][4][1], nxt_RX_PB_WM_XON[16][4][9:6], RX_PB_WM[16][4].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][5][0], nxt_RX_PB_WM_XON[16][5][5:0], RX_PB_WM[16][5].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][5][1], nxt_RX_PB_WM_XON[16][5][9:6], RX_PB_WM[16][5].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][6][0], nxt_RX_PB_WM_XON[16][6][5:0], RX_PB_WM[16][6].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][6][1], nxt_RX_PB_WM_XON[16][6][9:6], RX_PB_WM[16][6].XON[9:6])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 6'h0, up_RX_PB_WM_XON[16][7][0], nxt_RX_PB_WM_XON[16][7][5:0], RX_PB_WM[16][7].XON[5:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 4'h8, up_RX_PB_WM_XON[16][7][1], nxt_RX_PB_WM_XON[16][7][9:6], RX_PB_WM[16][7].XON[9:6])

// ----------------------------------------------------------------------
// RX_PB_WM.LOSSLESS x1 RW, using RW template.
logic [16:0][7:0][0:0] up_RX_PB_WM_LOSSLESS;
always_comb begin
 up_RX_PB_WM_LOSSLESS[0][0] =
    ({1{write_req_RX_PB_WM[0][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[0][1] =
    ({1{write_req_RX_PB_WM[0][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[0][2] =
    ({1{write_req_RX_PB_WM[0][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[0][3] =
    ({1{write_req_RX_PB_WM[0][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[0][4] =
    ({1{write_req_RX_PB_WM[0][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[0][5] =
    ({1{write_req_RX_PB_WM[0][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[0][6] =
    ({1{write_req_RX_PB_WM[0][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[0][7] =
    ({1{write_req_RX_PB_WM[0][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][0] =
    ({1{write_req_RX_PB_WM[1][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][1] =
    ({1{write_req_RX_PB_WM[1][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][2] =
    ({1{write_req_RX_PB_WM[1][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][3] =
    ({1{write_req_RX_PB_WM[1][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][4] =
    ({1{write_req_RX_PB_WM[1][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][5] =
    ({1{write_req_RX_PB_WM[1][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][6] =
    ({1{write_req_RX_PB_WM[1][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[1][7] =
    ({1{write_req_RX_PB_WM[1][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][0] =
    ({1{write_req_RX_PB_WM[2][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][1] =
    ({1{write_req_RX_PB_WM[2][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][2] =
    ({1{write_req_RX_PB_WM[2][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][3] =
    ({1{write_req_RX_PB_WM[2][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][4] =
    ({1{write_req_RX_PB_WM[2][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][5] =
    ({1{write_req_RX_PB_WM[2][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][6] =
    ({1{write_req_RX_PB_WM[2][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[2][7] =
    ({1{write_req_RX_PB_WM[2][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][0] =
    ({1{write_req_RX_PB_WM[3][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][1] =
    ({1{write_req_RX_PB_WM[3][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][2] =
    ({1{write_req_RX_PB_WM[3][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][3] =
    ({1{write_req_RX_PB_WM[3][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][4] =
    ({1{write_req_RX_PB_WM[3][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][5] =
    ({1{write_req_RX_PB_WM[3][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][6] =
    ({1{write_req_RX_PB_WM[3][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[3][7] =
    ({1{write_req_RX_PB_WM[3][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][0] =
    ({1{write_req_RX_PB_WM[4][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][1] =
    ({1{write_req_RX_PB_WM[4][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][2] =
    ({1{write_req_RX_PB_WM[4][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][3] =
    ({1{write_req_RX_PB_WM[4][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][4] =
    ({1{write_req_RX_PB_WM[4][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][5] =
    ({1{write_req_RX_PB_WM[4][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][6] =
    ({1{write_req_RX_PB_WM[4][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[4][7] =
    ({1{write_req_RX_PB_WM[4][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][0] =
    ({1{write_req_RX_PB_WM[5][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][1] =
    ({1{write_req_RX_PB_WM[5][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][2] =
    ({1{write_req_RX_PB_WM[5][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][3] =
    ({1{write_req_RX_PB_WM[5][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][4] =
    ({1{write_req_RX_PB_WM[5][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][5] =
    ({1{write_req_RX_PB_WM[5][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][6] =
    ({1{write_req_RX_PB_WM[5][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[5][7] =
    ({1{write_req_RX_PB_WM[5][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][0] =
    ({1{write_req_RX_PB_WM[6][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][1] =
    ({1{write_req_RX_PB_WM[6][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][2] =
    ({1{write_req_RX_PB_WM[6][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][3] =
    ({1{write_req_RX_PB_WM[6][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][4] =
    ({1{write_req_RX_PB_WM[6][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][5] =
    ({1{write_req_RX_PB_WM[6][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][6] =
    ({1{write_req_RX_PB_WM[6][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[6][7] =
    ({1{write_req_RX_PB_WM[6][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][0] =
    ({1{write_req_RX_PB_WM[7][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][1] =
    ({1{write_req_RX_PB_WM[7][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][2] =
    ({1{write_req_RX_PB_WM[7][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][3] =
    ({1{write_req_RX_PB_WM[7][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][4] =
    ({1{write_req_RX_PB_WM[7][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][5] =
    ({1{write_req_RX_PB_WM[7][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][6] =
    ({1{write_req_RX_PB_WM[7][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[7][7] =
    ({1{write_req_RX_PB_WM[7][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][0] =
    ({1{write_req_RX_PB_WM[8][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][1] =
    ({1{write_req_RX_PB_WM[8][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][2] =
    ({1{write_req_RX_PB_WM[8][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][3] =
    ({1{write_req_RX_PB_WM[8][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][4] =
    ({1{write_req_RX_PB_WM[8][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][5] =
    ({1{write_req_RX_PB_WM[8][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][6] =
    ({1{write_req_RX_PB_WM[8][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[8][7] =
    ({1{write_req_RX_PB_WM[8][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][0] =
    ({1{write_req_RX_PB_WM[9][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][1] =
    ({1{write_req_RX_PB_WM[9][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][2] =
    ({1{write_req_RX_PB_WM[9][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][3] =
    ({1{write_req_RX_PB_WM[9][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][4] =
    ({1{write_req_RX_PB_WM[9][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][5] =
    ({1{write_req_RX_PB_WM[9][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][6] =
    ({1{write_req_RX_PB_WM[9][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[9][7] =
    ({1{write_req_RX_PB_WM[9][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][0] =
    ({1{write_req_RX_PB_WM[10][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][1] =
    ({1{write_req_RX_PB_WM[10][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][2] =
    ({1{write_req_RX_PB_WM[10][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][3] =
    ({1{write_req_RX_PB_WM[10][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][4] =
    ({1{write_req_RX_PB_WM[10][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][5] =
    ({1{write_req_RX_PB_WM[10][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][6] =
    ({1{write_req_RX_PB_WM[10][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[10][7] =
    ({1{write_req_RX_PB_WM[10][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][0] =
    ({1{write_req_RX_PB_WM[11][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][1] =
    ({1{write_req_RX_PB_WM[11][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][2] =
    ({1{write_req_RX_PB_WM[11][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][3] =
    ({1{write_req_RX_PB_WM[11][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][4] =
    ({1{write_req_RX_PB_WM[11][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][5] =
    ({1{write_req_RX_PB_WM[11][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][6] =
    ({1{write_req_RX_PB_WM[11][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[11][7] =
    ({1{write_req_RX_PB_WM[11][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][0] =
    ({1{write_req_RX_PB_WM[12][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][1] =
    ({1{write_req_RX_PB_WM[12][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][2] =
    ({1{write_req_RX_PB_WM[12][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][3] =
    ({1{write_req_RX_PB_WM[12][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][4] =
    ({1{write_req_RX_PB_WM[12][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][5] =
    ({1{write_req_RX_PB_WM[12][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][6] =
    ({1{write_req_RX_PB_WM[12][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[12][7] =
    ({1{write_req_RX_PB_WM[12][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][0] =
    ({1{write_req_RX_PB_WM[13][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][1] =
    ({1{write_req_RX_PB_WM[13][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][2] =
    ({1{write_req_RX_PB_WM[13][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][3] =
    ({1{write_req_RX_PB_WM[13][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][4] =
    ({1{write_req_RX_PB_WM[13][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][5] =
    ({1{write_req_RX_PB_WM[13][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][6] =
    ({1{write_req_RX_PB_WM[13][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[13][7] =
    ({1{write_req_RX_PB_WM[13][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][0] =
    ({1{write_req_RX_PB_WM[14][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][1] =
    ({1{write_req_RX_PB_WM[14][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][2] =
    ({1{write_req_RX_PB_WM[14][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][3] =
    ({1{write_req_RX_PB_WM[14][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][4] =
    ({1{write_req_RX_PB_WM[14][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][5] =
    ({1{write_req_RX_PB_WM[14][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][6] =
    ({1{write_req_RX_PB_WM[14][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[14][7] =
    ({1{write_req_RX_PB_WM[14][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][0] =
    ({1{write_req_RX_PB_WM[15][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][1] =
    ({1{write_req_RX_PB_WM[15][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][2] =
    ({1{write_req_RX_PB_WM[15][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][3] =
    ({1{write_req_RX_PB_WM[15][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][4] =
    ({1{write_req_RX_PB_WM[15][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][5] =
    ({1{write_req_RX_PB_WM[15][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][6] =
    ({1{write_req_RX_PB_WM[15][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[15][7] =
    ({1{write_req_RX_PB_WM[15][7] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][0] =
    ({1{write_req_RX_PB_WM[16][0] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][1] =
    ({1{write_req_RX_PB_WM[16][1] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][2] =
    ({1{write_req_RX_PB_WM[16][2] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][3] =
    ({1{write_req_RX_PB_WM[16][3] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][4] =
    ({1{write_req_RX_PB_WM[16][4] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][5] =
    ({1{write_req_RX_PB_WM[16][5] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][6] =
    ({1{write_req_RX_PB_WM[16][6] }} &
    be[2:2]);
 up_RX_PB_WM_LOSSLESS[16][7] =
    ({1{write_req_RX_PB_WM[16][7] }} &
    be[2:2]);
end

logic [16:0][7:0][0:0] nxt_RX_PB_WM_LOSSLESS;
always_comb begin
 nxt_RX_PB_WM_LOSSLESS[0][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[0][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[0][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[0][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[0][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[0][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[0][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[0][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[1][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[2][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[3][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[4][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[5][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[6][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[7][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[8][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[9][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[10][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[11][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[12][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[13][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[14][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[15][7] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][0] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][1] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][2] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][3] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][4] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][5] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][6] = write_data[20:20];

 nxt_RX_PB_WM_LOSSLESS[16][7] = write_data[20:20];

end


`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][0][0], nxt_RX_PB_WM_LOSSLESS[0][0][0:0], RX_PB_WM[0][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][1][0], nxt_RX_PB_WM_LOSSLESS[0][1][0:0], RX_PB_WM[0][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][2][0], nxt_RX_PB_WM_LOSSLESS[0][2][0:0], RX_PB_WM[0][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][3][0], nxt_RX_PB_WM_LOSSLESS[0][3][0:0], RX_PB_WM[0][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][4][0], nxt_RX_PB_WM_LOSSLESS[0][4][0:0], RX_PB_WM[0][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][5][0], nxt_RX_PB_WM_LOSSLESS[0][5][0:0], RX_PB_WM[0][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][6][0], nxt_RX_PB_WM_LOSSLESS[0][6][0:0], RX_PB_WM[0][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[0][7][0], nxt_RX_PB_WM_LOSSLESS[0][7][0:0], RX_PB_WM[0][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][0][0], nxt_RX_PB_WM_LOSSLESS[1][0][0:0], RX_PB_WM[1][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][1][0], nxt_RX_PB_WM_LOSSLESS[1][1][0:0], RX_PB_WM[1][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][2][0], nxt_RX_PB_WM_LOSSLESS[1][2][0:0], RX_PB_WM[1][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][3][0], nxt_RX_PB_WM_LOSSLESS[1][3][0:0], RX_PB_WM[1][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][4][0], nxt_RX_PB_WM_LOSSLESS[1][4][0:0], RX_PB_WM[1][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][5][0], nxt_RX_PB_WM_LOSSLESS[1][5][0:0], RX_PB_WM[1][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][6][0], nxt_RX_PB_WM_LOSSLESS[1][6][0:0], RX_PB_WM[1][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[1][7][0], nxt_RX_PB_WM_LOSSLESS[1][7][0:0], RX_PB_WM[1][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][0][0], nxt_RX_PB_WM_LOSSLESS[2][0][0:0], RX_PB_WM[2][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][1][0], nxt_RX_PB_WM_LOSSLESS[2][1][0:0], RX_PB_WM[2][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][2][0], nxt_RX_PB_WM_LOSSLESS[2][2][0:0], RX_PB_WM[2][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][3][0], nxt_RX_PB_WM_LOSSLESS[2][3][0:0], RX_PB_WM[2][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][4][0], nxt_RX_PB_WM_LOSSLESS[2][4][0:0], RX_PB_WM[2][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][5][0], nxt_RX_PB_WM_LOSSLESS[2][5][0:0], RX_PB_WM[2][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][6][0], nxt_RX_PB_WM_LOSSLESS[2][6][0:0], RX_PB_WM[2][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[2][7][0], nxt_RX_PB_WM_LOSSLESS[2][7][0:0], RX_PB_WM[2][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][0][0], nxt_RX_PB_WM_LOSSLESS[3][0][0:0], RX_PB_WM[3][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][1][0], nxt_RX_PB_WM_LOSSLESS[3][1][0:0], RX_PB_WM[3][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][2][0], nxt_RX_PB_WM_LOSSLESS[3][2][0:0], RX_PB_WM[3][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][3][0], nxt_RX_PB_WM_LOSSLESS[3][3][0:0], RX_PB_WM[3][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][4][0], nxt_RX_PB_WM_LOSSLESS[3][4][0:0], RX_PB_WM[3][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][5][0], nxt_RX_PB_WM_LOSSLESS[3][5][0:0], RX_PB_WM[3][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][6][0], nxt_RX_PB_WM_LOSSLESS[3][6][0:0], RX_PB_WM[3][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[3][7][0], nxt_RX_PB_WM_LOSSLESS[3][7][0:0], RX_PB_WM[3][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][0][0], nxt_RX_PB_WM_LOSSLESS[4][0][0:0], RX_PB_WM[4][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][1][0], nxt_RX_PB_WM_LOSSLESS[4][1][0:0], RX_PB_WM[4][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][2][0], nxt_RX_PB_WM_LOSSLESS[4][2][0:0], RX_PB_WM[4][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][3][0], nxt_RX_PB_WM_LOSSLESS[4][3][0:0], RX_PB_WM[4][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][4][0], nxt_RX_PB_WM_LOSSLESS[4][4][0:0], RX_PB_WM[4][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][5][0], nxt_RX_PB_WM_LOSSLESS[4][5][0:0], RX_PB_WM[4][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][6][0], nxt_RX_PB_WM_LOSSLESS[4][6][0:0], RX_PB_WM[4][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[4][7][0], nxt_RX_PB_WM_LOSSLESS[4][7][0:0], RX_PB_WM[4][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][0][0], nxt_RX_PB_WM_LOSSLESS[5][0][0:0], RX_PB_WM[5][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][1][0], nxt_RX_PB_WM_LOSSLESS[5][1][0:0], RX_PB_WM[5][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][2][0], nxt_RX_PB_WM_LOSSLESS[5][2][0:0], RX_PB_WM[5][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][3][0], nxt_RX_PB_WM_LOSSLESS[5][3][0:0], RX_PB_WM[5][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][4][0], nxt_RX_PB_WM_LOSSLESS[5][4][0:0], RX_PB_WM[5][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][5][0], nxt_RX_PB_WM_LOSSLESS[5][5][0:0], RX_PB_WM[5][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][6][0], nxt_RX_PB_WM_LOSSLESS[5][6][0:0], RX_PB_WM[5][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[5][7][0], nxt_RX_PB_WM_LOSSLESS[5][7][0:0], RX_PB_WM[5][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][0][0], nxt_RX_PB_WM_LOSSLESS[6][0][0:0], RX_PB_WM[6][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][1][0], nxt_RX_PB_WM_LOSSLESS[6][1][0:0], RX_PB_WM[6][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][2][0], nxt_RX_PB_WM_LOSSLESS[6][2][0:0], RX_PB_WM[6][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][3][0], nxt_RX_PB_WM_LOSSLESS[6][3][0:0], RX_PB_WM[6][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][4][0], nxt_RX_PB_WM_LOSSLESS[6][4][0:0], RX_PB_WM[6][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][5][0], nxt_RX_PB_WM_LOSSLESS[6][5][0:0], RX_PB_WM[6][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][6][0], nxt_RX_PB_WM_LOSSLESS[6][6][0:0], RX_PB_WM[6][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[6][7][0], nxt_RX_PB_WM_LOSSLESS[6][7][0:0], RX_PB_WM[6][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][0][0], nxt_RX_PB_WM_LOSSLESS[7][0][0:0], RX_PB_WM[7][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][1][0], nxt_RX_PB_WM_LOSSLESS[7][1][0:0], RX_PB_WM[7][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][2][0], nxt_RX_PB_WM_LOSSLESS[7][2][0:0], RX_PB_WM[7][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][3][0], nxt_RX_PB_WM_LOSSLESS[7][3][0:0], RX_PB_WM[7][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][4][0], nxt_RX_PB_WM_LOSSLESS[7][4][0:0], RX_PB_WM[7][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][5][0], nxt_RX_PB_WM_LOSSLESS[7][5][0:0], RX_PB_WM[7][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][6][0], nxt_RX_PB_WM_LOSSLESS[7][6][0:0], RX_PB_WM[7][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[7][7][0], nxt_RX_PB_WM_LOSSLESS[7][7][0:0], RX_PB_WM[7][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][0][0], nxt_RX_PB_WM_LOSSLESS[8][0][0:0], RX_PB_WM[8][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][1][0], nxt_RX_PB_WM_LOSSLESS[8][1][0:0], RX_PB_WM[8][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][2][0], nxt_RX_PB_WM_LOSSLESS[8][2][0:0], RX_PB_WM[8][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][3][0], nxt_RX_PB_WM_LOSSLESS[8][3][0:0], RX_PB_WM[8][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][4][0], nxt_RX_PB_WM_LOSSLESS[8][4][0:0], RX_PB_WM[8][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][5][0], nxt_RX_PB_WM_LOSSLESS[8][5][0:0], RX_PB_WM[8][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][6][0], nxt_RX_PB_WM_LOSSLESS[8][6][0:0], RX_PB_WM[8][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[8][7][0], nxt_RX_PB_WM_LOSSLESS[8][7][0:0], RX_PB_WM[8][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][0][0], nxt_RX_PB_WM_LOSSLESS[9][0][0:0], RX_PB_WM[9][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][1][0], nxt_RX_PB_WM_LOSSLESS[9][1][0:0], RX_PB_WM[9][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][2][0], nxt_RX_PB_WM_LOSSLESS[9][2][0:0], RX_PB_WM[9][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][3][0], nxt_RX_PB_WM_LOSSLESS[9][3][0:0], RX_PB_WM[9][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][4][0], nxt_RX_PB_WM_LOSSLESS[9][4][0:0], RX_PB_WM[9][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][5][0], nxt_RX_PB_WM_LOSSLESS[9][5][0:0], RX_PB_WM[9][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][6][0], nxt_RX_PB_WM_LOSSLESS[9][6][0:0], RX_PB_WM[9][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[9][7][0], nxt_RX_PB_WM_LOSSLESS[9][7][0:0], RX_PB_WM[9][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][0][0], nxt_RX_PB_WM_LOSSLESS[10][0][0:0], RX_PB_WM[10][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][1][0], nxt_RX_PB_WM_LOSSLESS[10][1][0:0], RX_PB_WM[10][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][2][0], nxt_RX_PB_WM_LOSSLESS[10][2][0:0], RX_PB_WM[10][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][3][0], nxt_RX_PB_WM_LOSSLESS[10][3][0:0], RX_PB_WM[10][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][4][0], nxt_RX_PB_WM_LOSSLESS[10][4][0:0], RX_PB_WM[10][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][5][0], nxt_RX_PB_WM_LOSSLESS[10][5][0:0], RX_PB_WM[10][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][6][0], nxt_RX_PB_WM_LOSSLESS[10][6][0:0], RX_PB_WM[10][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[10][7][0], nxt_RX_PB_WM_LOSSLESS[10][7][0:0], RX_PB_WM[10][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][0][0], nxt_RX_PB_WM_LOSSLESS[11][0][0:0], RX_PB_WM[11][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][1][0], nxt_RX_PB_WM_LOSSLESS[11][1][0:0], RX_PB_WM[11][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][2][0], nxt_RX_PB_WM_LOSSLESS[11][2][0:0], RX_PB_WM[11][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][3][0], nxt_RX_PB_WM_LOSSLESS[11][3][0:0], RX_PB_WM[11][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][4][0], nxt_RX_PB_WM_LOSSLESS[11][4][0:0], RX_PB_WM[11][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][5][0], nxt_RX_PB_WM_LOSSLESS[11][5][0:0], RX_PB_WM[11][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][6][0], nxt_RX_PB_WM_LOSSLESS[11][6][0:0], RX_PB_WM[11][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[11][7][0], nxt_RX_PB_WM_LOSSLESS[11][7][0:0], RX_PB_WM[11][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][0][0], nxt_RX_PB_WM_LOSSLESS[12][0][0:0], RX_PB_WM[12][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][1][0], nxt_RX_PB_WM_LOSSLESS[12][1][0:0], RX_PB_WM[12][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][2][0], nxt_RX_PB_WM_LOSSLESS[12][2][0:0], RX_PB_WM[12][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][3][0], nxt_RX_PB_WM_LOSSLESS[12][3][0:0], RX_PB_WM[12][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][4][0], nxt_RX_PB_WM_LOSSLESS[12][4][0:0], RX_PB_WM[12][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][5][0], nxt_RX_PB_WM_LOSSLESS[12][5][0:0], RX_PB_WM[12][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][6][0], nxt_RX_PB_WM_LOSSLESS[12][6][0:0], RX_PB_WM[12][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[12][7][0], nxt_RX_PB_WM_LOSSLESS[12][7][0:0], RX_PB_WM[12][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][0][0], nxt_RX_PB_WM_LOSSLESS[13][0][0:0], RX_PB_WM[13][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][1][0], nxt_RX_PB_WM_LOSSLESS[13][1][0:0], RX_PB_WM[13][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][2][0], nxt_RX_PB_WM_LOSSLESS[13][2][0:0], RX_PB_WM[13][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][3][0], nxt_RX_PB_WM_LOSSLESS[13][3][0:0], RX_PB_WM[13][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][4][0], nxt_RX_PB_WM_LOSSLESS[13][4][0:0], RX_PB_WM[13][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][5][0], nxt_RX_PB_WM_LOSSLESS[13][5][0:0], RX_PB_WM[13][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][6][0], nxt_RX_PB_WM_LOSSLESS[13][6][0:0], RX_PB_WM[13][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[13][7][0], nxt_RX_PB_WM_LOSSLESS[13][7][0:0], RX_PB_WM[13][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][0][0], nxt_RX_PB_WM_LOSSLESS[14][0][0:0], RX_PB_WM[14][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][1][0], nxt_RX_PB_WM_LOSSLESS[14][1][0:0], RX_PB_WM[14][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][2][0], nxt_RX_PB_WM_LOSSLESS[14][2][0:0], RX_PB_WM[14][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][3][0], nxt_RX_PB_WM_LOSSLESS[14][3][0:0], RX_PB_WM[14][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][4][0], nxt_RX_PB_WM_LOSSLESS[14][4][0:0], RX_PB_WM[14][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][5][0], nxt_RX_PB_WM_LOSSLESS[14][5][0:0], RX_PB_WM[14][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][6][0], nxt_RX_PB_WM_LOSSLESS[14][6][0:0], RX_PB_WM[14][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[14][7][0], nxt_RX_PB_WM_LOSSLESS[14][7][0:0], RX_PB_WM[14][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][0][0], nxt_RX_PB_WM_LOSSLESS[15][0][0:0], RX_PB_WM[15][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][1][0], nxt_RX_PB_WM_LOSSLESS[15][1][0:0], RX_PB_WM[15][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][2][0], nxt_RX_PB_WM_LOSSLESS[15][2][0:0], RX_PB_WM[15][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][3][0], nxt_RX_PB_WM_LOSSLESS[15][3][0:0], RX_PB_WM[15][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][4][0], nxt_RX_PB_WM_LOSSLESS[15][4][0:0], RX_PB_WM[15][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][5][0], nxt_RX_PB_WM_LOSSLESS[15][5][0:0], RX_PB_WM[15][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][6][0], nxt_RX_PB_WM_LOSSLESS[15][6][0:0], RX_PB_WM[15][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[15][7][0], nxt_RX_PB_WM_LOSSLESS[15][7][0:0], RX_PB_WM[15][7].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][0][0], nxt_RX_PB_WM_LOSSLESS[16][0][0:0], RX_PB_WM[16][0].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][1][0], nxt_RX_PB_WM_LOSSLESS[16][1][0:0], RX_PB_WM[16][1].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][2][0], nxt_RX_PB_WM_LOSSLESS[16][2][0:0], RX_PB_WM[16][2].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][3][0], nxt_RX_PB_WM_LOSSLESS[16][3][0:0], RX_PB_WM[16][3].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][4][0], nxt_RX_PB_WM_LOSSLESS[16][4][0:0], RX_PB_WM[16][4].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][5][0], nxt_RX_PB_WM_LOSSLESS[16][5][0:0], RX_PB_WM[16][5].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][6][0], nxt_RX_PB_WM_LOSSLESS[16][6][0:0], RX_PB_WM[16][6].LOSSLESS[0:0])
`RTLGEN_MBY_RX_PB_EN_FF(gated_clk, rst_n, 1'h0, up_RX_PB_WM_LOSSLESS[16][7][0], nxt_RX_PB_WM_LOSSLESS[16][7][0:0], RX_PB_WM[16][7].LOSSLESS[0:0])
// Shared registers assignments


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_RX_PB_MEM) 
           RX_PB_PORT_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_RX_PB_MEM) 
           RX_PB_PORT_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_RX_PB_MEM) 
           RX_PB_PORT_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_PORT_CFG};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[0][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[0][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[1][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[1][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[2][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[2][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[3][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[3][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[4][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[4][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[5][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[5][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[6][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[6][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[7][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[7][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[8][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[8][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[9][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[9][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[10][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[10][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[11][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[11][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[12][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[12][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[13][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[13][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[14][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[14][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[15][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[15][7]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][0]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][0]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][1]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][1]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][2]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][2]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][3]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][3]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][4]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][4]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][5]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][5]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][6]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][6]};
                 default: read_data = '0;
              endcase
           end
           RX_PB_WM_DECODE_ADDR[16][7]: begin
              unique casez ({req_fid,req_bar})
                 {MBY_RX_PB_MAP_SB_FID,MBY_RX_PB_MAP_SB_BAR}: read_data = {RX_PB_WM[16][7]};
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    RX_PB_PORT_CFG.reserved0 = '0;
    RX_PB_WM[0][0].reserved0 = '0;
    RX_PB_WM[0][1].reserved0 = '0;
    RX_PB_WM[0][2].reserved0 = '0;
    RX_PB_WM[0][3].reserved0 = '0;
    RX_PB_WM[0][4].reserved0 = '0;
    RX_PB_WM[0][5].reserved0 = '0;
    RX_PB_WM[0][6].reserved0 = '0;
    RX_PB_WM[0][7].reserved0 = '0;
    RX_PB_WM[1][0].reserved0 = '0;
    RX_PB_WM[1][1].reserved0 = '0;
    RX_PB_WM[1][2].reserved0 = '0;
    RX_PB_WM[1][3].reserved0 = '0;
    RX_PB_WM[1][4].reserved0 = '0;
    RX_PB_WM[1][5].reserved0 = '0;
    RX_PB_WM[1][6].reserved0 = '0;
    RX_PB_WM[1][7].reserved0 = '0;
    RX_PB_WM[2][0].reserved0 = '0;
    RX_PB_WM[2][1].reserved0 = '0;
    RX_PB_WM[2][2].reserved0 = '0;
    RX_PB_WM[2][3].reserved0 = '0;
    RX_PB_WM[2][4].reserved0 = '0;
    RX_PB_WM[2][5].reserved0 = '0;
    RX_PB_WM[2][6].reserved0 = '0;
    RX_PB_WM[2][7].reserved0 = '0;
    RX_PB_WM[3][0].reserved0 = '0;
    RX_PB_WM[3][1].reserved0 = '0;
    RX_PB_WM[3][2].reserved0 = '0;
    RX_PB_WM[3][3].reserved0 = '0;
    RX_PB_WM[3][4].reserved0 = '0;
    RX_PB_WM[3][5].reserved0 = '0;
    RX_PB_WM[3][6].reserved0 = '0;
    RX_PB_WM[3][7].reserved0 = '0;
    RX_PB_WM[4][0].reserved0 = '0;
    RX_PB_WM[4][1].reserved0 = '0;
    RX_PB_WM[4][2].reserved0 = '0;
    RX_PB_WM[4][3].reserved0 = '0;
    RX_PB_WM[4][4].reserved0 = '0;
    RX_PB_WM[4][5].reserved0 = '0;
    RX_PB_WM[4][6].reserved0 = '0;
    RX_PB_WM[4][7].reserved0 = '0;
    RX_PB_WM[5][0].reserved0 = '0;
    RX_PB_WM[5][1].reserved0 = '0;
    RX_PB_WM[5][2].reserved0 = '0;
    RX_PB_WM[5][3].reserved0 = '0;
    RX_PB_WM[5][4].reserved0 = '0;
    RX_PB_WM[5][5].reserved0 = '0;
    RX_PB_WM[5][6].reserved0 = '0;
    RX_PB_WM[5][7].reserved0 = '0;
    RX_PB_WM[6][0].reserved0 = '0;
    RX_PB_WM[6][1].reserved0 = '0;
    RX_PB_WM[6][2].reserved0 = '0;
    RX_PB_WM[6][3].reserved0 = '0;
    RX_PB_WM[6][4].reserved0 = '0;
    RX_PB_WM[6][5].reserved0 = '0;
    RX_PB_WM[6][6].reserved0 = '0;
    RX_PB_WM[6][7].reserved0 = '0;
    RX_PB_WM[7][0].reserved0 = '0;
    RX_PB_WM[7][1].reserved0 = '0;
    RX_PB_WM[7][2].reserved0 = '0;
    RX_PB_WM[7][3].reserved0 = '0;
    RX_PB_WM[7][4].reserved0 = '0;
    RX_PB_WM[7][5].reserved0 = '0;
    RX_PB_WM[7][6].reserved0 = '0;
    RX_PB_WM[7][7].reserved0 = '0;
    RX_PB_WM[8][0].reserved0 = '0;
    RX_PB_WM[8][1].reserved0 = '0;
    RX_PB_WM[8][2].reserved0 = '0;
    RX_PB_WM[8][3].reserved0 = '0;
    RX_PB_WM[8][4].reserved0 = '0;
    RX_PB_WM[8][5].reserved0 = '0;
    RX_PB_WM[8][6].reserved0 = '0;
    RX_PB_WM[8][7].reserved0 = '0;
    RX_PB_WM[9][0].reserved0 = '0;
    RX_PB_WM[9][1].reserved0 = '0;
    RX_PB_WM[9][2].reserved0 = '0;
    RX_PB_WM[9][3].reserved0 = '0;
    RX_PB_WM[9][4].reserved0 = '0;
    RX_PB_WM[9][5].reserved0 = '0;
    RX_PB_WM[9][6].reserved0 = '0;
    RX_PB_WM[9][7].reserved0 = '0;
    RX_PB_WM[10][0].reserved0 = '0;
    RX_PB_WM[10][1].reserved0 = '0;
    RX_PB_WM[10][2].reserved0 = '0;
    RX_PB_WM[10][3].reserved0 = '0;
    RX_PB_WM[10][4].reserved0 = '0;
    RX_PB_WM[10][5].reserved0 = '0;
    RX_PB_WM[10][6].reserved0 = '0;
    RX_PB_WM[10][7].reserved0 = '0;
    RX_PB_WM[11][0].reserved0 = '0;
    RX_PB_WM[11][1].reserved0 = '0;
    RX_PB_WM[11][2].reserved0 = '0;
    RX_PB_WM[11][3].reserved0 = '0;
    RX_PB_WM[11][4].reserved0 = '0;
    RX_PB_WM[11][5].reserved0 = '0;
    RX_PB_WM[11][6].reserved0 = '0;
    RX_PB_WM[11][7].reserved0 = '0;
    RX_PB_WM[12][0].reserved0 = '0;
    RX_PB_WM[12][1].reserved0 = '0;
    RX_PB_WM[12][2].reserved0 = '0;
    RX_PB_WM[12][3].reserved0 = '0;
    RX_PB_WM[12][4].reserved0 = '0;
    RX_PB_WM[12][5].reserved0 = '0;
    RX_PB_WM[12][6].reserved0 = '0;
    RX_PB_WM[12][7].reserved0 = '0;
    RX_PB_WM[13][0].reserved0 = '0;
    RX_PB_WM[13][1].reserved0 = '0;
    RX_PB_WM[13][2].reserved0 = '0;
    RX_PB_WM[13][3].reserved0 = '0;
    RX_PB_WM[13][4].reserved0 = '0;
    RX_PB_WM[13][5].reserved0 = '0;
    RX_PB_WM[13][6].reserved0 = '0;
    RX_PB_WM[13][7].reserved0 = '0;
    RX_PB_WM[14][0].reserved0 = '0;
    RX_PB_WM[14][1].reserved0 = '0;
    RX_PB_WM[14][2].reserved0 = '0;
    RX_PB_WM[14][3].reserved0 = '0;
    RX_PB_WM[14][4].reserved0 = '0;
    RX_PB_WM[14][5].reserved0 = '0;
    RX_PB_WM[14][6].reserved0 = '0;
    RX_PB_WM[14][7].reserved0 = '0;
    RX_PB_WM[15][0].reserved0 = '0;
    RX_PB_WM[15][1].reserved0 = '0;
    RX_PB_WM[15][2].reserved0 = '0;
    RX_PB_WM[15][3].reserved0 = '0;
    RX_PB_WM[15][4].reserved0 = '0;
    RX_PB_WM[15][5].reserved0 = '0;
    RX_PB_WM[15][6].reserved0 = '0;
    RX_PB_WM[15][7].reserved0 = '0;
    RX_PB_WM[16][0].reserved0 = '0;
    RX_PB_WM[16][1].reserved0 = '0;
    RX_PB_WM[16][2].reserved0 = '0;
    RX_PB_WM[16][3].reserved0 = '0;
    RX_PB_WM[16][4].reserved0 = '0;
    RX_PB_WM[16][5].reserved0 = '0;
    RX_PB_WM[16][6].reserved0 = '0;
    RX_PB_WM[16][7].reserved0 = '0;
end

// end register RSVD init section }


// ======================================================================
// begin unit parity section {


// end unit parity section }


endmodule
//lintra pop
//lintra pop
