package mby_mgp_bfm_pkg;

   `include "uvm_macros.svh"
   import uvm_pkg::*;
   import shdv_base_pkg::*;

   `include "mby_mgp_defines.svh"
   `include "mby_mgp_mem_crdt_io.sv"
   `include "mby_mgp_flow_ctrl.sv"
   `include "mby_mgp_agent_cfg.sv"
   `include "mby_mgp_req_agent_cfg.sv"
   `include "mby_mgp_req_seq_item.sv"
   `include "mby_mgp_rdreq_drv.sv"
   `include "mby_mgp_rdreq_mon.sv"
   `include "mby_mgp_rdreq_agent.sv"
   `include "mby_mgp_wrreq_drv.sv"
   `include "mby_mgp_wrreq_mon.sv"
   `include "mby_mgp_wrreq_agent.sv"
   `include "mby_mgp_rdrsp_drv.sv"
   `include "mby_mgp_rdrsp_mon.sv"
   `include "mby_mgp_rdrsp_agent.sv"
   `include "mby_mgp_agent.sv"
   `include "mby_mgp_bfm.sv"

endpackage