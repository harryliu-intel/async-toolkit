/*
 ******************************************************************************
 *
 *                     I N T E L   C O R P O R A T I O N
 *
 *                         Copyright(c) 2016
 *
 *                         All Rights Reserved
 *
 ******************************************************************************
 *
 * File Name   : ti_macro_defines.svh
 *
 * Author      : Mat.Khir Md Haniffa
 *
 * Last Update : 2016.w34.1
 *
 * Description : List the macros used for test island connectivity.
 *               RTL hierarchies must not be hardcoded in this file, instead
 *               should reference fc_hier_defines_generated.sv, which is a
 *               collage generated file
 *
 ******************************************************************************
*/
// Macros used to ease IOSF-SB interface connectivity
`include "iosfsb_conn_defines.svh"

`define HVL_TOP              fc_hvl_top
`define HDL_TOP              fc_hdl_top
`define DUT_IF               `HDL_TOP.fctop_dut_if
`define soc                  `HDL_TOP.dut
`define FCSIG_IF             `HVL_TOP.fc_sig_if
`define HDL_TOP_LIB          `HDL_TOP``_lib
`define HDL_TOP_CFG          `HDL_TOP``_cfg
`define HVL_TOP_LIB          `HVL_TOP``_lib
`define HVL_TOP_CFG          `HVL_TOP``_cfg
`define HDL_TOP_REALMIA_CFG  `HDL_TOP``_realmia_cfg
`define RTL_STUB_LIB         soc_ip_stub_lib
`define FCGPIO_IF `HVL_TOP.fc_gpio_if1

// All RTL hierarchy related defines are generated from Collage output
//`ifdef SOCFC
//`include "soc_ip_hier_defines.sv"
//`include "fc_hier_defines_generated.sv"
//`endif

// <<< PMC TI param
// PMC_TOP needs to be pointing to pmc_pwell because of what is
// in Declarations.svh in pmc/verif/tb/include/Declarations.svh
`define PMU_WRAPPER1 soc.pargpio.pmu_wrapper1
// >>>

// <<< RTC
// >>>

// <<< FUSE
`define FUSE_TB_ROOT         `HVL_TOP
// >>>


// <<< GPIO
`ifndef GPCOMMSTUNIT_WRAPPER
`define GPCOMMSTUNIT_WRAPPER soc.pargpio.gpcommstunit_wrapper
`endif
`define MAX_COM_NUM            1
`define GPIOCOMMST_TOP         `GPCOMMSTUNIT_WRAPPER
// >>>

// <<< DFX
// >>>

// <<< Macro to set fuse/strap values
// >>>

// <<< PARTITION
// >>>

// <<< HSUART
//define   HSUART    `HSU_UARTIOSF_TOP
//define   HSUART_TI `HVL_TOP.hsuart_ti
// >>>

// <<< PSF
`ifndef psf0
`define psf0 `soc.parmain.psf0
`endif
`ifndef psf1
`define psf1 `soc.parmain.psf1
`endif
`define PSF20_DLC_PSF0_TOP     `psf0.i_psf20_top_psf0
`define PSF20_DLC_PSF1_TOP     `psf1.i_psf20_top_psf1
// >>>

// <<< IO_WIDGET
//`define IOW_TOP                `CPK_IO_WIDGET
// >>>

// <<< ICM
//`define ICM_TOP_RTL `icm_top
// >>>

// <<< PE / RDMA
//`define PE_FUNC_LOGIC `pe_top.pe_core_apr.pe_func_logic
// >>>

// <<< SB endpoints reset & clocks
// CHS autogenerated
// GP
`define USP_SB_CLK 0
`define USP_SB_RST_B 0
`define PSF0_SB_CLK `psf0.side_clk
`define PSF0_SB_RST_B `psf0.side_rst_b
`define VSP0_SB_CLK 0
`define VSP0_SB_RST_B 0
`define VSP1_SB_CLK 0
`define VSP1_SB_RST_B 0
`define VSP2_SB_CLK 0
`define VSP2_SB_RST_B 0
`define P2SB_SB_CLK 0
`define P2SB_SB_RST_B 0
`define IEH_SB_CLK 0
`define IEH_SB_RST_B 0
`define FUSE_GP_SB_CLK `fuse_top.fuse_side_clk
`define FUSE_GP_SB_RST_B `fuse_top.fuse_side_rst_b
`define DRNG_SB_CLK `fuse_top.drng_side_clk
`define DRNG_SB_RST_B `fuse_top.drng_side_rst_b
`define DTS_GP_SB_CLK 0
`define DTS_GP_SB_RST_B 0
`define PSF1_SB_CLK `psf1.side_clk
`define PSF1_SB_RST_B `psf1.side_rst_b
`define VSP3_SB_CLK 0
`define VSP3_SB_RST_B 0
`define VSP4_SB_CLK 0
`define VSP4_SB_RST_B 0
`define CPM_SB_CLK 0
`define CPM_SB_RST_B 0
`define HQM1_GP_SB_CLK 0
`define HQM1_GP_SB_RST_B 0
`define HQM2_GP_SB_CLK 0
`define HQM2_GP_SB_RST_B 0
`define ESPI_SB_CLK 0
`define ESPI_SB_RST_B 0
`define CCU_SB_CLK `ccu_top.ccu_side_clk
`define CCU_SB_RST_B `ccu_top.ccu_side_rst_b
`define EC_SB_CLK 0
`define EC_SB_RST_B 0
`define NPK_SB_CLK `northpeak.npk_side_clk
`define NPK_SB_RST_B `northpeak.npk_side_rst_b
`define RU_GP_SB_CLK 0
`define RU_GP_SB_RST_B 0
`define MGFIA_SB_CLK 0
`define MGFIA_SB_RST_B 0
`define MGPHY_GP_SB_CLK 0
`define MGPHY_GP_SB_RST_B 0
`define DSA_SB_CLK `dfxagg_top.dfxagg_side_clock
`define DSA_SB_RST_B `dfxagg_top.dfxagg_side_rst_b
`define TAP2SB0_SB_CLK 0
`define TAP2SB0_SB_RST_B 0
`define PLL_GP_SB_CLK 0
`define PLL_GP_SB_RST_B 0
`define FIVR_GP_SB_CLK 0
`define FIVR_GP_SB_RST_B 0
`define GPIO_SB_CLK `gpcomgpiocom0unit_wrapper.side_clk
`define GPIO_SB_RST_B `gpcomgpiocom0unit_wrapper.sbi_rst_b
`define PSV_GP_SB_CLK `sbr_gp1.sbr_clk
`define PSV_GP_SB_RST_B `sbr_gp1.sbr_rst_b
// PM
`define FIVR_PM_SB_CLK 0
`define FIVR_PM_SB_RST_B 0
`define FUSE_PM_SB_CLK 0
`define FUSE_PM_SB_RST_B 0
`define DTS_PM_SB_CLK 0
`define DTS_PM_SB_RST_B 0
`define MGPHY_PM_SB_CLK 0
`define MGPHY_PM_SB_RST_B 0
`define PSV_PM_SB_CLK 0
`define PSV_PM_SB_RST_B 0
`define PLL_PM_SB_CLK 0
`define PLL_PM_SB_RST_B 0
`define RU_PM_SB_CLK 0
`define RU_PM_SB_RST_B 0
`define TAP2SB1_SB_CLK 0
`define TAP2SB1_SB_RST_B 0
`define HQM1_PM_SB_CLK 0
`define HQM1_PM_SB_RST_B 0
`define HQM2_PM_SB_CLK 0
`define HQM2_PM_SB_RST_B 0
// >>>

// <<< NORTHPEAK
`ifndef northpeak
`define northpeak      `soc.parmain.northpeak
`endif
`define NORTHPEAK_INST_NAME     `northpeak
`define NPK_TTC_INST_NAME       `northpeak.i_npk_vnn_gated_wrapper.i_npk_ttc
`define NPK_TPH_INST_NAME       `northpeak.i_npk_vnn_gated_wrapper.i_npk_tph
// >>>


/*
 *  ----------------
 *    End of file
 *  ----------------
*/
// <<< VIM SETTINGS
// vim: ts=4 et
// >>>
