///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///
// -------------------------------------------------------------------
// -- Intel Proprietary
// -- Copyright (C) 2018 Intel Corporation
// -- All Rights Reserved
// -------------------------------------------------------------------
// -- Author : Jon Bagge <jon.bagge@intel.com>
// -- Project Name : Madison Bay
// -- Description : Egress to shared table memory interface
// --
// -------------------------------------------------------------------

interface egr_ppe_stm_if
();
logic           [7:0]   wen;    //per chunk write enables
logic   [1:0]   [7:0]   ren;    //per port, per chunk read enables
logic   [2:0]   [17:0]  addr;   //per port address (port 0 is write, 1-2 are read)
logic           [575:0] wdata;  //write data (including ECC bits)
logic   [1:0]   [575:0] rdata;  //read data (including ECC bits)

modport egr(
    output  wen,
    output  ren,
    output  addr,
    output  wdata,
    input   rdata
);

modport stm(
    input   wen,
    input   ren,
    input   addr,
    input   wdata,
    output  rdata
);

endinterface: egr_ppe_stm_if
