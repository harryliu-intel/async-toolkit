rtlgen_include_v12.vh