magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect 25 -3 35 -2
rect 25 -6 35 -5
rect 25 -10 27 -6
rect 25 -11 35 -10
rect 25 -14 35 -13
rect 29 -18 35 -14
rect 25 -19 35 -18
rect 25 -22 35 -21
rect 25 -26 27 -22
rect 25 -27 35 -26
rect 25 -30 35 -29
rect 29 -34 35 -30
rect 25 -35 35 -34
rect 25 -38 35 -37
rect 25 -42 27 -38
rect 25 -43 35 -42
rect 25 -46 35 -45
<< pdiffusion >>
rect 47 -7 53 -6
rect 47 -13 53 -9
rect 47 -19 53 -15
rect 47 -22 53 -21
rect 51 -26 53 -22
rect 47 -27 53 -26
rect 47 -33 53 -29
rect 47 -39 53 -35
rect 47 -42 53 -41
<< ntransistor >>
rect 25 -5 35 -3
rect 25 -13 35 -11
rect 25 -21 35 -19
rect 25 -29 35 -27
rect 25 -37 35 -35
rect 25 -45 35 -43
<< ptransistor >>
rect 47 -9 53 -7
rect 47 -15 53 -13
rect 47 -21 53 -19
rect 47 -29 53 -27
rect 47 -35 53 -33
rect 47 -41 53 -39
<< polysilicon >>
rect 22 -5 25 -3
rect 35 -5 45 -3
rect 43 -7 45 -5
rect 43 -9 47 -7
rect 53 -9 56 -7
rect 22 -13 25 -11
rect 35 -13 39 -11
rect 37 -15 47 -13
rect 53 -15 56 -13
rect 22 -21 25 -19
rect 35 -21 47 -19
rect 53 -21 56 -19
rect 22 -29 25 -27
rect 35 -29 47 -27
rect 53 -29 56 -27
rect 37 -35 47 -33
rect 53 -35 56 -33
rect 22 -37 25 -35
rect 35 -37 39 -35
rect 43 -41 47 -39
rect 53 -41 56 -39
rect 43 -43 45 -41
rect 22 -45 25 -43
rect 35 -45 45 -43
<< ndcontact >>
rect 25 -2 35 2
rect 27 -10 35 -6
rect 25 -18 29 -14
rect 27 -26 35 -22
rect 25 -34 29 -30
rect 27 -42 35 -38
rect 25 -50 35 -46
<< pdcontact >>
rect 47 -6 53 -2
rect 47 -26 51 -22
rect 47 -46 53 -42
<< metal1 >>
rect 25 -2 35 2
rect 47 -6 53 -2
rect 27 -10 35 -6
rect 25 -18 29 -14
rect 32 -22 35 -10
rect 27 -26 51 -22
rect 25 -34 29 -30
rect 32 -38 35 -26
rect 27 -42 35 -38
rect 47 -46 53 -42
rect 25 -50 35 -46
<< labels >>
rlabel space 21 -51 28 3 7 ^n
rlabel space 50 -47 56 -1 3 ^p
rlabel polysilicon 54 -28 54 -28 7 c
rlabel polysilicon 54 -34 54 -34 7 b
rlabel polysilicon 54 -40 54 -40 7 a
rlabel polysilicon 54 -20 54 -20 7 a
rlabel polysilicon 54 -14 54 -14 7 b
rlabel polysilicon 24 -44 24 -44 7 a
rlabel polysilicon 24 -20 24 -20 7 a
rlabel polysilicon 24 -36 24 -36 7 b
rlabel polysilicon 24 -12 24 -12 7 b
rlabel polysilicon 24 -28 24 -28 7 c
rlabel polysilicon 24 -4 24 -4 7 c
rlabel polysilicon 54 -8 54 -8 7 c
rlabel ndcontact 33 -8 33 -8 1 x
rlabel ndcontact 33 -24 33 -24 1 x
rlabel ndcontact 33 -40 33 -40 1 x
rlabel pdcontact 49 -24 49 -24 1 x
rlabel pdcontact 49 -44 49 -44 1 Vdd!
rlabel pdcontact 49 -4 49 -4 1 Vdd!
rlabel ndcontact 27 -16 27 -16 1 GND!
rlabel ndcontact 27 0 27 0 5 GND!
rlabel ndcontact 27 -32 27 -32 1 GND!
rlabel ndcontact 27 -48 27 -48 1 GND!
<< end >>
