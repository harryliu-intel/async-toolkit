magic
tech scmos
timestamp 970030488
<< ndiffusion >>
rect -24 49 -8 50
rect -24 41 -8 46
rect -24 33 -8 38
rect -24 25 -8 30
rect -24 21 -8 22
rect -24 12 -8 13
<< pdiffusion >>
rect 8 54 34 55
rect 8 50 34 51
rect 22 42 34 50
rect 8 41 34 42
rect 8 37 34 38
rect 8 28 34 29
rect 8 24 34 25
rect 8 13 24 16
rect 8 9 24 10
<< ntransistor >>
rect -24 46 -8 49
rect -24 38 -8 41
rect -24 30 -8 33
rect -24 22 -8 25
<< ptransistor >>
rect 8 51 34 54
rect 8 38 34 41
rect 8 25 34 28
rect 8 10 24 13
<< polysilicon >>
rect 3 51 8 54
rect 34 51 38 54
rect 3 49 6 51
rect -28 46 -24 49
rect -8 46 6 49
rect -28 38 -24 41
rect -8 38 8 41
rect 34 38 38 41
rect -28 30 -24 33
rect -8 30 6 33
rect 3 28 6 30
rect 3 25 8 28
rect 34 25 38 28
rect -28 22 -24 25
rect -8 22 -4 25
rect 4 10 8 13
rect 24 10 31 13
rect 28 9 31 10
<< ndcontact >>
rect -24 50 -8 58
rect -24 13 -8 21
<< pdcontact >>
rect 8 55 34 63
rect 8 42 22 50
rect 8 29 34 37
rect 8 16 34 24
rect 8 1 24 9
<< psubstratepcontact >>
rect -24 4 -8 12
<< nsubstratencontact >>
rect 43 51 51 59
<< polycontact >>
rect -36 46 -28 54
rect 38 38 46 46
rect 38 25 46 33
rect -36 17 -28 25
rect 28 1 36 9
<< metal1 >>
rect 21 61 34 63
rect 8 59 34 61
rect -24 50 -8 58
rect 8 55 51 59
rect 26 51 51 55
rect -36 46 -28 49
rect -16 42 22 50
rect -36 7 -28 25
rect -4 24 4 42
rect 26 37 34 51
rect 38 43 46 46
rect 8 29 34 37
rect 38 31 46 33
rect -24 7 -8 21
rect -4 19 34 24
rect 4 16 34 19
rect 8 7 24 9
rect -24 4 -21 7
rect 21 1 24 7
rect 28 7 36 9
<< m2contact >>
rect 3 61 21 67
rect -36 49 -28 55
rect 38 37 46 43
rect 38 25 46 31
rect -36 1 -28 7
rect -4 13 4 19
rect -21 1 -3 7
rect 3 1 21 7
rect 28 1 36 7
<< metal2 >>
rect -36 49 0 55
rect 0 37 46 43
rect 0 25 46 31
rect -6 13 6 19
rect -37 1 -26 7
rect 26 1 37 7
<< m3contact >>
rect 3 61 21 67
rect -21 1 -3 7
rect 3 1 21 7
<< metal3 >>
rect -21 -2 -3 70
rect 3 -2 21 70
<< labels >>
rlabel m2contact 12 5 12 5 1 Vdd!
rlabel metal1 12 20 12 20 1 x
rlabel metal1 12 59 12 59 5 Vdd!
rlabel metal1 12 33 12 33 1 Vdd!
rlabel metal1 12 46 12 46 5 x
rlabel metal1 -12 17 -12 17 1 GND!
rlabel metal1 -12 54 -12 54 1 x
rlabel polysilicon -25 47 -25 47 3 c
rlabel polysilicon -25 39 -25 39 3 b
rlabel polysilicon -25 31 -25 31 3 a
rlabel polysilicon -25 23 -25 23 3 _SReset!
rlabel polysilicon 35 52 35 52 1 c
rlabel polysilicon 35 26 35 26 1 a
rlabel polysilicon 35 39 35 39 1 b
rlabel polysilicon 25 12 25 12 5 _PReset!
rlabel metal2 32 4 32 4 1 _PReset!
rlabel metal2 -32 4 -32 4 3 _SReset!
rlabel metal2 0 16 0 16 1 x
rlabel metal2 0 25 0 31 3 a
rlabel metal2 0 49 0 55 7 c
rlabel space -38 0 -24 59 7 ^n
rlabel metal2 -26 1 -26 7 3 ^n
rlabel metal1 47 55 47 55 7 Vdd!
rlabel space 22 20 52 64 3 ^p
rlabel metal2 -32 52 -32 52 1 c
rlabel metal2 42 40 42 40 1 b
rlabel metal2 42 28 42 28 1 a
rlabel metal2 0 37 0 43 3 b
<< end >>
