///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_fwd_misc_map_pkg.vh                                
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template

`ifndef MBY_PPE_FWD_MISC_MAP_PKG_VH
`define MBY_PPE_FWD_MISC_MAP_PKG_VH

`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"

package mby_ppe_fwd_misc_map_pkg;

import rtlgen_pkg_mby_top_map::*;

typedef cfg_req_64bit_t mby_ppe_fwd_misc_map_cr_req_t;
typedef cfg_ack_64bit_t mby_ppe_fwd_misc_map_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} mby_ppe_fwd_misc_map_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [39:0] reserved0;  // RSVD
    logic [23:0] DESTINATION_MASK;  // RW
} FWD_PORT_CFG_2_t;

localparam FWD_PORT_CFG_2_REG_STRIDE = 48'h8;
localparam FWD_PORT_CFG_2_REG_ENTRIES = 256;
localparam FWD_PORT_CFG_2_CR_ADDR = 48'h0;
localparam FWD_PORT_CFG_2_SIZE = 64;
localparam FWD_PORT_CFG_2_DESTINATION_MASK_LO = 0;
localparam FWD_PORT_CFG_2_DESTINATION_MASK_HI = 23;
localparam FWD_PORT_CFG_2_DESTINATION_MASK_RESET = 24'hffffff;
localparam FWD_PORT_CFG_2_USEMASK = 64'hFFFFFF;
localparam FWD_PORT_CFG_2_RO_MASK = 64'h0;
localparam FWD_PORT_CFG_2_WO_MASK = 64'h0;
localparam FWD_PORT_CFG_2_RESET = 64'hFFFFFF;

typedef struct packed {
    logic [53:0] reserved0;  // RSVD
    logic  [0:0] IN_LAG;  // RW
    logic  [0:0] HASH_ROTATION;  // RW
    logic  [3:0] INDEX;  // RW
    logic  [3:0] LAG_SIZE;  // RW
} FWD_LAG_CFG_t;

localparam FWD_LAG_CFG_REG_STRIDE = 48'h8;
localparam FWD_LAG_CFG_REG_ENTRIES = 17;
localparam FWD_LAG_CFG_CR_ADDR = 48'h1000;
localparam FWD_LAG_CFG_SIZE = 64;
localparam FWD_LAG_CFG_IN_LAG_LO = 9;
localparam FWD_LAG_CFG_IN_LAG_HI = 9;
localparam FWD_LAG_CFG_IN_LAG_RESET = 1'h0;
localparam FWD_LAG_CFG_HASH_ROTATION_LO = 8;
localparam FWD_LAG_CFG_HASH_ROTATION_HI = 8;
localparam FWD_LAG_CFG_HASH_ROTATION_RESET = 1'h0;
localparam FWD_LAG_CFG_INDEX_LO = 4;
localparam FWD_LAG_CFG_INDEX_HI = 7;
localparam FWD_LAG_CFG_INDEX_RESET = 4'h0;
localparam FWD_LAG_CFG_LAG_SIZE_LO = 0;
localparam FWD_LAG_CFG_LAG_SIZE_HI = 3;
localparam FWD_LAG_CFG_LAG_SIZE_RESET = 4'h0;
localparam FWD_LAG_CFG_USEMASK = 64'h3FF;
localparam FWD_LAG_CFG_RO_MASK = 64'h0;
localparam FWD_LAG_CFG_WO_MASK = 64'h0;
localparam FWD_LAG_CFG_RESET = 64'h0;

typedef struct packed {
    logic [37:0] reserved0;  // RSVD
    logic  [0:0] LEARNING_ENABLE;  // RW
    logic  [0:0] FILTER_VLAN_INGRESS;  // RW
    logic [23:0] DESTINATION_MASK;  // RW
} FWD_PORT_CFG_1_t;

localparam FWD_PORT_CFG_1_REG_STRIDE = 48'h8;
localparam FWD_PORT_CFG_1_REG_ENTRIES = 17;
localparam FWD_PORT_CFG_1_CR_ADDR = 48'h1100;
localparam FWD_PORT_CFG_1_SIZE = 64;
localparam FWD_PORT_CFG_1_LEARNING_ENABLE_LO = 25;
localparam FWD_PORT_CFG_1_LEARNING_ENABLE_HI = 25;
localparam FWD_PORT_CFG_1_LEARNING_ENABLE_RESET = 1'h1;
localparam FWD_PORT_CFG_1_FILTER_VLAN_INGRESS_LO = 24;
localparam FWD_PORT_CFG_1_FILTER_VLAN_INGRESS_HI = 24;
localparam FWD_PORT_CFG_1_FILTER_VLAN_INGRESS_RESET = 1'h1;
localparam FWD_PORT_CFG_1_DESTINATION_MASK_LO = 0;
localparam FWD_PORT_CFG_1_DESTINATION_MASK_HI = 23;
localparam FWD_PORT_CFG_1_DESTINATION_MASK_RESET = 24'hffffff;
localparam FWD_PORT_CFG_1_USEMASK = 64'h3FFFFFF;
localparam FWD_PORT_CFG_1_RO_MASK = 64'h0;
localparam FWD_PORT_CFG_1_WO_MASK = 64'h0;
localparam FWD_PORT_CFG_1_RESET = 64'h3FFFFFF;

typedef struct packed {
    logic [58:0] reserved0;  // RSVD
    logic  [0:0] STORE_TRAP_ACTION;  // RW
    logic  [0:0] DROP_MAC_CTRL_ETHERTYPE;  // RW
    logic  [0:0] DROP_INVALID_SMAC;  // RW
    logic  [0:0] ENABLE_TRAP_PLUS_LOG;  // RW
    logic  [0:0] TRAP_MTU_VIOLATIONS;  // RW
} FWD_SYS_CFG_1_t;

localparam FWD_SYS_CFG_1_REG_STRIDE = 48'h8;
localparam FWD_SYS_CFG_1_REG_ENTRIES = 1;
localparam [47:0] FWD_SYS_CFG_1_CR_ADDR = 48'h1200;
localparam FWD_SYS_CFG_1_SIZE = 64;
localparam FWD_SYS_CFG_1_STORE_TRAP_ACTION_LO = 4;
localparam FWD_SYS_CFG_1_STORE_TRAP_ACTION_HI = 4;
localparam FWD_SYS_CFG_1_STORE_TRAP_ACTION_RESET = 1'h1;
localparam FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE_LO = 3;
localparam FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE_HI = 3;
localparam FWD_SYS_CFG_1_DROP_MAC_CTRL_ETHERTYPE_RESET = 1'h1;
localparam FWD_SYS_CFG_1_DROP_INVALID_SMAC_LO = 2;
localparam FWD_SYS_CFG_1_DROP_INVALID_SMAC_HI = 2;
localparam FWD_SYS_CFG_1_DROP_INVALID_SMAC_RESET = 1'h1;
localparam FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG_LO = 1;
localparam FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG_HI = 1;
localparam FWD_SYS_CFG_1_ENABLE_TRAP_PLUS_LOG_RESET = 1'h1;
localparam FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS_LO = 0;
localparam FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS_HI = 0;
localparam FWD_SYS_CFG_1_TRAP_MTU_VIOLATIONS_RESET = 1'h1;
localparam FWD_SYS_CFG_1_USEMASK = 64'h1F;
localparam FWD_SYS_CFG_1_RO_MASK = 64'h0;
localparam FWD_SYS_CFG_1_WO_MASK = 64'h0;
localparam FWD_SYS_CFG_1_RESET = 64'h1F;

typedef struct packed {
    logic [15:0] reserved0;  // RSVD
    logic [47:0] MAC_ADDR;  // RW
} FWD_CPU_MAC_t;

localparam FWD_CPU_MAC_REG_STRIDE = 48'h8;
localparam FWD_CPU_MAC_REG_ENTRIES = 1;
localparam [47:0] FWD_CPU_MAC_CR_ADDR = 48'h1208;
localparam FWD_CPU_MAC_SIZE = 64;
localparam FWD_CPU_MAC_MAC_ADDR_LO = 0;
localparam FWD_CPU_MAC_MAC_ADDR_HI = 47;
localparam FWD_CPU_MAC_MAC_ADDR_RESET = 48'h0;
localparam FWD_CPU_MAC_USEMASK = 64'hFFFFFFFFFFFF;
localparam FWD_CPU_MAC_RO_MASK = 64'h0;
localparam FWD_CPU_MAC_WO_MASK = 64'h0;
localparam FWD_CPU_MAC_RESET = 64'h0;

typedef struct packed {
    logic [60:0] reserved0;  // RSVD
    logic  [0:0] TRAP_IP_OPTIONS;  // RW
    logic  [1:0] TRAP_TTL1;  // RW
} FWD_SYS_CFG_ROUTER_t;

localparam FWD_SYS_CFG_ROUTER_REG_STRIDE = 48'h8;
localparam FWD_SYS_CFG_ROUTER_REG_ENTRIES = 1;
localparam [47:0] FWD_SYS_CFG_ROUTER_CR_ADDR = 48'h1210;
localparam FWD_SYS_CFG_ROUTER_SIZE = 64;
localparam FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS_LO = 2;
localparam FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS_HI = 2;
localparam FWD_SYS_CFG_ROUTER_TRAP_IP_OPTIONS_RESET = 1'h0;
localparam FWD_SYS_CFG_ROUTER_TRAP_TTL1_LO = 0;
localparam FWD_SYS_CFG_ROUTER_TRAP_TTL1_HI = 1;
localparam FWD_SYS_CFG_ROUTER_TRAP_TTL1_RESET = 2'h0;
localparam FWD_SYS_CFG_ROUTER_USEMASK = 64'h7;
localparam FWD_SYS_CFG_ROUTER_RO_MASK = 64'h0;
localparam FWD_SYS_CFG_ROUTER_WO_MASK = 64'h0;
localparam FWD_SYS_CFG_ROUTER_RESET = 64'h0;

typedef struct packed {
    logic [57:0] reserved0;  // RSVD
    logic  [5:0] MIRROR_PROFILE_IDX;  // RW
} FWD_RX_MIRROR_CFG_t;

localparam FWD_RX_MIRROR_CFG_REG_STRIDE = 48'h8;
localparam FWD_RX_MIRROR_CFG_REG_ENTRIES = 1;
localparam [47:0] FWD_RX_MIRROR_CFG_CR_ADDR = 48'h1218;
localparam FWD_RX_MIRROR_CFG_SIZE = 64;
localparam FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX_LO = 0;
localparam FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX_HI = 5;
localparam FWD_RX_MIRROR_CFG_MIRROR_PROFILE_IDX_RESET = 6'h0;
localparam FWD_RX_MIRROR_CFG_USEMASK = 64'h3F;
localparam FWD_RX_MIRROR_CFG_RO_MASK = 64'h0;
localparam FWD_RX_MIRROR_CFG_WO_MASK = 64'h0;
localparam FWD_RX_MIRROR_CFG_RESET = 64'h0;

typedef struct packed {
    logic [55:0] reserved0;  // RSVD
    logic  [5:0] MIRROR_PROFILE_IDX;  // RW
    logic  [1:0] MIRROR_SESSION;  // RW
} FWD_QCN_MIRROR_CFG_t;

localparam FWD_QCN_MIRROR_CFG_REG_STRIDE = 48'h8;
localparam FWD_QCN_MIRROR_CFG_REG_ENTRIES = 1;
localparam [47:0] FWD_QCN_MIRROR_CFG_CR_ADDR = 48'h1220;
localparam FWD_QCN_MIRROR_CFG_SIZE = 64;
localparam FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX_LO = 2;
localparam FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX_HI = 7;
localparam FWD_QCN_MIRROR_CFG_MIRROR_PROFILE_IDX_RESET = 6'h0;
localparam FWD_QCN_MIRROR_CFG_MIRROR_SESSION_LO = 0;
localparam FWD_QCN_MIRROR_CFG_MIRROR_SESSION_HI = 1;
localparam FWD_QCN_MIRROR_CFG_MIRROR_SESSION_RESET = 2'h0;
localparam FWD_QCN_MIRROR_CFG_USEMASK = 64'hFF;
localparam FWD_QCN_MIRROR_CFG_RO_MASK = 64'h0;
localparam FWD_QCN_MIRROR_CFG_WO_MASK = 64'h0;
localparam FWD_QCN_MIRROR_CFG_RESET = 64'h0;

typedef struct packed {
    logic  [1:0] ACTION_63;  // RW
    logic  [1:0] ACTION_62;  // RW
    logic  [1:0] ACTION_61;  // RW
    logic  [1:0] ACTION_60;  // RW
    logic  [1:0] ACTION_59;  // RW
    logic  [1:0] ACTION_58;  // RW
    logic  [1:0] ACTION_57;  // RW
    logic  [1:0] ACTION_56;  // RW
    logic  [1:0] ACTION_55;  // RW
    logic  [1:0] ACTION_54;  // RW
    logic  [1:0] ACTION_53;  // RW
    logic  [1:0] ACTION_52;  // RW
    logic  [1:0] ACTION_51;  // RW
    logic  [1:0] ACTION_50;  // RW
    logic  [1:0] ACTION_49;  // RW
    logic  [1:0] ACTION_48;  // RW
    logic  [1:0] ACTION_47;  // RW
    logic  [1:0] ACTION_46;  // RW
    logic  [1:0] ACTION_45;  // RW
    logic  [1:0] ACTION_44;  // RW
    logic  [1:0] ACTION_43;  // RW
    logic  [1:0] ACTION_42;  // RW
    logic  [1:0] ACTION_41;  // RW
    logic  [1:0] ACTION_40;  // RW
    logic  [1:0] ACTION_39;  // RW
    logic  [1:0] ACTION_38;  // RW
    logic  [1:0] ACTION_37;  // RW
    logic  [1:0] ACTION_36;  // RW
    logic  [1:0] ACTION_35;  // RW
    logic  [1:0] ACTION_34;  // RW
    logic  [1:0] ACTION_33;  // RW
    logic  [1:0] ACTION_32;  // RW
    logic  [1:0] ACTION_31;  // RW
    logic  [1:0] ACTION_30;  // RW
    logic  [1:0] ACTION_29;  // RW
    logic  [1:0] ACTION_28;  // RW
    logic  [1:0] ACTION_27;  // RW
    logic  [1:0] ACTION_26;  // RW
    logic  [1:0] ACTION_25;  // RW
    logic  [1:0] ACTION_24;  // RW
    logic  [1:0] ACTION_23;  // RW
    logic  [1:0] ACTION_22;  // RW
    logic  [1:0] ACTION_21;  // RW
    logic  [1:0] ACTION_20;  // RW
    logic  [1:0] ACTION_19;  // RW
    logic  [1:0] ACTION_18;  // RW
    logic  [1:0] ACTION_17;  // RW
    logic  [1:0] ACTION_16;  // RW
    logic  [1:0] ACTION_15;  // RW
    logic  [1:0] ACTION_14;  // RW
    logic  [1:0] ACTION_13;  // RW
    logic  [1:0] ACTION_12;  // RW
    logic  [1:0] ACTION_11;  // RW
    logic  [1:0] ACTION_10;  // RW
    logic  [1:0] ACTION_9;  // RW
    logic  [1:0] ACTION_8;  // RW
    logic  [1:0] ACTION_7;  // RW
    logic  [1:0] ACTION_6;  // RW
    logic  [1:0] ACTION_5;  // RW
    logic  [1:0] ACTION_4;  // RW
    logic  [1:0] ACTION_3;  // RW
    logic  [1:0] ACTION_2;  // RW
    logic  [1:0] ACTION_1;  // RW
    logic  [1:0] ACTION_0;  // RW
} FWD_IEEE_RESERVED_MAC_ACTION_t;

localparam FWD_IEEE_RESERVED_MAC_ACTION_REG_STRIDE = 48'h10;
localparam FWD_IEEE_RESERVED_MAC_ACTION_REG_ENTRIES = 1;
localparam [47:0] FWD_IEEE_RESERVED_MAC_ACTION_CR_ADDR = 48'h1230;
localparam FWD_IEEE_RESERVED_MAC_ACTION_SIZE = 128;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63_LO = 126;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63_HI = 127;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_63_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62_LO = 124;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62_HI = 125;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_62_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61_LO = 122;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61_HI = 123;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_61_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60_LO = 120;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60_HI = 121;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_60_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59_LO = 118;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59_HI = 119;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_59_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58_LO = 116;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58_HI = 117;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_58_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57_LO = 114;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57_HI = 115;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_57_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56_LO = 112;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56_HI = 113;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_56_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55_LO = 110;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55_HI = 111;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_55_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54_LO = 108;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54_HI = 109;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_54_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53_LO = 106;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53_HI = 107;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_53_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52_LO = 104;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52_HI = 105;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_52_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51_LO = 102;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51_HI = 103;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_51_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50_LO = 100;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50_HI = 101;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_50_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49_LO = 98;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49_HI = 99;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_49_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48_LO = 96;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48_HI = 97;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_48_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47_LO = 94;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47_HI = 95;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_47_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46_LO = 92;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46_HI = 93;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_46_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45_LO = 90;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45_HI = 91;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_45_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44_LO = 88;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44_HI = 89;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_44_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43_LO = 86;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43_HI = 87;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_43_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42_LO = 84;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42_HI = 85;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_42_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41_LO = 82;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41_HI = 83;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_41_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40_LO = 80;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40_HI = 81;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_40_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39_LO = 78;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39_HI = 79;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_39_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38_LO = 76;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38_HI = 77;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_38_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37_LO = 74;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37_HI = 75;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_37_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36_LO = 72;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36_HI = 73;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_36_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35_LO = 70;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35_HI = 71;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_35_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34_LO = 68;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34_HI = 69;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_34_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33_LO = 66;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33_HI = 67;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_33_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32_LO = 64;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32_HI = 65;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_32_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31_LO = 62;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31_HI = 63;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_31_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30_LO = 60;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30_HI = 61;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_30_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29_LO = 58;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29_HI = 59;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_29_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28_LO = 56;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28_HI = 57;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_28_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27_LO = 54;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27_HI = 55;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_27_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26_LO = 52;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26_HI = 53;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_26_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25_LO = 50;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25_HI = 51;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_25_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24_LO = 48;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24_HI = 49;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_24_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23_LO = 46;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23_HI = 47;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_23_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22_LO = 44;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22_HI = 45;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_22_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21_LO = 42;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21_HI = 43;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_21_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20_LO = 40;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20_HI = 41;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_20_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19_LO = 38;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19_HI = 39;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_19_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18_LO = 36;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18_HI = 37;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_18_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17_LO = 34;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17_HI = 35;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_17_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16_LO = 32;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16_HI = 33;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_16_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15_LO = 30;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15_HI = 31;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_15_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14_LO = 28;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14_HI = 29;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_14_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13_LO = 26;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13_HI = 27;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_13_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12_LO = 24;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12_HI = 25;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_12_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11_LO = 22;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11_HI = 23;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_11_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10_LO = 20;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10_HI = 21;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_10_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9_LO = 18;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9_HI = 19;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_9_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8_LO = 16;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8_HI = 17;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_8_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7_LO = 14;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7_HI = 15;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_7_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6_LO = 12;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6_HI = 13;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_6_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5_LO = 10;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5_HI = 11;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_5_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4_LO = 8;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4_HI = 9;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_4_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3_LO = 6;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3_HI = 7;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_3_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2_LO = 4;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2_HI = 5;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_2_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1_LO = 2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1_HI = 3;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_1_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0_LO = 0;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0_HI = 1;
localparam FWD_IEEE_RESERVED_MAC_ACTION_ACTION_0_RESET = 2'h2;
localparam FWD_IEEE_RESERVED_MAC_ACTION_USEMASK = 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
localparam FWD_IEEE_RESERVED_MAC_ACTION_RO_MASK = 128'h0;
localparam FWD_IEEE_RESERVED_MAC_ACTION_WO_MASK = 128'h0;
localparam FWD_IEEE_RESERVED_MAC_ACTION_RESET = 128'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;

typedef struct packed {
    logic [63:0] SELECT;  // RW
} FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_t;

localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_REG_STRIDE = 48'h8;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_REG_ENTRIES = 1;
localparam [47:0] FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_CR_ADDR = 48'h1340;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SIZE = 64;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT_LO = 0;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT_HI = 63;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_SELECT_RESET = 64'h0;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_RO_MASK = 64'h0;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_WO_MASK = 64'h0;
localparam FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_RESET = 64'h0;

typedef struct packed {
    logic [60:0] reserved0;  // RSVD
    logic  [2:0] TRAP_TC;  // RW
} FWD_IEEE_RESERVED_MAC_CFG_t;

localparam FWD_IEEE_RESERVED_MAC_CFG_REG_STRIDE = 48'h8;
localparam FWD_IEEE_RESERVED_MAC_CFG_REG_ENTRIES = 1;
localparam [47:0] FWD_IEEE_RESERVED_MAC_CFG_CR_ADDR = 48'h1350;
localparam FWD_IEEE_RESERVED_MAC_CFG_SIZE = 64;
localparam FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC_LO = 0;
localparam FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC_HI = 2;
localparam FWD_IEEE_RESERVED_MAC_CFG_TRAP_TC_RESET = 3'h0;
localparam FWD_IEEE_RESERVED_MAC_CFG_USEMASK = 64'h7;
localparam FWD_IEEE_RESERVED_MAC_CFG_RO_MASK = 64'h0;
localparam FWD_IEEE_RESERVED_MAC_CFG_WO_MASK = 64'h0;
localparam FWD_IEEE_RESERVED_MAC_CFG_RESET = 64'h0;

typedef struct packed {
    logic [57:0] reserved0;  // RSVD
    logic  [0:0] MA_TCN;  // RO/V
    logic  [0:0] WB_FIFO_PERR;  // RW/1C/V
    logic  [0:0] TRIGGER;  // RO/V
    logic  [0:0] TCAM_ERR;  // RO/V
    logic  [0:0] ENTRY_COUNT;  // RO/V
    logic  [0:0] SHELL_CTRL_U_ERR;  // RW/1C/V
} FWD_IP_t;

localparam FWD_IP_REG_STRIDE = 48'h8;
localparam FWD_IP_REG_ENTRIES = 1;
localparam [47:0] FWD_IP_CR_ADDR = 48'h1360;
localparam FWD_IP_SIZE = 64;
localparam FWD_IP_MA_TCN_LO = 5;
localparam FWD_IP_MA_TCN_HI = 5;
localparam FWD_IP_MA_TCN_RESET = 1'h0;
localparam FWD_IP_WB_FIFO_PERR_LO = 4;
localparam FWD_IP_WB_FIFO_PERR_HI = 4;
localparam FWD_IP_WB_FIFO_PERR_RESET = 1'h0;
localparam FWD_IP_TRIGGER_LO = 3;
localparam FWD_IP_TRIGGER_HI = 3;
localparam FWD_IP_TRIGGER_RESET = 1'h0;
localparam FWD_IP_TCAM_ERR_LO = 2;
localparam FWD_IP_TCAM_ERR_HI = 2;
localparam FWD_IP_TCAM_ERR_RESET = 1'h0;
localparam FWD_IP_ENTRY_COUNT_LO = 1;
localparam FWD_IP_ENTRY_COUNT_HI = 1;
localparam FWD_IP_ENTRY_COUNT_RESET = 1'h0;
localparam FWD_IP_SHELL_CTRL_U_ERR_LO = 0;
localparam FWD_IP_SHELL_CTRL_U_ERR_HI = 0;
localparam FWD_IP_SHELL_CTRL_U_ERR_RESET = 1'h0;
localparam FWD_IP_USEMASK = 64'h3F;
localparam FWD_IP_RO_MASK = 64'h2E;
localparam FWD_IP_WO_MASK = 64'h0;
localparam FWD_IP_RESET = 64'h0;

typedef struct packed {
    logic [57:0] reserved0;  // RSVD
    logic  [0:0] MA_TCN;  // RO/V
    logic  [0:0] WB_FIFO_PERR;  // RW
    logic  [0:0] TRIGGER;  // RW
    logic  [0:0] TCAM_ERR;  // RW
    logic  [0:0] ENTRY_COUNT;  // RW
    logic  [0:0] SHELL_CTRL_U_ERR;  // RW
} FWD_IM_t;

localparam FWD_IM_REG_STRIDE = 48'h8;
localparam FWD_IM_REG_ENTRIES = 1;
localparam [47:0] FWD_IM_CR_ADDR = 48'h1370;
localparam FWD_IM_SIZE = 64;
localparam FWD_IM_MA_TCN_LO = 5;
localparam FWD_IM_MA_TCN_HI = 5;
localparam FWD_IM_MA_TCN_RESET = 1'h0;
localparam FWD_IM_WB_FIFO_PERR_LO = 4;
localparam FWD_IM_WB_FIFO_PERR_HI = 4;
localparam FWD_IM_WB_FIFO_PERR_RESET = 1'h1;
localparam FWD_IM_TRIGGER_LO = 3;
localparam FWD_IM_TRIGGER_HI = 3;
localparam FWD_IM_TRIGGER_RESET = 1'h1;
localparam FWD_IM_TCAM_ERR_LO = 2;
localparam FWD_IM_TCAM_ERR_HI = 2;
localparam FWD_IM_TCAM_ERR_RESET = 1'h1;
localparam FWD_IM_ENTRY_COUNT_LO = 1;
localparam FWD_IM_ENTRY_COUNT_HI = 1;
localparam FWD_IM_ENTRY_COUNT_RESET = 1'h1;
localparam FWD_IM_SHELL_CTRL_U_ERR_LO = 0;
localparam FWD_IM_SHELL_CTRL_U_ERR_HI = 0;
localparam FWD_IM_SHELL_CTRL_U_ERR_RESET = 1'h1;
localparam FWD_IM_USEMASK = 64'h3F;
localparam FWD_IM_RO_MASK = 64'h20;
localparam FWD_IM_WO_MASK = 64'h0;
localparam FWD_IM_RESET = 64'h1F;

typedef struct packed {
    FWD_SYS_CFG_1_t  FWD_SYS_CFG_1;
    FWD_CPU_MAC_t  FWD_CPU_MAC;
    FWD_SYS_CFG_ROUTER_t  FWD_SYS_CFG_ROUTER;
    FWD_RX_MIRROR_CFG_t  FWD_RX_MIRROR_CFG;
    FWD_QCN_MIRROR_CFG_t  FWD_QCN_MIRROR_CFG;
    FWD_IEEE_RESERVED_MAC_ACTION_t  FWD_IEEE_RESERVED_MAC_ACTION;
    FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY_t  FWD_IEEE_RESERVED_MAC_TRAP_PRIORITY;
    FWD_IEEE_RESERVED_MAC_CFG_t  FWD_IEEE_RESERVED_MAC_CFG;
    FWD_IP_t  FWD_IP;
    FWD_IM_t  FWD_IM;
} mby_ppe_fwd_misc_map_registers_t;

// ===================================================
// load

typedef struct packed {
    logic  [0:0] WB_FIFO_PERR;  // RW/1C/V
    logic  [0:0] SHELL_CTRL_U_ERR;  // RW/1C/V
} load_FWD_IP_t;

typedef struct packed {
    load_FWD_IP_t  FWD_IP;
} mby_ppe_fwd_misc_map_load_t;

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

typedef struct packed {
    logic  [0:0] MA_TCN;  // RO/V
    logic  [0:0] WB_FIFO_PERR;  // RW/1C/V
    logic  [0:0] TRIGGER;  // RO/V
    logic  [0:0] TCAM_ERR;  // RO/V
    logic  [0:0] ENTRY_COUNT;  // RO/V
    logic  [0:0] SHELL_CTRL_U_ERR;  // RW/1C/V
} new_FWD_IP_t;

typedef struct packed {
    logic  [0:0] MA_TCN;  // RO/V
} new_FWD_IM_t;

typedef struct packed {
    new_FWD_IP_t  FWD_IP;
    new_FWD_IM_t  FWD_IM;
} mby_ppe_fwd_misc_map_new_t;

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

typedef logic [7:0] we_FWD_PORT_CFG_2_t;

typedef logic [7:0] we_FWD_LAG_CFG_t;

typedef logic [7:0] we_FWD_PORT_CFG_1_t;

typedef struct packed {
    we_FWD_PORT_CFG_2_t FWD_PORT_CFG_2;
    we_FWD_LAG_CFG_t FWD_LAG_CFG;
    we_FWD_PORT_CFG_1_t FWD_PORT_CFG_1;
} mby_ppe_fwd_misc_map_handcoded_t;

typedef logic [7:0] re_FWD_PORT_CFG_2_t;

typedef logic [7:0] re_FWD_LAG_CFG_t;

typedef logic [7:0] re_FWD_PORT_CFG_1_t;

typedef struct packed {
    re_FWD_PORT_CFG_2_t FWD_PORT_CFG_2;
    re_FWD_LAG_CFG_t FWD_LAG_CFG;
    re_FWD_PORT_CFG_1_t FWD_PORT_CFG_1;
} mby_ppe_fwd_misc_map_hc_re_t;

typedef logic handcode_rvalid_FWD_PORT_CFG_2_t;

typedef logic handcode_rvalid_FWD_LAG_CFG_t;

typedef logic handcode_rvalid_FWD_PORT_CFG_1_t;

typedef struct packed {
    handcode_rvalid_FWD_PORT_CFG_2_t FWD_PORT_CFG_2;
    handcode_rvalid_FWD_LAG_CFG_t FWD_LAG_CFG;
    handcode_rvalid_FWD_PORT_CFG_1_t FWD_PORT_CFG_1;
} mby_ppe_fwd_misc_map_hc_rvalid_t;

typedef logic handcode_wvalid_FWD_PORT_CFG_2_t;

typedef logic handcode_wvalid_FWD_LAG_CFG_t;

typedef logic handcode_wvalid_FWD_PORT_CFG_1_t;

typedef struct packed {
    handcode_wvalid_FWD_PORT_CFG_2_t FWD_PORT_CFG_2;
    handcode_wvalid_FWD_LAG_CFG_t FWD_LAG_CFG;
    handcode_wvalid_FWD_PORT_CFG_1_t FWD_PORT_CFG_1;
} mby_ppe_fwd_misc_map_hc_wvalid_t;

typedef logic handcode_error_FWD_PORT_CFG_2_t;

typedef logic handcode_error_FWD_LAG_CFG_t;

typedef logic handcode_error_FWD_PORT_CFG_1_t;

typedef struct packed {
    handcode_error_FWD_PORT_CFG_2_t FWD_PORT_CFG_2;
    handcode_error_FWD_LAG_CFG_t FWD_LAG_CFG;
    handcode_error_FWD_PORT_CFG_1_t FWD_PORT_CFG_1;
} mby_ppe_fwd_misc_map_hc_error_t;

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

typedef struct packed {
    FWD_PORT_CFG_2_t FWD_PORT_CFG_2;
    FWD_LAG_CFG_t FWD_LAG_CFG;
    FWD_PORT_CFG_1_t FWD_PORT_CFG_1;
} mby_ppe_fwd_misc_map_hc_reg_read_t;

typedef struct packed {
    FWD_PORT_CFG_2_t FWD_PORT_CFG_2;
    FWD_LAG_CFG_t FWD_LAG_CFG;
    FWD_PORT_CFG_1_t FWD_PORT_CFG_1;
} mby_ppe_fwd_misc_map_hc_reg_write_t;

// ===================================================
// RW/V2 Structure

// ===================================================
// Watch Signals Structure


endpackage: mby_ppe_fwd_misc_map_pkg

`endif // MBY_PPE_FWD_MISC_MAP_PKG_VH
