magic
tech scmos
timestamp 962519129
<< ndiffusion >>
rect 115 136 123 137
rect 115 130 123 134
rect 137 130 141 131
rect 115 124 123 128
rect 115 121 123 122
rect 115 117 117 121
rect 115 116 123 117
rect 137 124 141 128
rect 137 121 141 122
rect 137 116 141 117
rect 115 110 123 114
rect 137 110 141 114
rect 115 104 123 108
rect 137 107 141 108
rect 137 102 141 103
rect 115 101 123 102
rect 115 97 117 101
rect 115 96 123 97
rect 115 93 123 94
rect 119 90 123 93
rect 137 96 141 100
rect 137 93 141 94
rect 137 88 141 89
rect 137 82 141 86
rect 137 79 141 80
<< pdiffusion >>
rect 153 130 157 131
rect 171 130 183 131
rect 153 124 157 128
rect 171 124 183 128
rect 153 121 157 122
rect 153 116 157 117
rect 153 110 157 114
rect 171 121 183 122
rect 181 117 183 121
rect 171 116 183 117
rect 171 110 183 114
rect 153 107 157 108
rect 153 102 157 103
rect 171 107 183 108
rect 181 103 183 107
rect 171 102 183 103
rect 153 96 157 100
rect 171 99 183 100
rect 171 96 179 99
rect 153 93 157 94
rect 153 88 157 89
rect 153 82 157 86
rect 171 86 175 88
rect 171 82 183 86
rect 153 79 157 80
rect 171 79 183 80
<< ntransistor >>
rect 115 134 123 136
rect 115 128 123 130
rect 137 128 141 130
rect 115 122 123 124
rect 137 122 141 124
rect 115 114 123 116
rect 137 114 141 116
rect 115 108 123 110
rect 137 108 141 110
rect 115 102 123 104
rect 137 100 141 102
rect 115 94 123 96
rect 137 94 141 96
rect 137 86 141 88
rect 137 80 141 82
<< ptransistor >>
rect 153 128 157 130
rect 171 128 183 130
rect 153 122 157 124
rect 171 122 183 124
rect 153 114 157 116
rect 171 114 183 116
rect 153 108 157 110
rect 171 108 183 110
rect 153 100 157 102
rect 171 100 183 102
rect 153 94 157 96
rect 153 86 157 88
rect 153 80 157 82
rect 171 80 183 82
<< polysilicon >>
rect 112 134 115 136
rect 123 134 126 136
rect 112 128 115 130
rect 123 128 137 130
rect 141 128 153 130
rect 157 128 171 130
rect 183 128 186 130
rect 111 122 115 124
rect 123 122 126 124
rect 111 118 113 122
rect 129 116 131 128
rect 134 122 137 124
rect 141 122 153 124
rect 157 122 165 124
rect 168 122 171 124
rect 183 122 187 124
rect 113 114 115 116
rect 123 114 126 116
rect 129 114 137 116
rect 141 114 153 116
rect 157 114 160 116
rect 163 110 165 122
rect 185 118 187 122
rect 168 114 171 116
rect 183 114 185 116
rect 112 108 115 110
rect 123 108 137 110
rect 141 108 153 110
rect 157 108 171 110
rect 183 108 186 110
rect 112 102 115 104
rect 123 102 126 104
rect 129 100 137 102
rect 141 100 153 102
rect 157 100 160 102
rect 168 100 171 102
rect 183 100 187 102
rect 111 94 115 96
rect 123 94 126 96
rect 111 86 113 94
rect 129 88 131 100
rect 134 94 137 96
rect 141 94 153 96
rect 157 94 165 96
rect 129 86 137 88
rect 141 86 153 88
rect 157 86 160 88
rect 111 84 117 86
rect 163 82 165 94
rect 185 92 187 100
rect 181 90 187 92
rect 134 80 137 82
rect 141 80 153 82
rect 157 80 165 82
rect 168 80 171 82
rect 183 80 186 82
<< ndcontact >>
rect 115 137 123 141
rect 137 131 141 135
rect 117 117 123 121
rect 137 117 141 121
rect 137 103 141 107
rect 117 97 123 101
rect 115 89 119 93
rect 137 89 141 93
rect 137 75 141 79
<< pdcontact >>
rect 153 131 157 135
rect 171 131 183 135
rect 153 117 157 121
rect 171 117 181 121
rect 153 103 157 107
rect 171 103 181 107
rect 179 95 183 99
rect 153 89 157 93
rect 171 88 175 92
rect 153 75 157 79
rect 171 75 183 79
<< polycontact >>
rect 109 114 113 118
rect 185 114 189 118
rect 117 82 121 86
rect 177 88 181 92
<< metal1 >>
rect 115 137 123 141
rect 119 135 123 137
rect 119 131 141 135
rect 153 131 183 135
rect 109 114 113 118
rect 117 117 181 121
rect 110 93 113 114
rect 128 103 141 107
rect 128 101 132 103
rect 117 97 132 101
rect 145 93 149 117
rect 185 114 189 118
rect 153 103 181 107
rect 185 99 188 114
rect 179 95 188 99
rect 110 89 119 93
rect 137 92 157 93
rect 122 89 181 92
rect 110 79 113 89
rect 122 86 125 89
rect 171 88 181 89
rect 117 83 125 86
rect 185 85 188 95
rect 117 82 121 83
rect 129 82 188 85
rect 129 79 132 82
rect 110 76 132 79
rect 137 75 141 79
rect 153 75 183 79
<< labels >>
rlabel polysilicon 170 101 170 101 5 x
rlabel polysilicon 184 81 184 81 7 _PReset!
rlabel polysilicon 158 101 158 101 3 b
rlabel polysilicon 158 115 158 115 3 b
rlabel polysilicon 158 129 158 129 3 b
rlabel polysilicon 158 87 158 87 3 b
rlabel polysilicon 158 123 158 123 3 a
rlabel polysilicon 158 109 158 109 3 a
rlabel polysilicon 158 81 158 81 3 a
rlabel polysilicon 158 95 158 95 3 a
rlabel polysilicon 136 95 136 95 3 a
rlabel polysilicon 136 81 136 81 3 a
rlabel polysilicon 136 109 136 109 3 a
rlabel polysilicon 136 123 136 123 3 a
rlabel polysilicon 136 87 136 87 3 b
rlabel polysilicon 136 129 136 129 3 b
rlabel polysilicon 136 115 136 115 3 b
rlabel polysilicon 136 101 136 101 3 b
rlabel polysilicon 114 103 114 103 1 _SReset!
rlabel polysilicon 124 95 124 95 5 x
rlabel polysilicon 114 135 114 135 3 _SReset!
rlabel space 109 74 138 142 7 ^n
rlabel space 156 74 189 136 3 ^p
rlabel pdcontact 177 133 177 133 5 Vdd!
rlabel pdcontact 177 77 177 77 1 Vdd!
rlabel pdcontact 176 105 176 105 1 Vdd!
rlabel pdcontact 176 119 176 119 1 x
rlabel pdcontact 155 77 155 77 1 Vdd!
rlabel pdcontact 155 133 155 133 5 Vdd!
rlabel pdcontact 155 119 155 119 1 x
rlabel pdcontact 155 91 155 91 1 x
rlabel pdcontact 155 105 155 105 1 Vdd!
rlabel ndcontact 139 105 139 105 1 GND!
rlabel ndcontact 139 91 139 91 1 x
rlabel ndcontact 139 119 139 119 1 x
rlabel ndcontact 139 77 139 77 1 GND!
rlabel ndcontact 139 133 139 133 5 GND!
rlabel ndcontact 120 99 120 99 1 GND!
rlabel ndcontact 120 119 120 119 1 x
rlabel ndcontact 119 139 119 139 5 GND!
<< end >>
