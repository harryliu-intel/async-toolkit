.SUBCKT g1ibd08ffaa0d08x5  
.ENDS g1ibd08ffaa0d08x5

.SUBCKT g1iclkbfiaa2n06x5  
.ENDS g1iclkbfiaa2n06x5

.SUBCKT g1ictree2aa2n04x5  
.ENDS g1ictree2aa2n04x5

.SUBCKT g1idivertaa2d04x5  
.ENDS g1idivertaa2d04x5

.SUBCKT g1icutsnkaa2n04x5  
.ENDS g1icutsnkaa2n04x5

.SUBCKT g1ixor002aa2n04x5  
.ENDS g1ixor002aa2n04x5

.SUBCKT g1itd1004aa0d04x5  
.ENDS g1itd1004aa0d04x5

.SUBCKT g1itd1008aa0d04x5  
.ENDS g1itd1008aa0d04x5

.SUBCKT g1itilo00aa2n02x5  
.ENDS g1itilo00aa2n02x5

.SUBCKT g1itihi00aa2n02x5  
.ENDS g1itihi00aa2n02x5

.SUBCKT g1idl1006aa0d04x5  
.ENDS g1idl1006aa0d04x5

.SUBCKT g1ibd07ffaa0d08x5  
.ENDS g1ibd07ffaa0d08x5

.SUBCKT g1ibfn000aa2n12x5  
.ENDS g1ibfn000aa2n12x5

.SUBCKT g1ilsn000aa2n04x5  
.ENDS g1ilsn000aa2n04x5

.SUBCKT g1idl1004aa0d04x5  
.ENDS g1idl1004aa0d04x5

.SUBCKT g1ibfn000aa2n24x5  
.ENDS g1ibfn000aa2n24x5

.SUBCKT g1ibfn000aa2n08x5  
.ENDS g1ibfn000aa2n08x5

.SUBCKT g1iltny00aa2n02x5  
.ENDS g1iltny00aa2n02x5

.SUBCKT g1ibfn000aa2n02x5  
.ENDS g1ibfn000aa2n02x5

.SUBCKT g1ibfn000aa2n04x5  
.ENDS g1ibfn000aa2n04x5

.SUBCKT g1ixor002aa2n02x5  
.ENDS g1ixor002aa2n02x5

.SUBCKT g1iand002aa2n02x5  
.ENDS g1iand002aa2n02x5

.SUBCKT g1ixnr002aa2n02x5  
.ENDS g1ixnr002aa2n02x5

.SUBCKT g1iorn002aa2n02x5  
.ENDS g1iorn002aa2n02x5

.SUBCKT g1irm0023aa2d02x5  
.ENDS g1irm0023aa2d02x5

.SUBCKT g1ixor003ba2n01x1  
.ENDS g1ixor003ba2n01x1

.SUBCKT g1imbn022aa2n01x1  
.ENDS g1imbn022aa2n01x1

.SUBCKT g1iaoi012aa2n02x5  
.ENDS g1iaoi012aa2n02x5

.SUBCKT g1ioai012aa2n02x5  
.ENDS g1ioai012aa2n02x5

.SUBCKT g1ikpginvaa2n01x5  
.ENDS g1ikpginvaa2n01x5

.SUBCKT g1ikpgcmbaa2n02x5  
.ENDS g1ikpgcmbaa2n02x5

.SUBCKT g1ioai012aa2n01x1  
.ENDS g1ioai012aa2n01x1

.SUBCKT g1iaoi012aa2n01x1  
.ENDS g1iaoi012aa2n01x1

.SUBCKT g1iinv000aa2n02x5  
.ENDS g1iinv000aa2n02x5

.SUBCKT g1ikpgencaa2n02x5  
.ENDS g1ikpgencaa2n02x5

.SUBCKT g1inorb02aa2n01x1  
.ENDS g1inorb02aa2n01x1

.SUBCKT g1ixor002aa2n01x1  
.ENDS g1ixor002aa2n01x1

.SUBCKT g1ixnr002aa2n01x1  
.ENDS g1ixnr002aa2n01x1

.SUBCKT g1ikpgcmbaa2n01x5  
.ENDS g1ikpgcmbaa2n01x5

.SUBCKT g1ioao003aa2n02x5  
.ENDS g1ioao003aa2n02x5

.SUBCKT g1ibfm201aa2n02x5  
.ENDS g1ibfm201aa2n02x5

.SUBCKT g1ibfm201aa2n04x5  
.ENDS g1ibfm201aa2n04x5

.SUBCKT g1iltny00aa2n01x5  
.ENDS g1iltny00aa2n01x5

.SUBCKT core_D_crypto_D_bitcoin_D_stage_D_TEST_U_4_U_STAGES_D_1000  
.ENDS core_D_crypto_D_bitcoin_D_stage_D_TEST_U_4_U_STAGES_D_1000

