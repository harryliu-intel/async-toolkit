magic
tech scmos
timestamp 965421252
use s_c2 s_c2_0
timestamp 962795507
transform 1 0 -76 0 1 -22
box -112 289 -70 318
use m_c2 m_c2_0
timestamp 963604341
transform 1 0 254 0 1 -49
box -157 315 3 367
use l_c2 l_c2_0
timestamp 965420547
transform 1 0 392 0 1 280
box -43 -15 83 80
use s_c2_rhi s_c2_rhi_0
timestamp 965421252
transform 1 0 -34 0 1 58
box -154 65 13 102
use m_c2_rhi m_c2_rhi_0
timestamp 964630225
transform 1 0 176 0 1 105
box -79 17 81 85
use l_c2_rhi l_c2_rhi_0
timestamp 965420787
transform 1 0 289 0 1 179
box 59 -57 186 69
use s_c2_phi s_c2_phi_0
timestamp 965421252
transform 1 0 -63 0 1 -103
box -125 85 37 120
use m_c2_phi m_c2_phi_0
timestamp 963604341
transform 1 0 124 0 1 -43
box -27 24 133 92
use l_c2_phi l_c2_phi_0
timestamp 965420787
transform 1 0 263 0 1 -47
box 84 44 213 138
use s_2and2c2 s_2and2c2_0
timestamp 965071231
transform 1 0 -63 0 1 -299
box -126 90 -62 152
use m_2and2c2 m_2and2c2_0
timestamp 965071348
transform 1 0 91 0 1 -218
box 6 9 120 137
use s_2and2c2_rhi s_2and2c2_rhi_0
timestamp 965421252
transform 1 0 -12 0 1 -500
box -177 91 18 154
use m_2and2c2_rhi m_2and2c2_rhi_0
timestamp 965071231
transform 1 0 -22 0 1 -439
box 119 30 246 172
use s_and2c2 s_and2c2_0
timestamp 965071231
transform 1 0 -55 0 1 -1104
box -134 548 -70 597
use m_and2c2 m_and2c2_0
timestamp 965071231
transform 1 0 101 0 1 -585
box -4 29 121 140
use s_and2c2_rhi s_and2c2_rhi_0
timestamp 965421252
transform 1 0 -24 0 1 -1261
box -165 560 21 615
use m_and2c2_rhi m_and2c2_rhi_0
timestamp 965071231
transform 1 0 123 0 1 -747
box -26 46 115 160
use l_and2c2_rhi l_and2c2_rhi_0
timestamp 964081429
transform 1 0 258 0 1 -702
box 79 -2 244 165
<< end >>
