///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_trig_apply_misc_map.sv                             
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_trig_apply_misc_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_RSTD


module rtlgen_mby_ppe_trig_apply_misc_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_trig_apply_misc_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_PH2_FF
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_trig_apply_misc_map ( //lintra s-2096
    // Clocks
    gated_clk,
    rtl_clk,

    // Resets
    rst_n,


    // Register Inputs
    load_MA_TCN_IP,
    load_TRIGGER_IP,

    new_MA_TCN_IP,
    new_TRIGGER_IP,
    new_TRIGGER_RATE_LIM_EMPTY,

    handcode_reg_rdata_MA_TCN_DATA_0,
    handcode_reg_rdata_MA_TCN_DATA_1,
    handcode_reg_rdata_MA_TCN_DEQUEUE,
    handcode_reg_rdata_MA_TCN_FIFO_0,
    handcode_reg_rdata_MA_TCN_FIFO_1,
    handcode_reg_rdata_MA_TCN_PTR_HEAD,
    handcode_reg_rdata_MA_TCN_PTR_TAIL,
    handcode_reg_rdata_TRIGGER_ACTION_METADATA_MASK,
    handcode_reg_rdata_TRIGGER_RATE_LIM_CFG_2,

    handcode_rvalid_MA_TCN_DATA_0,
    handcode_rvalid_MA_TCN_DATA_1,
    handcode_rvalid_MA_TCN_DEQUEUE,
    handcode_rvalid_MA_TCN_FIFO_0,
    handcode_rvalid_MA_TCN_FIFO_1,
    handcode_rvalid_MA_TCN_PTR_HEAD,
    handcode_rvalid_MA_TCN_PTR_TAIL,
    handcode_rvalid_TRIGGER_ACTION_METADATA_MASK,
    handcode_rvalid_TRIGGER_RATE_LIM_CFG_2,

    handcode_wvalid_MA_TCN_DATA_0,
    handcode_wvalid_MA_TCN_DATA_1,
    handcode_wvalid_MA_TCN_DEQUEUE,
    handcode_wvalid_MA_TCN_FIFO_0,
    handcode_wvalid_MA_TCN_FIFO_1,
    handcode_wvalid_MA_TCN_PTR_HEAD,
    handcode_wvalid_MA_TCN_PTR_TAIL,
    handcode_wvalid_TRIGGER_ACTION_METADATA_MASK,
    handcode_wvalid_TRIGGER_RATE_LIM_CFG_2,

    handcode_error_MA_TCN_DATA_0,
    handcode_error_MA_TCN_DATA_1,
    handcode_error_MA_TCN_DEQUEUE,
    handcode_error_MA_TCN_FIFO_0,
    handcode_error_MA_TCN_FIFO_1,
    handcode_error_MA_TCN_PTR_HEAD,
    handcode_error_MA_TCN_PTR_TAIL,
    handcode_error_TRIGGER_ACTION_METADATA_MASK,
    handcode_error_TRIGGER_RATE_LIM_CFG_2,


    // Register Outputs
    MA_TCN_IM,
    MA_TCN_IP,
    MA_TCN_USAGE,
    MA_TCN_WM,
    TRIGGER_IM,
    TRIGGER_IP,
    TRIGGER_RATE_LIM_EMPTY,


    // Register signals for HandCoded registers
    handcode_reg_wdata_MA_TCN_DATA_0,
    handcode_reg_wdata_MA_TCN_DATA_1,
    handcode_reg_wdata_MA_TCN_DEQUEUE,
    handcode_reg_wdata_MA_TCN_FIFO_0,
    handcode_reg_wdata_MA_TCN_FIFO_1,
    handcode_reg_wdata_MA_TCN_PTR_HEAD,
    handcode_reg_wdata_MA_TCN_PTR_TAIL,
    handcode_reg_wdata_TRIGGER_ACTION_METADATA_MASK,
    handcode_reg_wdata_TRIGGER_RATE_LIM_CFG_2,

    we_MA_TCN_DATA_0,
    we_MA_TCN_DATA_1,
    we_MA_TCN_DEQUEUE,
    we_MA_TCN_FIFO_0,
    we_MA_TCN_FIFO_1,
    we_MA_TCN_PTR_HEAD,
    we_MA_TCN_PTR_TAIL,
    we_TRIGGER_ACTION_METADATA_MASK,
    we_TRIGGER_RATE_LIM_CFG_2,

    re_MA_TCN_DATA_0,
    re_MA_TCN_DATA_1,
    re_MA_TCN_DEQUEUE,
    re_MA_TCN_FIFO_0,
    re_MA_TCN_FIFO_1,
    re_MA_TCN_PTR_HEAD,
    re_MA_TCN_PTR_TAIL,
    re_TRIGGER_ACTION_METADATA_MASK,
    re_TRIGGER_RATE_LIM_CFG_2,




    // Config Access
    req,
    ack
    

);

import mby_ppe_trig_apply_misc_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:0] MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET = {MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] TRIG_APPLY_MISC_SB_BAR = 3'b0;
parameter [7:0] TRIG_APPLY_MISC_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
`define TRIGGER_IP_CR_ADDR_def(INDEX) TRIGGER_IP_CR_ADDR``INDEX``[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
`define TRIGGER_IM_CR_ADDR_def(INDEX) TRIGGER_IM_CR_ADDR``INDEX``[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
`define MA_TCN_WM_CR_ADDR_def(INDEX) MA_TCN_WM_CR_ADDR``INDEX``[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
`define MA_TCN_USAGE_CR_ADDR_def(INDEX) MA_TCN_USAGE_CR_ADDR``INDEX``[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]
localparam [1:0][MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] TRIGGER_IP_DECODE_ADDR = {`TRIGGER_IP_CR_ADDR_def([1]),`TRIGGER_IP_CR_ADDR_def([0])};
localparam [1:0][MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] TRIGGER_IM_DECODE_ADDR = {`TRIGGER_IM_CR_ADDR_def([1]),`TRIGGER_IM_CR_ADDR_def([0])};
localparam [MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] TRIGGER_RATE_LIM_EMPTY_DECODE_ADDR = TRIGGER_RATE_LIM_EMPTY_CR_ADDR[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MA_TCN_IP_DECODE_ADDR = MA_TCN_IP_CR_ADDR[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MA_TCN_IM_DECODE_ADDR = MA_TCN_IM_CR_ADDR[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_TRIG_APPLY_MISC_MAP_OFFSET[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [16:0][MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MA_TCN_WM_DECODE_ADDR = {`MA_TCN_WM_CR_ADDR_def([16]),`MA_TCN_WM_CR_ADDR_def([15]),`MA_TCN_WM_CR_ADDR_def([14]),`MA_TCN_WM_CR_ADDR_def([13]),`MA_TCN_WM_CR_ADDR_def([12]),`MA_TCN_WM_CR_ADDR_def([11]),`MA_TCN_WM_CR_ADDR_def([10]),`MA_TCN_WM_CR_ADDR_def([9]),`MA_TCN_WM_CR_ADDR_def([8]),`MA_TCN_WM_CR_ADDR_def([7]),`MA_TCN_WM_CR_ADDR_def([6]),`MA_TCN_WM_CR_ADDR_def([5]),`MA_TCN_WM_CR_ADDR_def([4]),`MA_TCN_WM_CR_ADDR_def([3]),`MA_TCN_WM_CR_ADDR_def([2]),`MA_TCN_WM_CR_ADDR_def([1]),`MA_TCN_WM_CR_ADDR_def([0])};
localparam [16:0][MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MA_TCN_USAGE_DECODE_ADDR = {`MA_TCN_USAGE_CR_ADDR_def([16]),`MA_TCN_USAGE_CR_ADDR_def([15]),`MA_TCN_USAGE_CR_ADDR_def([14]),`MA_TCN_USAGE_CR_ADDR_def([13]),`MA_TCN_USAGE_CR_ADDR_def([12]),`MA_TCN_USAGE_CR_ADDR_def([11]),`MA_TCN_USAGE_CR_ADDR_def([10]),`MA_TCN_USAGE_CR_ADDR_def([9]),`MA_TCN_USAGE_CR_ADDR_def([8]),`MA_TCN_USAGE_CR_ADDR_def([7]),`MA_TCN_USAGE_CR_ADDR_def([6]),`MA_TCN_USAGE_CR_ADDR_def([5]),`MA_TCN_USAGE_CR_ADDR_def([4]),`MA_TCN_USAGE_CR_ADDR_def([3]),`MA_TCN_USAGE_CR_ADDR_def([2]),`MA_TCN_USAGE_CR_ADDR_def([1]),`MA_TCN_USAGE_CR_ADDR_def([0])};

    // Clocks
input logic  gated_clk;
input logic  rtl_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input load_MA_TCN_IP_t  load_MA_TCN_IP;
input load_TRIGGER_IP_t [1:0] load_TRIGGER_IP;

input new_MA_TCN_IP_t  new_MA_TCN_IP;
input new_TRIGGER_IP_t [1:0] new_TRIGGER_IP;
input new_TRIGGER_RATE_LIM_EMPTY_t  new_TRIGGER_RATE_LIM_EMPTY;

input MA_TCN_DATA_0_t  handcode_reg_rdata_MA_TCN_DATA_0;
input MA_TCN_DATA_1_t  handcode_reg_rdata_MA_TCN_DATA_1;
input MA_TCN_DEQUEUE_t  handcode_reg_rdata_MA_TCN_DEQUEUE;
input MA_TCN_FIFO_0_t  handcode_reg_rdata_MA_TCN_FIFO_0;
input MA_TCN_FIFO_1_t  handcode_reg_rdata_MA_TCN_FIFO_1;
input MA_TCN_PTR_HEAD_t  handcode_reg_rdata_MA_TCN_PTR_HEAD;
input MA_TCN_PTR_TAIL_t  handcode_reg_rdata_MA_TCN_PTR_TAIL;
input TRIGGER_ACTION_METADATA_MASK_t  handcode_reg_rdata_TRIGGER_ACTION_METADATA_MASK;
input TRIGGER_RATE_LIM_CFG_2_t  handcode_reg_rdata_TRIGGER_RATE_LIM_CFG_2;

input handcode_rvalid_MA_TCN_DATA_0_t  handcode_rvalid_MA_TCN_DATA_0;
input handcode_rvalid_MA_TCN_DATA_1_t  handcode_rvalid_MA_TCN_DATA_1;
input handcode_rvalid_MA_TCN_DEQUEUE_t  handcode_rvalid_MA_TCN_DEQUEUE;
input handcode_rvalid_MA_TCN_FIFO_0_t  handcode_rvalid_MA_TCN_FIFO_0;
input handcode_rvalid_MA_TCN_FIFO_1_t  handcode_rvalid_MA_TCN_FIFO_1;
input handcode_rvalid_MA_TCN_PTR_HEAD_t  handcode_rvalid_MA_TCN_PTR_HEAD;
input handcode_rvalid_MA_TCN_PTR_TAIL_t  handcode_rvalid_MA_TCN_PTR_TAIL;
input handcode_rvalid_TRIGGER_ACTION_METADATA_MASK_t  handcode_rvalid_TRIGGER_ACTION_METADATA_MASK;
input handcode_rvalid_TRIGGER_RATE_LIM_CFG_2_t  handcode_rvalid_TRIGGER_RATE_LIM_CFG_2;

input handcode_wvalid_MA_TCN_DATA_0_t  handcode_wvalid_MA_TCN_DATA_0;
input handcode_wvalid_MA_TCN_DATA_1_t  handcode_wvalid_MA_TCN_DATA_1;
input handcode_wvalid_MA_TCN_DEQUEUE_t  handcode_wvalid_MA_TCN_DEQUEUE;
input handcode_wvalid_MA_TCN_FIFO_0_t  handcode_wvalid_MA_TCN_FIFO_0;
input handcode_wvalid_MA_TCN_FIFO_1_t  handcode_wvalid_MA_TCN_FIFO_1;
input handcode_wvalid_MA_TCN_PTR_HEAD_t  handcode_wvalid_MA_TCN_PTR_HEAD;
input handcode_wvalid_MA_TCN_PTR_TAIL_t  handcode_wvalid_MA_TCN_PTR_TAIL;
input handcode_wvalid_TRIGGER_ACTION_METADATA_MASK_t  handcode_wvalid_TRIGGER_ACTION_METADATA_MASK;
input handcode_wvalid_TRIGGER_RATE_LIM_CFG_2_t  handcode_wvalid_TRIGGER_RATE_LIM_CFG_2;

input handcode_error_MA_TCN_DATA_0_t  handcode_error_MA_TCN_DATA_0;
input handcode_error_MA_TCN_DATA_1_t  handcode_error_MA_TCN_DATA_1;
input handcode_error_MA_TCN_DEQUEUE_t  handcode_error_MA_TCN_DEQUEUE;
input handcode_error_MA_TCN_FIFO_0_t  handcode_error_MA_TCN_FIFO_0;
input handcode_error_MA_TCN_FIFO_1_t  handcode_error_MA_TCN_FIFO_1;
input handcode_error_MA_TCN_PTR_HEAD_t  handcode_error_MA_TCN_PTR_HEAD;
input handcode_error_MA_TCN_PTR_TAIL_t  handcode_error_MA_TCN_PTR_TAIL;
input handcode_error_TRIGGER_ACTION_METADATA_MASK_t  handcode_error_TRIGGER_ACTION_METADATA_MASK;
input handcode_error_TRIGGER_RATE_LIM_CFG_2_t  handcode_error_TRIGGER_RATE_LIM_CFG_2;


    // Register Outputs
output MA_TCN_IM_t  MA_TCN_IM;
output MA_TCN_IP_t  MA_TCN_IP;
output MA_TCN_USAGE_t [16:0] MA_TCN_USAGE;
output MA_TCN_WM_t [16:0] MA_TCN_WM;
output TRIGGER_IM_t [1:0] TRIGGER_IM;
output TRIGGER_IP_t [1:0] TRIGGER_IP;
output TRIGGER_RATE_LIM_EMPTY_t  TRIGGER_RATE_LIM_EMPTY;


    // Register signals for HandCoded registers
output MA_TCN_DATA_0_t  handcode_reg_wdata_MA_TCN_DATA_0;
output MA_TCN_DATA_1_t  handcode_reg_wdata_MA_TCN_DATA_1;
output MA_TCN_DEQUEUE_t  handcode_reg_wdata_MA_TCN_DEQUEUE;
output MA_TCN_FIFO_0_t  handcode_reg_wdata_MA_TCN_FIFO_0;
output MA_TCN_FIFO_1_t  handcode_reg_wdata_MA_TCN_FIFO_1;
output MA_TCN_PTR_HEAD_t  handcode_reg_wdata_MA_TCN_PTR_HEAD;
output MA_TCN_PTR_TAIL_t  handcode_reg_wdata_MA_TCN_PTR_TAIL;
output TRIGGER_ACTION_METADATA_MASK_t  handcode_reg_wdata_TRIGGER_ACTION_METADATA_MASK;
output TRIGGER_RATE_LIM_CFG_2_t  handcode_reg_wdata_TRIGGER_RATE_LIM_CFG_2;

output we_MA_TCN_DATA_0_t  we_MA_TCN_DATA_0;
output we_MA_TCN_DATA_1_t  we_MA_TCN_DATA_1;
output we_MA_TCN_DEQUEUE_t  we_MA_TCN_DEQUEUE;
output we_MA_TCN_FIFO_0_t  we_MA_TCN_FIFO_0;
output we_MA_TCN_FIFO_1_t  we_MA_TCN_FIFO_1;
output we_MA_TCN_PTR_HEAD_t  we_MA_TCN_PTR_HEAD;
output we_MA_TCN_PTR_TAIL_t  we_MA_TCN_PTR_TAIL;
output we_TRIGGER_ACTION_METADATA_MASK_t  we_TRIGGER_ACTION_METADATA_MASK;
output we_TRIGGER_RATE_LIM_CFG_2_t  we_TRIGGER_RATE_LIM_CFG_2;

output re_MA_TCN_DATA_0_t  re_MA_TCN_DATA_0;
output re_MA_TCN_DATA_1_t  re_MA_TCN_DATA_1;
output re_MA_TCN_DEQUEUE_t  re_MA_TCN_DEQUEUE;
output re_MA_TCN_FIFO_0_t  re_MA_TCN_FIFO_0;
output re_MA_TCN_FIFO_1_t  re_MA_TCN_FIFO_1;
output re_MA_TCN_PTR_HEAD_t  re_MA_TCN_PTR_HEAD;
output re_MA_TCN_PTR_TAIL_t  re_MA_TCN_PTR_TAIL;
output re_TRIGGER_ACTION_METADATA_MASK_t  re_TRIGGER_ACTION_METADATA_MASK;
output re_TRIGGER_RATE_LIM_CFG_2_t  re_TRIGGER_RATE_LIM_CFG_2;




    // Config Access
input mby_ppe_trig_apply_misc_map_cr_req_t  req;
output mby_ppe_trig_apply_misc_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_trig_apply_misc_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_TRIG_APPLY_MISC_MAP_MEM;
assign case_req_addr_MBY_PPE_TRIG_APPLY_MISC_MAP_MEM = req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_trig_apply_misc;
always_comb begin : sb_fid_cond_trig_apply_misc_BLOCK
    unique casez (req_fid) 
		TRIG_APPLY_MISC_SB_FID: sb_fid_cond_trig_apply_misc = 1;
		default: sb_fid_cond_trig_apply_misc = 0;
    endcase 
end


logic sb_bar_cond_trig_apply_misc;
always_comb begin : sb_bar_cond_trig_apply_misc_BLOCK
    unique casez (req_bar) 
		TRIG_APPLY_MISC_SB_BAR: sb_bar_cond_trig_apply_misc = 1;
		default: sb_bar_cond_trig_apply_misc = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// TRIGGER_RATE_LIM_CFG_2 using HANDCODED_REG template.
logic addr_decode_TRIGGER_RATE_LIM_CFG_2;
logic write_req_TRIGGER_RATE_LIM_CFG_2;
logic read_req_TRIGGER_RATE_LIM_CFG_2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'b0???,1'b?}: 
         addr_decode_TRIGGER_RATE_LIM_CFG_2 = req.valid;
      default: 
         addr_decode_TRIGGER_RATE_LIM_CFG_2 = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_RATE_LIM_CFG_2 = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_RATE_LIM_CFG_2 ;
always_comb read_req_TRIGGER_RATE_LIM_CFG_2  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_RATE_LIM_CFG_2 ;

always_comb we_TRIGGER_RATE_LIM_CFG_2 = {8{write_req_TRIGGER_RATE_LIM_CFG_2}} & be;
always_comb re_TRIGGER_RATE_LIM_CFG_2 = {8{read_req_TRIGGER_RATE_LIM_CFG_2}} & be;
always_comb handcode_reg_wdata_TRIGGER_RATE_LIM_CFG_2 = write_data;


// ----------------------------------------------------------------------
// TRIGGER_ACTION_METADATA_MASK using HANDCODED_REG template.
logic addr_decode_TRIGGER_ACTION_METADATA_MASK;
logic write_req_TRIGGER_ACTION_METADATA_MASK;
logic read_req_TRIGGER_ACTION_METADATA_MASK;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'b10??,1'b?}: 
         addr_decode_TRIGGER_ACTION_METADATA_MASK = req.valid;
      default: 
         addr_decode_TRIGGER_ACTION_METADATA_MASK = 1'b0; 
   endcase
end

always_comb write_req_TRIGGER_ACTION_METADATA_MASK = f_IsMEMWr(req_opcode) && addr_decode_TRIGGER_ACTION_METADATA_MASK ;
always_comb read_req_TRIGGER_ACTION_METADATA_MASK  = f_IsMEMRd(req_opcode) && addr_decode_TRIGGER_ACTION_METADATA_MASK ;

always_comb we_TRIGGER_ACTION_METADATA_MASK = {8{write_req_TRIGGER_ACTION_METADATA_MASK}} & be;
always_comb re_TRIGGER_ACTION_METADATA_MASK = {8{read_req_TRIGGER_ACTION_METADATA_MASK}} & be;
always_comb handcode_reg_wdata_TRIGGER_ACTION_METADATA_MASK = write_data;


//---------------------------------------------------------------------
// TRIGGER_IP Address Decode
logic [1:0] addr_decode_TRIGGER_IP;
logic [1:0] write_req_TRIGGER_IP;
always_comb begin
   addr_decode_TRIGGER_IP[0] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == TRIGGER_IP_DECODE_ADDR[0]) && req.valid ;
   addr_decode_TRIGGER_IP[1] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == TRIGGER_IP_DECODE_ADDR[1]) && req.valid ;
   write_req_TRIGGER_IP[0] = IsMEMWr && addr_decode_TRIGGER_IP[0] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_TRIGGER_IP[1] = IsMEMWr && addr_decode_TRIGGER_IP[1] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
end

// ----------------------------------------------------------------------
// TRIGGER_IP.PENDING x8 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [1:0][47:0] req_up_TRIGGER_IP_PENDING;
always_comb begin
 req_up_TRIGGER_IP_PENDING[0][7:0] = 
   {8{write_req_TRIGGER_IP[0] & be[0]}}
;
 req_up_TRIGGER_IP_PENDING[0][15:8] = 
   {8{write_req_TRIGGER_IP[0] & be[1]}}
;
 req_up_TRIGGER_IP_PENDING[0][23:16] = 
   {8{write_req_TRIGGER_IP[0] & be[2]}}
;
 req_up_TRIGGER_IP_PENDING[0][31:24] = 
   {8{write_req_TRIGGER_IP[0] & be[3]}}
;
 req_up_TRIGGER_IP_PENDING[0][39:32] = 
   {8{write_req_TRIGGER_IP[0] & be[4]}}
;
 req_up_TRIGGER_IP_PENDING[0][47:40] = 
   {8{write_req_TRIGGER_IP[0] & be[5]}}
;
 req_up_TRIGGER_IP_PENDING[1][7:0] = 
   {8{write_req_TRIGGER_IP[1] & be[0]}}
;
 req_up_TRIGGER_IP_PENDING[1][15:8] = 
   {8{write_req_TRIGGER_IP[1] & be[1]}}
;
 req_up_TRIGGER_IP_PENDING[1][23:16] = 
   {8{write_req_TRIGGER_IP[1] & be[2]}}
;
 req_up_TRIGGER_IP_PENDING[1][31:24] = 
   {8{write_req_TRIGGER_IP[1] & be[3]}}
;
 req_up_TRIGGER_IP_PENDING[1][39:32] = 
   {8{write_req_TRIGGER_IP[1] & be[4]}}
;
 req_up_TRIGGER_IP_PENDING[1][47:40] = 
   {8{write_req_TRIGGER_IP[1] & be[5]}}
;
end

logic [1:0][47:0] clr_TRIGGER_IP_PENDING;
always_comb begin
 clr_TRIGGER_IP_PENDING[0] = write_data[47:0] & req_up_TRIGGER_IP_PENDING[0];

 clr_TRIGGER_IP_PENDING[1] = write_data[47:0] & req_up_TRIGGER_IP_PENDING[1];

end
logic [1:0][47:0] swwr_TRIGGER_IP_PENDING;
logic [1:0][47:0] sw_nxt_TRIGGER_IP_PENDING;
always_comb begin
 swwr_TRIGGER_IP_PENDING[0] = clr_TRIGGER_IP_PENDING[0];
 sw_nxt_TRIGGER_IP_PENDING[0] = {48{1'b0}};

 swwr_TRIGGER_IP_PENDING[1] = clr_TRIGGER_IP_PENDING[1];
 sw_nxt_TRIGGER_IP_PENDING[1] = {48{1'b0}};

end
logic [1:0][47:0] up_TRIGGER_IP_PENDING;
logic [1:0][47:0] nxt_TRIGGER_IP_PENDING;
always_comb begin
 up_TRIGGER_IP_PENDING[0] = 
   swwr_TRIGGER_IP_PENDING[0] | {48{load_TRIGGER_IP[0].PENDING}};
 up_TRIGGER_IP_PENDING[1] = 
   swwr_TRIGGER_IP_PENDING[1] | {48{load_TRIGGER_IP[1].PENDING}};
end
always_comb begin
 nxt_TRIGGER_IP_PENDING[0][0] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[0] :
    sw_nxt_TRIGGER_IP_PENDING[0][0];
 nxt_TRIGGER_IP_PENDING[0][1] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[1] :
    sw_nxt_TRIGGER_IP_PENDING[0][1];
 nxt_TRIGGER_IP_PENDING[0][2] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[2] :
    sw_nxt_TRIGGER_IP_PENDING[0][2];
 nxt_TRIGGER_IP_PENDING[0][3] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[3] :
    sw_nxt_TRIGGER_IP_PENDING[0][3];
 nxt_TRIGGER_IP_PENDING[0][4] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[4] :
    sw_nxt_TRIGGER_IP_PENDING[0][4];
 nxt_TRIGGER_IP_PENDING[0][5] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[5] :
    sw_nxt_TRIGGER_IP_PENDING[0][5];
 nxt_TRIGGER_IP_PENDING[0][6] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[6] :
    sw_nxt_TRIGGER_IP_PENDING[0][6];
 nxt_TRIGGER_IP_PENDING[0][7] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[7] :
    sw_nxt_TRIGGER_IP_PENDING[0][7];
 nxt_TRIGGER_IP_PENDING[0][8] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[8] :
    sw_nxt_TRIGGER_IP_PENDING[0][8];
 nxt_TRIGGER_IP_PENDING[0][9] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[9] :
    sw_nxt_TRIGGER_IP_PENDING[0][9];
 nxt_TRIGGER_IP_PENDING[0][10] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[10] :
    sw_nxt_TRIGGER_IP_PENDING[0][10];
 nxt_TRIGGER_IP_PENDING[0][11] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[11] :
    sw_nxt_TRIGGER_IP_PENDING[0][11];
 nxt_TRIGGER_IP_PENDING[0][12] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[12] :
    sw_nxt_TRIGGER_IP_PENDING[0][12];
 nxt_TRIGGER_IP_PENDING[0][13] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[13] :
    sw_nxt_TRIGGER_IP_PENDING[0][13];
 nxt_TRIGGER_IP_PENDING[0][14] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[14] :
    sw_nxt_TRIGGER_IP_PENDING[0][14];
 nxt_TRIGGER_IP_PENDING[0][15] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[15] :
    sw_nxt_TRIGGER_IP_PENDING[0][15];
 nxt_TRIGGER_IP_PENDING[0][16] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[16] :
    sw_nxt_TRIGGER_IP_PENDING[0][16];
 nxt_TRIGGER_IP_PENDING[0][17] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[17] :
    sw_nxt_TRIGGER_IP_PENDING[0][17];
 nxt_TRIGGER_IP_PENDING[0][18] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[18] :
    sw_nxt_TRIGGER_IP_PENDING[0][18];
 nxt_TRIGGER_IP_PENDING[0][19] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[19] :
    sw_nxt_TRIGGER_IP_PENDING[0][19];
 nxt_TRIGGER_IP_PENDING[0][20] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[20] :
    sw_nxt_TRIGGER_IP_PENDING[0][20];
 nxt_TRIGGER_IP_PENDING[0][21] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[21] :
    sw_nxt_TRIGGER_IP_PENDING[0][21];
 nxt_TRIGGER_IP_PENDING[0][22] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[22] :
    sw_nxt_TRIGGER_IP_PENDING[0][22];
 nxt_TRIGGER_IP_PENDING[0][23] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[23] :
    sw_nxt_TRIGGER_IP_PENDING[0][23];
 nxt_TRIGGER_IP_PENDING[0][24] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[24] :
    sw_nxt_TRIGGER_IP_PENDING[0][24];
 nxt_TRIGGER_IP_PENDING[0][25] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[25] :
    sw_nxt_TRIGGER_IP_PENDING[0][25];
 nxt_TRIGGER_IP_PENDING[0][26] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[26] :
    sw_nxt_TRIGGER_IP_PENDING[0][26];
 nxt_TRIGGER_IP_PENDING[0][27] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[27] :
    sw_nxt_TRIGGER_IP_PENDING[0][27];
 nxt_TRIGGER_IP_PENDING[0][28] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[28] :
    sw_nxt_TRIGGER_IP_PENDING[0][28];
 nxt_TRIGGER_IP_PENDING[0][29] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[29] :
    sw_nxt_TRIGGER_IP_PENDING[0][29];
 nxt_TRIGGER_IP_PENDING[0][30] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[30] :
    sw_nxt_TRIGGER_IP_PENDING[0][30];
 nxt_TRIGGER_IP_PENDING[0][31] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[31] :
    sw_nxt_TRIGGER_IP_PENDING[0][31];
 nxt_TRIGGER_IP_PENDING[0][32] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[32] :
    sw_nxt_TRIGGER_IP_PENDING[0][32];
 nxt_TRIGGER_IP_PENDING[0][33] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[33] :
    sw_nxt_TRIGGER_IP_PENDING[0][33];
 nxt_TRIGGER_IP_PENDING[0][34] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[34] :
    sw_nxt_TRIGGER_IP_PENDING[0][34];
 nxt_TRIGGER_IP_PENDING[0][35] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[35] :
    sw_nxt_TRIGGER_IP_PENDING[0][35];
 nxt_TRIGGER_IP_PENDING[0][36] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[36] :
    sw_nxt_TRIGGER_IP_PENDING[0][36];
 nxt_TRIGGER_IP_PENDING[0][37] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[37] :
    sw_nxt_TRIGGER_IP_PENDING[0][37];
 nxt_TRIGGER_IP_PENDING[0][38] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[38] :
    sw_nxt_TRIGGER_IP_PENDING[0][38];
 nxt_TRIGGER_IP_PENDING[0][39] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[39] :
    sw_nxt_TRIGGER_IP_PENDING[0][39];
 nxt_TRIGGER_IP_PENDING[0][40] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[40] :
    sw_nxt_TRIGGER_IP_PENDING[0][40];
 nxt_TRIGGER_IP_PENDING[0][41] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[41] :
    sw_nxt_TRIGGER_IP_PENDING[0][41];
 nxt_TRIGGER_IP_PENDING[0][42] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[42] :
    sw_nxt_TRIGGER_IP_PENDING[0][42];
 nxt_TRIGGER_IP_PENDING[0][43] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[43] :
    sw_nxt_TRIGGER_IP_PENDING[0][43];
 nxt_TRIGGER_IP_PENDING[0][44] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[44] :
    sw_nxt_TRIGGER_IP_PENDING[0][44];
 nxt_TRIGGER_IP_PENDING[0][45] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[45] :
    sw_nxt_TRIGGER_IP_PENDING[0][45];
 nxt_TRIGGER_IP_PENDING[0][46] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[46] :
    sw_nxt_TRIGGER_IP_PENDING[0][46];
 nxt_TRIGGER_IP_PENDING[0][47] = 
    load_TRIGGER_IP[0].PENDING ?
    new_TRIGGER_IP[0].PENDING[47] :
    sw_nxt_TRIGGER_IP_PENDING[0][47];
 nxt_TRIGGER_IP_PENDING[1][0] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[0] :
    sw_nxt_TRIGGER_IP_PENDING[1][0];
 nxt_TRIGGER_IP_PENDING[1][1] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[1] :
    sw_nxt_TRIGGER_IP_PENDING[1][1];
 nxt_TRIGGER_IP_PENDING[1][2] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[2] :
    sw_nxt_TRIGGER_IP_PENDING[1][2];
 nxt_TRIGGER_IP_PENDING[1][3] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[3] :
    sw_nxt_TRIGGER_IP_PENDING[1][3];
 nxt_TRIGGER_IP_PENDING[1][4] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[4] :
    sw_nxt_TRIGGER_IP_PENDING[1][4];
 nxt_TRIGGER_IP_PENDING[1][5] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[5] :
    sw_nxt_TRIGGER_IP_PENDING[1][5];
 nxt_TRIGGER_IP_PENDING[1][6] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[6] :
    sw_nxt_TRIGGER_IP_PENDING[1][6];
 nxt_TRIGGER_IP_PENDING[1][7] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[7] :
    sw_nxt_TRIGGER_IP_PENDING[1][7];
 nxt_TRIGGER_IP_PENDING[1][8] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[8] :
    sw_nxt_TRIGGER_IP_PENDING[1][8];
 nxt_TRIGGER_IP_PENDING[1][9] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[9] :
    sw_nxt_TRIGGER_IP_PENDING[1][9];
 nxt_TRIGGER_IP_PENDING[1][10] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[10] :
    sw_nxt_TRIGGER_IP_PENDING[1][10];
 nxt_TRIGGER_IP_PENDING[1][11] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[11] :
    sw_nxt_TRIGGER_IP_PENDING[1][11];
 nxt_TRIGGER_IP_PENDING[1][12] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[12] :
    sw_nxt_TRIGGER_IP_PENDING[1][12];
 nxt_TRIGGER_IP_PENDING[1][13] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[13] :
    sw_nxt_TRIGGER_IP_PENDING[1][13];
 nxt_TRIGGER_IP_PENDING[1][14] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[14] :
    sw_nxt_TRIGGER_IP_PENDING[1][14];
 nxt_TRIGGER_IP_PENDING[1][15] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[15] :
    sw_nxt_TRIGGER_IP_PENDING[1][15];
 nxt_TRIGGER_IP_PENDING[1][16] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[16] :
    sw_nxt_TRIGGER_IP_PENDING[1][16];
 nxt_TRIGGER_IP_PENDING[1][17] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[17] :
    sw_nxt_TRIGGER_IP_PENDING[1][17];
 nxt_TRIGGER_IP_PENDING[1][18] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[18] :
    sw_nxt_TRIGGER_IP_PENDING[1][18];
 nxt_TRIGGER_IP_PENDING[1][19] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[19] :
    sw_nxt_TRIGGER_IP_PENDING[1][19];
 nxt_TRIGGER_IP_PENDING[1][20] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[20] :
    sw_nxt_TRIGGER_IP_PENDING[1][20];
 nxt_TRIGGER_IP_PENDING[1][21] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[21] :
    sw_nxt_TRIGGER_IP_PENDING[1][21];
 nxt_TRIGGER_IP_PENDING[1][22] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[22] :
    sw_nxt_TRIGGER_IP_PENDING[1][22];
 nxt_TRIGGER_IP_PENDING[1][23] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[23] :
    sw_nxt_TRIGGER_IP_PENDING[1][23];
 nxt_TRIGGER_IP_PENDING[1][24] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[24] :
    sw_nxt_TRIGGER_IP_PENDING[1][24];
 nxt_TRIGGER_IP_PENDING[1][25] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[25] :
    sw_nxt_TRIGGER_IP_PENDING[1][25];
 nxt_TRIGGER_IP_PENDING[1][26] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[26] :
    sw_nxt_TRIGGER_IP_PENDING[1][26];
 nxt_TRIGGER_IP_PENDING[1][27] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[27] :
    sw_nxt_TRIGGER_IP_PENDING[1][27];
 nxt_TRIGGER_IP_PENDING[1][28] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[28] :
    sw_nxt_TRIGGER_IP_PENDING[1][28];
 nxt_TRIGGER_IP_PENDING[1][29] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[29] :
    sw_nxt_TRIGGER_IP_PENDING[1][29];
 nxt_TRIGGER_IP_PENDING[1][30] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[30] :
    sw_nxt_TRIGGER_IP_PENDING[1][30];
 nxt_TRIGGER_IP_PENDING[1][31] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[31] :
    sw_nxt_TRIGGER_IP_PENDING[1][31];
 nxt_TRIGGER_IP_PENDING[1][32] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[32] :
    sw_nxt_TRIGGER_IP_PENDING[1][32];
 nxt_TRIGGER_IP_PENDING[1][33] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[33] :
    sw_nxt_TRIGGER_IP_PENDING[1][33];
 nxt_TRIGGER_IP_PENDING[1][34] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[34] :
    sw_nxt_TRIGGER_IP_PENDING[1][34];
 nxt_TRIGGER_IP_PENDING[1][35] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[35] :
    sw_nxt_TRIGGER_IP_PENDING[1][35];
 nxt_TRIGGER_IP_PENDING[1][36] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[36] :
    sw_nxt_TRIGGER_IP_PENDING[1][36];
 nxt_TRIGGER_IP_PENDING[1][37] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[37] :
    sw_nxt_TRIGGER_IP_PENDING[1][37];
 nxt_TRIGGER_IP_PENDING[1][38] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[38] :
    sw_nxt_TRIGGER_IP_PENDING[1][38];
 nxt_TRIGGER_IP_PENDING[1][39] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[39] :
    sw_nxt_TRIGGER_IP_PENDING[1][39];
 nxt_TRIGGER_IP_PENDING[1][40] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[40] :
    sw_nxt_TRIGGER_IP_PENDING[1][40];
 nxt_TRIGGER_IP_PENDING[1][41] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[41] :
    sw_nxt_TRIGGER_IP_PENDING[1][41];
 nxt_TRIGGER_IP_PENDING[1][42] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[42] :
    sw_nxt_TRIGGER_IP_PENDING[1][42];
 nxt_TRIGGER_IP_PENDING[1][43] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[43] :
    sw_nxt_TRIGGER_IP_PENDING[1][43];
 nxt_TRIGGER_IP_PENDING[1][44] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[44] :
    sw_nxt_TRIGGER_IP_PENDING[1][44];
 nxt_TRIGGER_IP_PENDING[1][45] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[45] :
    sw_nxt_TRIGGER_IP_PENDING[1][45];
 nxt_TRIGGER_IP_PENDING[1][46] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[46] :
    sw_nxt_TRIGGER_IP_PENDING[1][46];
 nxt_TRIGGER_IP_PENDING[1][47] = 
    load_TRIGGER_IP[1].PENDING ?
    new_TRIGGER_IP[1].PENDING[47] :
    sw_nxt_TRIGGER_IP_PENDING[1][47];
end



`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][0], nxt_TRIGGER_IP_PENDING[0][0], TRIGGER_IP[0].PENDING[0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][1], nxt_TRIGGER_IP_PENDING[0][1], TRIGGER_IP[0].PENDING[1])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][2], nxt_TRIGGER_IP_PENDING[0][2], TRIGGER_IP[0].PENDING[2])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][3], nxt_TRIGGER_IP_PENDING[0][3], TRIGGER_IP[0].PENDING[3])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][4], nxt_TRIGGER_IP_PENDING[0][4], TRIGGER_IP[0].PENDING[4])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][5], nxt_TRIGGER_IP_PENDING[0][5], TRIGGER_IP[0].PENDING[5])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][6], nxt_TRIGGER_IP_PENDING[0][6], TRIGGER_IP[0].PENDING[6])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][7], nxt_TRIGGER_IP_PENDING[0][7], TRIGGER_IP[0].PENDING[7])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][8], nxt_TRIGGER_IP_PENDING[0][8], TRIGGER_IP[0].PENDING[8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][9], nxt_TRIGGER_IP_PENDING[0][9], TRIGGER_IP[0].PENDING[9])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][10], nxt_TRIGGER_IP_PENDING[0][10], TRIGGER_IP[0].PENDING[10])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][11], nxt_TRIGGER_IP_PENDING[0][11], TRIGGER_IP[0].PENDING[11])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][12], nxt_TRIGGER_IP_PENDING[0][12], TRIGGER_IP[0].PENDING[12])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][13], nxt_TRIGGER_IP_PENDING[0][13], TRIGGER_IP[0].PENDING[13])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][14], nxt_TRIGGER_IP_PENDING[0][14], TRIGGER_IP[0].PENDING[14])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][15], nxt_TRIGGER_IP_PENDING[0][15], TRIGGER_IP[0].PENDING[15])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][16], nxt_TRIGGER_IP_PENDING[0][16], TRIGGER_IP[0].PENDING[16])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][17], nxt_TRIGGER_IP_PENDING[0][17], TRIGGER_IP[0].PENDING[17])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][18], nxt_TRIGGER_IP_PENDING[0][18], TRIGGER_IP[0].PENDING[18])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][19], nxt_TRIGGER_IP_PENDING[0][19], TRIGGER_IP[0].PENDING[19])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][20], nxt_TRIGGER_IP_PENDING[0][20], TRIGGER_IP[0].PENDING[20])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][21], nxt_TRIGGER_IP_PENDING[0][21], TRIGGER_IP[0].PENDING[21])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][22], nxt_TRIGGER_IP_PENDING[0][22], TRIGGER_IP[0].PENDING[22])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][23], nxt_TRIGGER_IP_PENDING[0][23], TRIGGER_IP[0].PENDING[23])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][24], nxt_TRIGGER_IP_PENDING[0][24], TRIGGER_IP[0].PENDING[24])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][25], nxt_TRIGGER_IP_PENDING[0][25], TRIGGER_IP[0].PENDING[25])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][26], nxt_TRIGGER_IP_PENDING[0][26], TRIGGER_IP[0].PENDING[26])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][27], nxt_TRIGGER_IP_PENDING[0][27], TRIGGER_IP[0].PENDING[27])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][28], nxt_TRIGGER_IP_PENDING[0][28], TRIGGER_IP[0].PENDING[28])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][29], nxt_TRIGGER_IP_PENDING[0][29], TRIGGER_IP[0].PENDING[29])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][30], nxt_TRIGGER_IP_PENDING[0][30], TRIGGER_IP[0].PENDING[30])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][31], nxt_TRIGGER_IP_PENDING[0][31], TRIGGER_IP[0].PENDING[31])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][32], nxt_TRIGGER_IP_PENDING[0][32], TRIGGER_IP[0].PENDING[32])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][33], nxt_TRIGGER_IP_PENDING[0][33], TRIGGER_IP[0].PENDING[33])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][34], nxt_TRIGGER_IP_PENDING[0][34], TRIGGER_IP[0].PENDING[34])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][35], nxt_TRIGGER_IP_PENDING[0][35], TRIGGER_IP[0].PENDING[35])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][36], nxt_TRIGGER_IP_PENDING[0][36], TRIGGER_IP[0].PENDING[36])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][37], nxt_TRIGGER_IP_PENDING[0][37], TRIGGER_IP[0].PENDING[37])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][38], nxt_TRIGGER_IP_PENDING[0][38], TRIGGER_IP[0].PENDING[38])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][39], nxt_TRIGGER_IP_PENDING[0][39], TRIGGER_IP[0].PENDING[39])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][40], nxt_TRIGGER_IP_PENDING[0][40], TRIGGER_IP[0].PENDING[40])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][41], nxt_TRIGGER_IP_PENDING[0][41], TRIGGER_IP[0].PENDING[41])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][42], nxt_TRIGGER_IP_PENDING[0][42], TRIGGER_IP[0].PENDING[42])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][43], nxt_TRIGGER_IP_PENDING[0][43], TRIGGER_IP[0].PENDING[43])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][44], nxt_TRIGGER_IP_PENDING[0][44], TRIGGER_IP[0].PENDING[44])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][45], nxt_TRIGGER_IP_PENDING[0][45], TRIGGER_IP[0].PENDING[45])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][46], nxt_TRIGGER_IP_PENDING[0][46], TRIGGER_IP[0].PENDING[46])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[0][47], nxt_TRIGGER_IP_PENDING[0][47], TRIGGER_IP[0].PENDING[47])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][0], nxt_TRIGGER_IP_PENDING[1][0], TRIGGER_IP[1].PENDING[0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][1], nxt_TRIGGER_IP_PENDING[1][1], TRIGGER_IP[1].PENDING[1])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][2], nxt_TRIGGER_IP_PENDING[1][2], TRIGGER_IP[1].PENDING[2])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][3], nxt_TRIGGER_IP_PENDING[1][3], TRIGGER_IP[1].PENDING[3])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][4], nxt_TRIGGER_IP_PENDING[1][4], TRIGGER_IP[1].PENDING[4])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][5], nxt_TRIGGER_IP_PENDING[1][5], TRIGGER_IP[1].PENDING[5])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][6], nxt_TRIGGER_IP_PENDING[1][6], TRIGGER_IP[1].PENDING[6])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][7], nxt_TRIGGER_IP_PENDING[1][7], TRIGGER_IP[1].PENDING[7])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][8], nxt_TRIGGER_IP_PENDING[1][8], TRIGGER_IP[1].PENDING[8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][9], nxt_TRIGGER_IP_PENDING[1][9], TRIGGER_IP[1].PENDING[9])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][10], nxt_TRIGGER_IP_PENDING[1][10], TRIGGER_IP[1].PENDING[10])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][11], nxt_TRIGGER_IP_PENDING[1][11], TRIGGER_IP[1].PENDING[11])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][12], nxt_TRIGGER_IP_PENDING[1][12], TRIGGER_IP[1].PENDING[12])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][13], nxt_TRIGGER_IP_PENDING[1][13], TRIGGER_IP[1].PENDING[13])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][14], nxt_TRIGGER_IP_PENDING[1][14], TRIGGER_IP[1].PENDING[14])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][15], nxt_TRIGGER_IP_PENDING[1][15], TRIGGER_IP[1].PENDING[15])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][16], nxt_TRIGGER_IP_PENDING[1][16], TRIGGER_IP[1].PENDING[16])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][17], nxt_TRIGGER_IP_PENDING[1][17], TRIGGER_IP[1].PENDING[17])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][18], nxt_TRIGGER_IP_PENDING[1][18], TRIGGER_IP[1].PENDING[18])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][19], nxt_TRIGGER_IP_PENDING[1][19], TRIGGER_IP[1].PENDING[19])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][20], nxt_TRIGGER_IP_PENDING[1][20], TRIGGER_IP[1].PENDING[20])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][21], nxt_TRIGGER_IP_PENDING[1][21], TRIGGER_IP[1].PENDING[21])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][22], nxt_TRIGGER_IP_PENDING[1][22], TRIGGER_IP[1].PENDING[22])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][23], nxt_TRIGGER_IP_PENDING[1][23], TRIGGER_IP[1].PENDING[23])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][24], nxt_TRIGGER_IP_PENDING[1][24], TRIGGER_IP[1].PENDING[24])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][25], nxt_TRIGGER_IP_PENDING[1][25], TRIGGER_IP[1].PENDING[25])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][26], nxt_TRIGGER_IP_PENDING[1][26], TRIGGER_IP[1].PENDING[26])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][27], nxt_TRIGGER_IP_PENDING[1][27], TRIGGER_IP[1].PENDING[27])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][28], nxt_TRIGGER_IP_PENDING[1][28], TRIGGER_IP[1].PENDING[28])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][29], nxt_TRIGGER_IP_PENDING[1][29], TRIGGER_IP[1].PENDING[29])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][30], nxt_TRIGGER_IP_PENDING[1][30], TRIGGER_IP[1].PENDING[30])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][31], nxt_TRIGGER_IP_PENDING[1][31], TRIGGER_IP[1].PENDING[31])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][32], nxt_TRIGGER_IP_PENDING[1][32], TRIGGER_IP[1].PENDING[32])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][33], nxt_TRIGGER_IP_PENDING[1][33], TRIGGER_IP[1].PENDING[33])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][34], nxt_TRIGGER_IP_PENDING[1][34], TRIGGER_IP[1].PENDING[34])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][35], nxt_TRIGGER_IP_PENDING[1][35], TRIGGER_IP[1].PENDING[35])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][36], nxt_TRIGGER_IP_PENDING[1][36], TRIGGER_IP[1].PENDING[36])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][37], nxt_TRIGGER_IP_PENDING[1][37], TRIGGER_IP[1].PENDING[37])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][38], nxt_TRIGGER_IP_PENDING[1][38], TRIGGER_IP[1].PENDING[38])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][39], nxt_TRIGGER_IP_PENDING[1][39], TRIGGER_IP[1].PENDING[39])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][40], nxt_TRIGGER_IP_PENDING[1][40], TRIGGER_IP[1].PENDING[40])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][41], nxt_TRIGGER_IP_PENDING[1][41], TRIGGER_IP[1].PENDING[41])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][42], nxt_TRIGGER_IP_PENDING[1][42], TRIGGER_IP[1].PENDING[42])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][43], nxt_TRIGGER_IP_PENDING[1][43], TRIGGER_IP[1].PENDING[43])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][44], nxt_TRIGGER_IP_PENDING[1][44], TRIGGER_IP[1].PENDING[44])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][45], nxt_TRIGGER_IP_PENDING[1][45], TRIGGER_IP[1].PENDING[45])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][46], nxt_TRIGGER_IP_PENDING[1][46], TRIGGER_IP[1].PENDING[46])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_TRIGGER_IP_PENDING[1][47], nxt_TRIGGER_IP_PENDING[1][47], TRIGGER_IP[1].PENDING[47])

//---------------------------------------------------------------------
// TRIGGER_IM Address Decode
logic [1:0] addr_decode_TRIGGER_IM;
logic [1:0] write_req_TRIGGER_IM;
always_comb begin
   addr_decode_TRIGGER_IM[0] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == TRIGGER_IM_DECODE_ADDR[0]) && req.valid ;
   addr_decode_TRIGGER_IM[1] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == TRIGGER_IM_DECODE_ADDR[1]) && req.valid ;
   write_req_TRIGGER_IM[0] = IsMEMWr && addr_decode_TRIGGER_IM[0] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_TRIGGER_IM[1] = IsMEMWr && addr_decode_TRIGGER_IM[1] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
end

// ----------------------------------------------------------------------
// TRIGGER_IM.MASK x8 RW, using RW template.
logic [1:0][5:0] up_TRIGGER_IM_MASK;
always_comb begin
 up_TRIGGER_IM_MASK[0] =
    ({6{write_req_TRIGGER_IM[0] }} &
    be[5:0]);
 up_TRIGGER_IM_MASK[1] =
    ({6{write_req_TRIGGER_IM[1] }} &
    be[5:0]);
end

logic [1:0][47:0] nxt_TRIGGER_IM_MASK;
always_comb begin
 nxt_TRIGGER_IM_MASK[0] = write_data[47:0];

 nxt_TRIGGER_IM_MASK[1] = write_data[47:0];

end


`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[0][0], nxt_TRIGGER_IM_MASK[0][7:0], TRIGGER_IM[0].MASK[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[0][1], nxt_TRIGGER_IM_MASK[0][15:8], TRIGGER_IM[0].MASK[15:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[0][2], nxt_TRIGGER_IM_MASK[0][23:16], TRIGGER_IM[0].MASK[23:16])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[0][3], nxt_TRIGGER_IM_MASK[0][31:24], TRIGGER_IM[0].MASK[31:24])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[0][4], nxt_TRIGGER_IM_MASK[0][39:32], TRIGGER_IM[0].MASK[39:32])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[0][5], nxt_TRIGGER_IM_MASK[0][47:40], TRIGGER_IM[0].MASK[47:40])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[1][0], nxt_TRIGGER_IM_MASK[1][7:0], TRIGGER_IM[1].MASK[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[1][1], nxt_TRIGGER_IM_MASK[1][15:8], TRIGGER_IM[1].MASK[15:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[1][2], nxt_TRIGGER_IM_MASK[1][23:16], TRIGGER_IM[1].MASK[23:16])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[1][3], nxt_TRIGGER_IM_MASK[1][31:24], TRIGGER_IM[1].MASK[31:24])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[1][4], nxt_TRIGGER_IM_MASK[1][39:32], TRIGGER_IM[1].MASK[39:32])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'hFF, up_TRIGGER_IM_MASK[1][5], nxt_TRIGGER_IM_MASK[1][47:40], TRIGGER_IM[1].MASK[47:40])

//---------------------------------------------------------------------
// TRIGGER_RATE_LIM_EMPTY Address Decode
// ----------------------------------------------------------------------
// TRIGGER_RATE_LIM_EMPTY.EMPTY x8 RO/V, using RO/V template.
assign TRIGGER_RATE_LIM_EMPTY.EMPTY = new_TRIGGER_RATE_LIM_EMPTY.EMPTY;




// ----------------------------------------------------------------------
// MA_TCN_FIFO_0 using HANDCODED_REG template.
logic addr_decode_MA_TCN_FIFO_0;
logic write_req_MA_TCN_FIFO_0;
logic read_req_MA_TCN_FIFO_0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h1?,1'b?},
      {40'b1?,4'h?,1'b?},
      {40'b1??,4'h?,1'b?},
      {40'b1???,4'h?,1'b?},
      {44'h10?,1'b?}:
          addr_decode_MA_TCN_FIFO_0 = req.valid;
      default: 
         addr_decode_MA_TCN_FIFO_0 = 1'b0; 
   endcase
end

always_comb write_req_MA_TCN_FIFO_0 = f_IsMEMWr(req_opcode) && addr_decode_MA_TCN_FIFO_0 ;
always_comb read_req_MA_TCN_FIFO_0  = f_IsMEMRd(req_opcode) && addr_decode_MA_TCN_FIFO_0 ;

always_comb we_MA_TCN_FIFO_0 = {8{write_req_MA_TCN_FIFO_0}} & be;
always_comb re_MA_TCN_FIFO_0 = {8{read_req_MA_TCN_FIFO_0}} & be;
always_comb handcode_reg_wdata_MA_TCN_FIFO_0 = write_data;


// ----------------------------------------------------------------------
// MA_TCN_FIFO_1 using HANDCODED_REG template.
logic addr_decode_MA_TCN_FIFO_1;
logic write_req_MA_TCN_FIFO_1;
logic read_req_MA_TCN_FIFO_1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h11?,1'b?},
      {36'h1,4'b001?,4'h?,1'b?},
      {36'h1,4'b01??,4'h?,1'b?},
      {36'h1,4'b1???,4'h?,1'b?},
      {44'h20?,1'b?}:
          addr_decode_MA_TCN_FIFO_1 = req.valid;
      default: 
         addr_decode_MA_TCN_FIFO_1 = 1'b0; 
   endcase
end

always_comb write_req_MA_TCN_FIFO_1 = f_IsMEMWr(req_opcode) && addr_decode_MA_TCN_FIFO_1 ;
always_comb read_req_MA_TCN_FIFO_1  = f_IsMEMRd(req_opcode) && addr_decode_MA_TCN_FIFO_1 ;

always_comb we_MA_TCN_FIFO_1 = {8{write_req_MA_TCN_FIFO_1}} & be;
always_comb re_MA_TCN_FIFO_1 = {8{read_req_MA_TCN_FIFO_1}} & be;
always_comb handcode_reg_wdata_MA_TCN_FIFO_1 = write_data;


// ----------------------------------------------------------------------
// MA_TCN_DEQUEUE using HANDCODED_REG template.
logic addr_decode_MA_TCN_DEQUEUE;
logic write_req_MA_TCN_DEQUEUE;
logic read_req_MA_TCN_DEQUEUE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h210,1'b0}: 
         addr_decode_MA_TCN_DEQUEUE = req.valid;
      default: 
         addr_decode_MA_TCN_DEQUEUE = 1'b0; 
   endcase
end

always_comb write_req_MA_TCN_DEQUEUE = f_IsMEMWr(req_opcode) && addr_decode_MA_TCN_DEQUEUE ;
always_comb read_req_MA_TCN_DEQUEUE  = f_IsMEMRd(req_opcode) && addr_decode_MA_TCN_DEQUEUE ;

always_comb we_MA_TCN_DEQUEUE = {8{write_req_MA_TCN_DEQUEUE}} & be;
always_comb re_MA_TCN_DEQUEUE = {8{read_req_MA_TCN_DEQUEUE}} & be;
always_comb handcode_reg_wdata_MA_TCN_DEQUEUE = write_data;


// ----------------------------------------------------------------------
// MA_TCN_DATA_0 using HANDCODED_REG template.
logic addr_decode_MA_TCN_DATA_0;
logic write_req_MA_TCN_DATA_0;
logic read_req_MA_TCN_DATA_0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h210,1'b1}: 
         addr_decode_MA_TCN_DATA_0 = req.valid;
      default: 
         addr_decode_MA_TCN_DATA_0 = 1'b0; 
   endcase
end

always_comb write_req_MA_TCN_DATA_0 = f_IsMEMWr(req_opcode) && addr_decode_MA_TCN_DATA_0 ;
always_comb read_req_MA_TCN_DATA_0  = f_IsMEMRd(req_opcode) && addr_decode_MA_TCN_DATA_0 ;

always_comb we_MA_TCN_DATA_0 = {8{write_req_MA_TCN_DATA_0}} & be;
always_comb re_MA_TCN_DATA_0 = {8{read_req_MA_TCN_DATA_0}} & be;
always_comb handcode_reg_wdata_MA_TCN_DATA_0 = write_data;


// ----------------------------------------------------------------------
// MA_TCN_DATA_1 using HANDCODED_REG template.
logic addr_decode_MA_TCN_DATA_1;
logic write_req_MA_TCN_DATA_1;
logic read_req_MA_TCN_DATA_1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h211,1'b0}: 
         addr_decode_MA_TCN_DATA_1 = req.valid;
      default: 
         addr_decode_MA_TCN_DATA_1 = 1'b0; 
   endcase
end

always_comb write_req_MA_TCN_DATA_1 = f_IsMEMWr(req_opcode) && addr_decode_MA_TCN_DATA_1 ;
always_comb read_req_MA_TCN_DATA_1  = f_IsMEMRd(req_opcode) && addr_decode_MA_TCN_DATA_1 ;

always_comb we_MA_TCN_DATA_1 = {8{write_req_MA_TCN_DATA_1}} & be;
always_comb re_MA_TCN_DATA_1 = {8{read_req_MA_TCN_DATA_1}} & be;
always_comb handcode_reg_wdata_MA_TCN_DATA_1 = write_data;


// ----------------------------------------------------------------------
// MA_TCN_PTR_HEAD using HANDCODED_REG template.
logic addr_decode_MA_TCN_PTR_HEAD;
logic write_req_MA_TCN_PTR_HEAD;
logic read_req_MA_TCN_PTR_HEAD;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h211,1'b1}: 
         addr_decode_MA_TCN_PTR_HEAD = req.valid;
      default: 
         addr_decode_MA_TCN_PTR_HEAD = 1'b0; 
   endcase
end

always_comb write_req_MA_TCN_PTR_HEAD = f_IsMEMWr(req_opcode) && addr_decode_MA_TCN_PTR_HEAD ;
always_comb read_req_MA_TCN_PTR_HEAD  = f_IsMEMRd(req_opcode) && addr_decode_MA_TCN_PTR_HEAD ;

always_comb we_MA_TCN_PTR_HEAD = {8{write_req_MA_TCN_PTR_HEAD}} & be;
always_comb re_MA_TCN_PTR_HEAD = {8{read_req_MA_TCN_PTR_HEAD}} & be;
always_comb handcode_reg_wdata_MA_TCN_PTR_HEAD = write_data;


// ----------------------------------------------------------------------
// MA_TCN_PTR_TAIL using HANDCODED_REG template.
logic addr_decode_MA_TCN_PTR_TAIL;
logic write_req_MA_TCN_PTR_TAIL;
logic read_req_MA_TCN_PTR_TAIL;

always_comb begin 
   unique casez (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h212,1'b0}: 
         addr_decode_MA_TCN_PTR_TAIL = req.valid;
      default: 
         addr_decode_MA_TCN_PTR_TAIL = 1'b0; 
   endcase
end

always_comb write_req_MA_TCN_PTR_TAIL = f_IsMEMWr(req_opcode) && addr_decode_MA_TCN_PTR_TAIL ;
always_comb read_req_MA_TCN_PTR_TAIL  = f_IsMEMRd(req_opcode) && addr_decode_MA_TCN_PTR_TAIL ;

always_comb we_MA_TCN_PTR_TAIL = {8{write_req_MA_TCN_PTR_TAIL}} & be;
always_comb re_MA_TCN_PTR_TAIL = {8{read_req_MA_TCN_PTR_TAIL}} & be;
always_comb handcode_reg_wdata_MA_TCN_PTR_TAIL = write_data;


//---------------------------------------------------------------------
// MA_TCN_IP Address Decode
logic  addr_decode_MA_TCN_IP;
logic  write_req_MA_TCN_IP;
always_comb begin
   addr_decode_MA_TCN_IP = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_IP_DECODE_ADDR) && req.valid ;
   write_req_MA_TCN_IP = IsMEMWr && addr_decode_MA_TCN_IP && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
end

// ----------------------------------------------------------------------
// MA_TCN_IP.TCN_OVERFLOW x1 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [0:0] req_up_MA_TCN_IP_TCN_OVERFLOW;
always_comb begin
 req_up_MA_TCN_IP_TCN_OVERFLOW[0:0] = 
   {1{write_req_MA_TCN_IP & be[0]}}
;
end

logic [0:0] clr_MA_TCN_IP_TCN_OVERFLOW;
always_comb begin
 clr_MA_TCN_IP_TCN_OVERFLOW = write_data[0:0] & req_up_MA_TCN_IP_TCN_OVERFLOW;

end
logic [0:0] swwr_MA_TCN_IP_TCN_OVERFLOW;
logic [0:0] sw_nxt_MA_TCN_IP_TCN_OVERFLOW;
always_comb begin
 swwr_MA_TCN_IP_TCN_OVERFLOW = clr_MA_TCN_IP_TCN_OVERFLOW;
 sw_nxt_MA_TCN_IP_TCN_OVERFLOW = {1{1'b0}};

end
logic [0:0] up_MA_TCN_IP_TCN_OVERFLOW;
logic [0:0] nxt_MA_TCN_IP_TCN_OVERFLOW;
always_comb begin
 up_MA_TCN_IP_TCN_OVERFLOW = 
   swwr_MA_TCN_IP_TCN_OVERFLOW | {1{load_MA_TCN_IP.TCN_OVERFLOW}};
end
always_comb begin
 nxt_MA_TCN_IP_TCN_OVERFLOW[0] = 
    load_MA_TCN_IP.TCN_OVERFLOW ?
    new_MA_TCN_IP.TCN_OVERFLOW[0] :
    sw_nxt_MA_TCN_IP_TCN_OVERFLOW[0];
end



`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_MA_TCN_IP_TCN_OVERFLOW[0], nxt_MA_TCN_IP_TCN_OVERFLOW[0], MA_TCN_IP.TCN_OVERFLOW[0])

// ----------------------------------------------------------------------
// MA_TCN_IP.PENDING_EVENTS x1 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [0:0] req_up_MA_TCN_IP_PENDING_EVENTS;
always_comb begin
 req_up_MA_TCN_IP_PENDING_EVENTS[0:0] = 
   {1{write_req_MA_TCN_IP & be[0]}}
;
end

logic [0:0] clr_MA_TCN_IP_PENDING_EVENTS;
always_comb begin
 clr_MA_TCN_IP_PENDING_EVENTS = write_data[1:1] & req_up_MA_TCN_IP_PENDING_EVENTS;

end
logic [0:0] swwr_MA_TCN_IP_PENDING_EVENTS;
logic [0:0] sw_nxt_MA_TCN_IP_PENDING_EVENTS;
always_comb begin
 swwr_MA_TCN_IP_PENDING_EVENTS = clr_MA_TCN_IP_PENDING_EVENTS;
 sw_nxt_MA_TCN_IP_PENDING_EVENTS = {1{1'b0}};

end
logic [0:0] up_MA_TCN_IP_PENDING_EVENTS;
logic [0:0] nxt_MA_TCN_IP_PENDING_EVENTS;
always_comb begin
 up_MA_TCN_IP_PENDING_EVENTS = 
   swwr_MA_TCN_IP_PENDING_EVENTS | {1{load_MA_TCN_IP.PENDING_EVENTS}};
end
always_comb begin
 nxt_MA_TCN_IP_PENDING_EVENTS[0] = 
    load_MA_TCN_IP.PENDING_EVENTS ?
    new_MA_TCN_IP.PENDING_EVENTS[0] :
    sw_nxt_MA_TCN_IP_PENDING_EVENTS[0];
end



`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_MA_TCN_IP_PENDING_EVENTS[0], nxt_MA_TCN_IP_PENDING_EVENTS[0], MA_TCN_IP.PENDING_EVENTS[0])

//---------------------------------------------------------------------
// MA_TCN_IM Address Decode
logic  addr_decode_MA_TCN_IM;
logic  write_req_MA_TCN_IM;
always_comb begin
   addr_decode_MA_TCN_IM = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_IM_DECODE_ADDR) && req.valid ;
   write_req_MA_TCN_IM = IsMEMWr && addr_decode_MA_TCN_IM && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
end

// ----------------------------------------------------------------------
// MA_TCN_IM.TCN_OVERFLOW x1 RW, using RW template.
logic [0:0] up_MA_TCN_IM_TCN_OVERFLOW;
always_comb begin
 up_MA_TCN_IM_TCN_OVERFLOW =
    ({1{write_req_MA_TCN_IM }} &
    be[0:0]);
end

logic [0:0] nxt_MA_TCN_IM_TCN_OVERFLOW;
always_comb begin
 nxt_MA_TCN_IM_TCN_OVERFLOW = write_data[0:0];

end


`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MA_TCN_IM_TCN_OVERFLOW[0], nxt_MA_TCN_IM_TCN_OVERFLOW[0:0], MA_TCN_IM.TCN_OVERFLOW[0:0])

// ----------------------------------------------------------------------
// MA_TCN_IM.PENDING_EVENTS x1 RW, using RW template.
logic [0:0] up_MA_TCN_IM_PENDING_EVENTS;
always_comb begin
 up_MA_TCN_IM_PENDING_EVENTS =
    ({1{write_req_MA_TCN_IM }} &
    be[0:0]);
end

logic [0:0] nxt_MA_TCN_IM_PENDING_EVENTS;
always_comb begin
 nxt_MA_TCN_IM_PENDING_EVENTS = write_data[1:1];

end


`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MA_TCN_IM_PENDING_EVENTS[0], nxt_MA_TCN_IM_PENDING_EVENTS[0:0], MA_TCN_IM.PENDING_EVENTS[0:0])

//---------------------------------------------------------------------
// MA_TCN_WM Address Decode
logic [16:0] addr_decode_MA_TCN_WM;
logic [16:0] write_req_MA_TCN_WM;
always_comb begin
   addr_decode_MA_TCN_WM[0] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[0]) && req.valid ;
   addr_decode_MA_TCN_WM[1] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[1]) && req.valid ;
   addr_decode_MA_TCN_WM[2] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[2]) && req.valid ;
   addr_decode_MA_TCN_WM[3] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[3]) && req.valid ;
   addr_decode_MA_TCN_WM[4] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[4]) && req.valid ;
   addr_decode_MA_TCN_WM[5] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[5]) && req.valid ;
   addr_decode_MA_TCN_WM[6] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[6]) && req.valid ;
   addr_decode_MA_TCN_WM[7] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[7]) && req.valid ;
   addr_decode_MA_TCN_WM[8] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[8]) && req.valid ;
   addr_decode_MA_TCN_WM[9] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[9]) && req.valid ;
   addr_decode_MA_TCN_WM[10] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[10]) && req.valid ;
   addr_decode_MA_TCN_WM[11] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[11]) && req.valid ;
   addr_decode_MA_TCN_WM[12] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[12]) && req.valid ;
   addr_decode_MA_TCN_WM[13] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[13]) && req.valid ;
   addr_decode_MA_TCN_WM[14] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[14]) && req.valid ;
   addr_decode_MA_TCN_WM[15] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[15]) && req.valid ;
   addr_decode_MA_TCN_WM[16] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_WM_DECODE_ADDR[16]) && req.valid ;
   write_req_MA_TCN_WM[0] = IsMEMWr && addr_decode_MA_TCN_WM[0] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[1] = IsMEMWr && addr_decode_MA_TCN_WM[1] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[2] = IsMEMWr && addr_decode_MA_TCN_WM[2] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[3] = IsMEMWr && addr_decode_MA_TCN_WM[3] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[4] = IsMEMWr && addr_decode_MA_TCN_WM[4] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[5] = IsMEMWr && addr_decode_MA_TCN_WM[5] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[6] = IsMEMWr && addr_decode_MA_TCN_WM[6] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[7] = IsMEMWr && addr_decode_MA_TCN_WM[7] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[8] = IsMEMWr && addr_decode_MA_TCN_WM[8] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[9] = IsMEMWr && addr_decode_MA_TCN_WM[9] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[10] = IsMEMWr && addr_decode_MA_TCN_WM[10] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[11] = IsMEMWr && addr_decode_MA_TCN_WM[11] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[12] = IsMEMWr && addr_decode_MA_TCN_WM[12] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[13] = IsMEMWr && addr_decode_MA_TCN_WM[13] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[14] = IsMEMWr && addr_decode_MA_TCN_WM[14] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[15] = IsMEMWr && addr_decode_MA_TCN_WM[15] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_WM[16] = IsMEMWr && addr_decode_MA_TCN_WM[16] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
end

// ----------------------------------------------------------------------
// MA_TCN_WM.WM x1 RW, using RW template.
logic [16:0][1:0] up_MA_TCN_WM_WM;
always_comb begin
 up_MA_TCN_WM_WM[0] =
    ({2{write_req_MA_TCN_WM[0] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[1] =
    ({2{write_req_MA_TCN_WM[1] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[2] =
    ({2{write_req_MA_TCN_WM[2] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[3] =
    ({2{write_req_MA_TCN_WM[3] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[4] =
    ({2{write_req_MA_TCN_WM[4] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[5] =
    ({2{write_req_MA_TCN_WM[5] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[6] =
    ({2{write_req_MA_TCN_WM[6] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[7] =
    ({2{write_req_MA_TCN_WM[7] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[8] =
    ({2{write_req_MA_TCN_WM[8] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[9] =
    ({2{write_req_MA_TCN_WM[9] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[10] =
    ({2{write_req_MA_TCN_WM[10] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[11] =
    ({2{write_req_MA_TCN_WM[11] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[12] =
    ({2{write_req_MA_TCN_WM[12] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[13] =
    ({2{write_req_MA_TCN_WM[13] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[14] =
    ({2{write_req_MA_TCN_WM[14] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[15] =
    ({2{write_req_MA_TCN_WM[15] }} &
    be[1:0]);
 up_MA_TCN_WM_WM[16] =
    ({2{write_req_MA_TCN_WM[16] }} &
    be[1:0]);
end

logic [16:0][8:0] nxt_MA_TCN_WM_WM;
always_comb begin
 nxt_MA_TCN_WM_WM[0] = write_data[8:0];

 nxt_MA_TCN_WM_WM[1] = write_data[8:0];

 nxt_MA_TCN_WM_WM[2] = write_data[8:0];

 nxt_MA_TCN_WM_WM[3] = write_data[8:0];

 nxt_MA_TCN_WM_WM[4] = write_data[8:0];

 nxt_MA_TCN_WM_WM[5] = write_data[8:0];

 nxt_MA_TCN_WM_WM[6] = write_data[8:0];

 nxt_MA_TCN_WM_WM[7] = write_data[8:0];

 nxt_MA_TCN_WM_WM[8] = write_data[8:0];

 nxt_MA_TCN_WM_WM[9] = write_data[8:0];

 nxt_MA_TCN_WM_WM[10] = write_data[8:0];

 nxt_MA_TCN_WM_WM[11] = write_data[8:0];

 nxt_MA_TCN_WM_WM[12] = write_data[8:0];

 nxt_MA_TCN_WM_WM[13] = write_data[8:0];

 nxt_MA_TCN_WM_WM[14] = write_data[8:0];

 nxt_MA_TCN_WM_WM[15] = write_data[8:0];

 nxt_MA_TCN_WM_WM[16] = write_data[8:0];

end


`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[0][0], nxt_MA_TCN_WM_WM[0][7:0], MA_TCN_WM[0].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[0][1], nxt_MA_TCN_WM_WM[0][8:8], MA_TCN_WM[0].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[1][0], nxt_MA_TCN_WM_WM[1][7:0], MA_TCN_WM[1].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[1][1], nxt_MA_TCN_WM_WM[1][8:8], MA_TCN_WM[1].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[2][0], nxt_MA_TCN_WM_WM[2][7:0], MA_TCN_WM[2].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[2][1], nxt_MA_TCN_WM_WM[2][8:8], MA_TCN_WM[2].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[3][0], nxt_MA_TCN_WM_WM[3][7:0], MA_TCN_WM[3].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[3][1], nxt_MA_TCN_WM_WM[3][8:8], MA_TCN_WM[3].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[4][0], nxt_MA_TCN_WM_WM[4][7:0], MA_TCN_WM[4].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[4][1], nxt_MA_TCN_WM_WM[4][8:8], MA_TCN_WM[4].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[5][0], nxt_MA_TCN_WM_WM[5][7:0], MA_TCN_WM[5].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[5][1], nxt_MA_TCN_WM_WM[5][8:8], MA_TCN_WM[5].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[6][0], nxt_MA_TCN_WM_WM[6][7:0], MA_TCN_WM[6].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[6][1], nxt_MA_TCN_WM_WM[6][8:8], MA_TCN_WM[6].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[7][0], nxt_MA_TCN_WM_WM[7][7:0], MA_TCN_WM[7].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[7][1], nxt_MA_TCN_WM_WM[7][8:8], MA_TCN_WM[7].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[8][0], nxt_MA_TCN_WM_WM[8][7:0], MA_TCN_WM[8].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[8][1], nxt_MA_TCN_WM_WM[8][8:8], MA_TCN_WM[8].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[9][0], nxt_MA_TCN_WM_WM[9][7:0], MA_TCN_WM[9].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[9][1], nxt_MA_TCN_WM_WM[9][8:8], MA_TCN_WM[9].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[10][0], nxt_MA_TCN_WM_WM[10][7:0], MA_TCN_WM[10].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[10][1], nxt_MA_TCN_WM_WM[10][8:8], MA_TCN_WM[10].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[11][0], nxt_MA_TCN_WM_WM[11][7:0], MA_TCN_WM[11].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[11][1], nxt_MA_TCN_WM_WM[11][8:8], MA_TCN_WM[11].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[12][0], nxt_MA_TCN_WM_WM[12][7:0], MA_TCN_WM[12].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[12][1], nxt_MA_TCN_WM_WM[12][8:8], MA_TCN_WM[12].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[13][0], nxt_MA_TCN_WM_WM[13][7:0], MA_TCN_WM[13].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[13][1], nxt_MA_TCN_WM_WM[13][8:8], MA_TCN_WM[13].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[14][0], nxt_MA_TCN_WM_WM[14][7:0], MA_TCN_WM[14].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[14][1], nxt_MA_TCN_WM_WM[14][8:8], MA_TCN_WM[14].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[15][0], nxt_MA_TCN_WM_WM[15][7:0], MA_TCN_WM[15].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[15][1], nxt_MA_TCN_WM_WM[15][8:8], MA_TCN_WM[15].WM[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h1E, up_MA_TCN_WM_WM[16][0], nxt_MA_TCN_WM_WM[16][7:0], MA_TCN_WM[16].WM[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_WM_WM[16][1], nxt_MA_TCN_WM_WM[16][8:8], MA_TCN_WM[16].WM[8:8])

//---------------------------------------------------------------------
// MA_TCN_USAGE Address Decode
logic [16:0] addr_decode_MA_TCN_USAGE;
logic [16:0] write_req_MA_TCN_USAGE;
always_comb begin
   addr_decode_MA_TCN_USAGE[0] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[0]) && req.valid ;
   addr_decode_MA_TCN_USAGE[1] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[1]) && req.valid ;
   addr_decode_MA_TCN_USAGE[2] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[2]) && req.valid ;
   addr_decode_MA_TCN_USAGE[3] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[3]) && req.valid ;
   addr_decode_MA_TCN_USAGE[4] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[4]) && req.valid ;
   addr_decode_MA_TCN_USAGE[5] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[5]) && req.valid ;
   addr_decode_MA_TCN_USAGE[6] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[6]) && req.valid ;
   addr_decode_MA_TCN_USAGE[7] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[7]) && req.valid ;
   addr_decode_MA_TCN_USAGE[8] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[8]) && req.valid ;
   addr_decode_MA_TCN_USAGE[9] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[9]) && req.valid ;
   addr_decode_MA_TCN_USAGE[10] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[10]) && req.valid ;
   addr_decode_MA_TCN_USAGE[11] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[11]) && req.valid ;
   addr_decode_MA_TCN_USAGE[12] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[12]) && req.valid ;
   addr_decode_MA_TCN_USAGE[13] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[13]) && req.valid ;
   addr_decode_MA_TCN_USAGE[14] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[14]) && req.valid ;
   addr_decode_MA_TCN_USAGE[15] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[15]) && req.valid ;
   addr_decode_MA_TCN_USAGE[16] = (req_addr[MBY_PPE_TRIG_APPLY_MISC_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MA_TCN_USAGE_DECODE_ADDR[16]) && req.valid ;
   write_req_MA_TCN_USAGE[0] = IsMEMWr && addr_decode_MA_TCN_USAGE[0] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[1] = IsMEMWr && addr_decode_MA_TCN_USAGE[1] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[2] = IsMEMWr && addr_decode_MA_TCN_USAGE[2] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[3] = IsMEMWr && addr_decode_MA_TCN_USAGE[3] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[4] = IsMEMWr && addr_decode_MA_TCN_USAGE[4] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[5] = IsMEMWr && addr_decode_MA_TCN_USAGE[5] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[6] = IsMEMWr && addr_decode_MA_TCN_USAGE[6] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[7] = IsMEMWr && addr_decode_MA_TCN_USAGE[7] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[8] = IsMEMWr && addr_decode_MA_TCN_USAGE[8] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[9] = IsMEMWr && addr_decode_MA_TCN_USAGE[9] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[10] = IsMEMWr && addr_decode_MA_TCN_USAGE[10] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[11] = IsMEMWr && addr_decode_MA_TCN_USAGE[11] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[12] = IsMEMWr && addr_decode_MA_TCN_USAGE[12] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[13] = IsMEMWr && addr_decode_MA_TCN_USAGE[13] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[14] = IsMEMWr && addr_decode_MA_TCN_USAGE[14] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[15] = IsMEMWr && addr_decode_MA_TCN_USAGE[15] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
   write_req_MA_TCN_USAGE[16] = IsMEMWr && addr_decode_MA_TCN_USAGE[16] && sb_fid_cond_trig_apply_misc && sb_bar_cond_trig_apply_misc;
end

// ----------------------------------------------------------------------
// MA_TCN_USAGE.USAGE x1 RW, using RW template.
logic [16:0][1:0] up_MA_TCN_USAGE_USAGE;
always_comb begin
 up_MA_TCN_USAGE_USAGE[0] =
    ({2{write_req_MA_TCN_USAGE[0] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[1] =
    ({2{write_req_MA_TCN_USAGE[1] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[2] =
    ({2{write_req_MA_TCN_USAGE[2] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[3] =
    ({2{write_req_MA_TCN_USAGE[3] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[4] =
    ({2{write_req_MA_TCN_USAGE[4] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[5] =
    ({2{write_req_MA_TCN_USAGE[5] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[6] =
    ({2{write_req_MA_TCN_USAGE[6] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[7] =
    ({2{write_req_MA_TCN_USAGE[7] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[8] =
    ({2{write_req_MA_TCN_USAGE[8] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[9] =
    ({2{write_req_MA_TCN_USAGE[9] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[10] =
    ({2{write_req_MA_TCN_USAGE[10] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[11] =
    ({2{write_req_MA_TCN_USAGE[11] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[12] =
    ({2{write_req_MA_TCN_USAGE[12] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[13] =
    ({2{write_req_MA_TCN_USAGE[13] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[14] =
    ({2{write_req_MA_TCN_USAGE[14] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[15] =
    ({2{write_req_MA_TCN_USAGE[15] }} &
    be[1:0]);
 up_MA_TCN_USAGE_USAGE[16] =
    ({2{write_req_MA_TCN_USAGE[16] }} &
    be[1:0]);
end

logic [16:0][8:0] nxt_MA_TCN_USAGE_USAGE;
always_comb begin
 nxt_MA_TCN_USAGE_USAGE[0] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[1] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[2] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[3] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[4] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[5] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[6] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[7] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[8] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[9] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[10] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[11] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[12] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[13] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[14] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[15] = write_data[8:0];

 nxt_MA_TCN_USAGE_USAGE[16] = write_data[8:0];

end


`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[0][0], nxt_MA_TCN_USAGE_USAGE[0][7:0], MA_TCN_USAGE[0].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[0][1], nxt_MA_TCN_USAGE_USAGE[0][8:8], MA_TCN_USAGE[0].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[1][0], nxt_MA_TCN_USAGE_USAGE[1][7:0], MA_TCN_USAGE[1].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[1][1], nxt_MA_TCN_USAGE_USAGE[1][8:8], MA_TCN_USAGE[1].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[2][0], nxt_MA_TCN_USAGE_USAGE[2][7:0], MA_TCN_USAGE[2].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[2][1], nxt_MA_TCN_USAGE_USAGE[2][8:8], MA_TCN_USAGE[2].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[3][0], nxt_MA_TCN_USAGE_USAGE[3][7:0], MA_TCN_USAGE[3].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[3][1], nxt_MA_TCN_USAGE_USAGE[3][8:8], MA_TCN_USAGE[3].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[4][0], nxt_MA_TCN_USAGE_USAGE[4][7:0], MA_TCN_USAGE[4].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[4][1], nxt_MA_TCN_USAGE_USAGE[4][8:8], MA_TCN_USAGE[4].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[5][0], nxt_MA_TCN_USAGE_USAGE[5][7:0], MA_TCN_USAGE[5].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[5][1], nxt_MA_TCN_USAGE_USAGE[5][8:8], MA_TCN_USAGE[5].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[6][0], nxt_MA_TCN_USAGE_USAGE[6][7:0], MA_TCN_USAGE[6].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[6][1], nxt_MA_TCN_USAGE_USAGE[6][8:8], MA_TCN_USAGE[6].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[7][0], nxt_MA_TCN_USAGE_USAGE[7][7:0], MA_TCN_USAGE[7].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[7][1], nxt_MA_TCN_USAGE_USAGE[7][8:8], MA_TCN_USAGE[7].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[8][0], nxt_MA_TCN_USAGE_USAGE[8][7:0], MA_TCN_USAGE[8].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[8][1], nxt_MA_TCN_USAGE_USAGE[8][8:8], MA_TCN_USAGE[8].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[9][0], nxt_MA_TCN_USAGE_USAGE[9][7:0], MA_TCN_USAGE[9].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[9][1], nxt_MA_TCN_USAGE_USAGE[9][8:8], MA_TCN_USAGE[9].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[10][0], nxt_MA_TCN_USAGE_USAGE[10][7:0], MA_TCN_USAGE[10].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[10][1], nxt_MA_TCN_USAGE_USAGE[10][8:8], MA_TCN_USAGE[10].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[11][0], nxt_MA_TCN_USAGE_USAGE[11][7:0], MA_TCN_USAGE[11].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[11][1], nxt_MA_TCN_USAGE_USAGE[11][8:8], MA_TCN_USAGE[11].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[12][0], nxt_MA_TCN_USAGE_USAGE[12][7:0], MA_TCN_USAGE[12].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[12][1], nxt_MA_TCN_USAGE_USAGE[12][8:8], MA_TCN_USAGE[12].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[13][0], nxt_MA_TCN_USAGE_USAGE[13][7:0], MA_TCN_USAGE[13].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[13][1], nxt_MA_TCN_USAGE_USAGE[13][8:8], MA_TCN_USAGE[13].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[14][0], nxt_MA_TCN_USAGE_USAGE[14][7:0], MA_TCN_USAGE[14].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[14][1], nxt_MA_TCN_USAGE_USAGE[14][8:8], MA_TCN_USAGE[14].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[15][0], nxt_MA_TCN_USAGE_USAGE[15][7:0], MA_TCN_USAGE[15].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[15][1], nxt_MA_TCN_USAGE_USAGE[15][8:8], MA_TCN_USAGE[15].USAGE[8:8])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 8'h0, up_MA_TCN_USAGE_USAGE[16][0], nxt_MA_TCN_USAGE_USAGE[16][7:0], MA_TCN_USAGE[16].USAGE[7:0])
`RTLGEN_MBY_PPE_TRIG_APPLY_MISC_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_MA_TCN_USAGE_USAGE[16][1], nxt_MA_TCN_USAGE_USAGE[16][8:8], MA_TCN_USAGE[16].USAGE[8:8])

// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_TRIG_APPLY_MISC_MAP_MEM) 
           {44'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_RATE_LIM_CFG_2;
                    ack.read_miss = handcode_error_TRIGGER_RATE_LIM_CFG_2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'b10??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_TRIGGER_ACTION_METADATA_MASK;
                    ack.read_miss = handcode_error_TRIGGER_ACTION_METADATA_MASK;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           TRIGGER_IP_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           TRIGGER_IP_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           TRIGGER_IM_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           TRIGGER_IM_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           TRIGGER_RATE_LIM_EMPTY_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h1?,1'b?},
           {40'b1?,4'h?,1'b?},
           {40'b1??,4'h?,1'b?},
           {40'b1???,4'h?,1'b?},
           {44'h10?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MA_TCN_FIFO_0;
                    ack.read_miss = handcode_error_MA_TCN_FIFO_0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h11?,1'b?},
           {36'h1,4'b001?,4'h?,1'b?},
           {36'h1,4'b01??,4'h?,1'b?},
           {36'h1,4'b1???,4'h?,1'b?},
           {44'h20?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MA_TCN_FIFO_1;
                    ack.read_miss = handcode_error_MA_TCN_FIFO_1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h210,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MA_TCN_DEQUEUE;
                    ack.read_miss = handcode_error_MA_TCN_DEQUEUE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h210,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MA_TCN_DATA_0;
                    ack.read_miss = handcode_error_MA_TCN_DATA_0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h211,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MA_TCN_DATA_1;
                    ack.read_miss = handcode_error_MA_TCN_DATA_1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h211,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MA_TCN_PTR_HEAD;
                    ack.read_miss = handcode_error_MA_TCN_PTR_HEAD;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h212,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MA_TCN_PTR_TAIL;
                    ack.read_miss = handcode_error_MA_TCN_PTR_TAIL;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_TRIG_APPLY_MISC_MAP_MEM) 
           {44'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_RATE_LIM_CFG_2;
                    ack.write_miss = handcode_error_TRIGGER_RATE_LIM_CFG_2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'b10??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_TRIGGER_ACTION_METADATA_MASK;
                    ack.write_miss = handcode_error_TRIGGER_ACTION_METADATA_MASK;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           TRIGGER_IP_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           TRIGGER_IP_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           TRIGGER_IM_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           TRIGGER_IM_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           TRIGGER_RATE_LIM_EMPTY_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h1?,1'b?},
           {40'b1?,4'h?,1'b?},
           {40'b1??,4'h?,1'b?},
           {40'b1???,4'h?,1'b?},
           {44'h10?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MA_TCN_FIFO_0;
                    ack.write_miss = handcode_error_MA_TCN_FIFO_0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h11?,1'b?},
           {36'h1,4'b001?,4'h?,1'b?},
           {36'h1,4'b01??,4'h?,1'b?},
           {36'h1,4'b1???,4'h?,1'b?},
           {44'h20?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MA_TCN_FIFO_1;
                    ack.write_miss = handcode_error_MA_TCN_FIFO_1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h210,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MA_TCN_DEQUEUE;
                    ack.write_miss = handcode_error_MA_TCN_DEQUEUE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h210,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MA_TCN_DATA_0;
                    ack.write_miss = handcode_error_MA_TCN_DATA_0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h211,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MA_TCN_DATA_1;
                    ack.write_miss = handcode_error_MA_TCN_DATA_1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h211,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MA_TCN_PTR_HEAD;
                    ack.write_miss = handcode_error_MA_TCN_PTR_HEAD;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h212,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MA_TCN_PTR_TAIL;
                    ack.write_miss = handcode_error_MA_TCN_PTR_TAIL;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_TRIG_APPLY_MISC_MAP_MEM) 
           {44'b0???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_RATE_LIM_CFG_2;
                 default: read_data = '0;
              endcase
           end
           {44'b10??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_TRIGGER_ACTION_METADATA_MASK;
                 default: read_data = '0;
              endcase
           end
           TRIGGER_IP_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {TRIGGER_IP[0]};
                 default: read_data = '0;
              endcase
           end
           TRIGGER_IP_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {TRIGGER_IP[1]};
                 default: read_data = '0;
              endcase
           end
           TRIGGER_IM_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {TRIGGER_IM[0]};
                 default: read_data = '0;
              endcase
           end
           TRIGGER_IM_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {TRIGGER_IM[1]};
                 default: read_data = '0;
              endcase
           end
           TRIGGER_RATE_LIM_EMPTY_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {TRIGGER_RATE_LIM_EMPTY};
                 default: read_data = '0;
              endcase
           end
           {44'h1?,1'b?},
           {40'b1?,4'h?,1'b?},
           {40'b1??,4'h?,1'b?},
           {40'b1???,4'h?,1'b?},
           {44'h10?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_MA_TCN_FIFO_0;
                 default: read_data = '0;
              endcase
           end
           {44'h11?,1'b?},
           {36'h1,4'b001?,4'h?,1'b?},
           {36'h1,4'b01??,4'h?,1'b?},
           {36'h1,4'b1???,4'h?,1'b?},
           {44'h20?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_MA_TCN_FIFO_1;
                 default: read_data = '0;
              endcase
           end
           {44'h210,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_MA_TCN_DEQUEUE;
                 default: read_data = '0;
              endcase
           end
           {44'h210,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_MA_TCN_DATA_0;
                 default: read_data = '0;
              endcase
           end
           {44'h211,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_MA_TCN_DATA_1;
                 default: read_data = '0;
              endcase
           end
           {44'h211,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_MA_TCN_PTR_HEAD;
                 default: read_data = '0;
              endcase
           end
           {44'h212,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = handcode_reg_rdata_MA_TCN_PTR_TAIL;
                 default: read_data = '0;
              endcase
           end
           MA_TCN_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_IP};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_IM};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[0]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[1]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[2]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[3]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[4]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[5]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[6]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[7]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[8]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[9]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[10]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[11]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[12]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[13]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[14]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[15]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_WM_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_WM[16]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[0]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[0]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[1]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[1]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[2]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[2]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[3]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[3]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[4]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[4]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[5]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[5]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[6]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[6]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[7]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[7]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[8]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[8]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[9]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[9]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[10]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[10]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[11]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[11]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[12]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[12]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[13]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[13]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[14]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[14]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[15]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[15]};
                 default: read_data = '0;
              endcase
           end
           MA_TCN_USAGE_DECODE_ADDR[16]: begin
              unique casez ({req_fid,req_bar})
                 {TRIG_APPLY_MISC_SB_FID,TRIG_APPLY_MISC_SB_BAR}: read_data = {MA_TCN_USAGE[16]};
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    TRIGGER_IP[0].reserved0 = '0;
    TRIGGER_IP[1].reserved0 = '0;
    TRIGGER_IM[0].reserved0 = '0;
    TRIGGER_IM[1].reserved0 = '0;
    TRIGGER_RATE_LIM_EMPTY.reserved0 = '0;
    MA_TCN_IP.reserved0 = '0;
    MA_TCN_IM.reserved0 = '0;
    MA_TCN_WM[0].reserved0 = '0;
    MA_TCN_WM[1].reserved0 = '0;
    MA_TCN_WM[2].reserved0 = '0;
    MA_TCN_WM[3].reserved0 = '0;
    MA_TCN_WM[4].reserved0 = '0;
    MA_TCN_WM[5].reserved0 = '0;
    MA_TCN_WM[6].reserved0 = '0;
    MA_TCN_WM[7].reserved0 = '0;
    MA_TCN_WM[8].reserved0 = '0;
    MA_TCN_WM[9].reserved0 = '0;
    MA_TCN_WM[10].reserved0 = '0;
    MA_TCN_WM[11].reserved0 = '0;
    MA_TCN_WM[12].reserved0 = '0;
    MA_TCN_WM[13].reserved0 = '0;
    MA_TCN_WM[14].reserved0 = '0;
    MA_TCN_WM[15].reserved0 = '0;
    MA_TCN_WM[16].reserved0 = '0;
    MA_TCN_USAGE[0].reserved0 = '0;
    MA_TCN_USAGE[1].reserved0 = '0;
    MA_TCN_USAGE[2].reserved0 = '0;
    MA_TCN_USAGE[3].reserved0 = '0;
    MA_TCN_USAGE[4].reserved0 = '0;
    MA_TCN_USAGE[5].reserved0 = '0;
    MA_TCN_USAGE[6].reserved0 = '0;
    MA_TCN_USAGE[7].reserved0 = '0;
    MA_TCN_USAGE[8].reserved0 = '0;
    MA_TCN_USAGE[9].reserved0 = '0;
    MA_TCN_USAGE[10].reserved0 = '0;
    MA_TCN_USAGE[11].reserved0 = '0;
    MA_TCN_USAGE[12].reserved0 = '0;
    MA_TCN_USAGE[13].reserved0 = '0;
    MA_TCN_USAGE[14].reserved0 = '0;
    MA_TCN_USAGE[15].reserved0 = '0;
    MA_TCN_USAGE[16].reserved0 = '0;
end

// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
