magic
tech scmos
timestamp 970031125
<< ndiffusion >>
rect -34 459 -8 460
rect -34 455 -8 456
rect -34 447 -22 455
rect -34 446 -8 447
rect -34 442 -8 443
rect -34 433 -8 434
rect -34 429 -8 430
<< pdiffusion >>
rect 8 458 24 459
rect 8 449 24 450
rect 8 441 24 446
rect 8 433 24 438
rect 8 429 24 430
<< ntransistor >>
rect -34 456 -8 459
rect -34 443 -8 446
rect -34 430 -8 433
<< ptransistor >>
rect 8 446 24 449
rect 8 438 24 441
rect 8 430 24 433
<< polysilicon >>
rect -38 456 -34 459
rect -8 456 6 459
rect 3 449 6 456
rect 3 446 8 449
rect 24 446 28 449
rect -38 443 -34 446
rect -8 443 -3 446
rect -6 441 -3 443
rect -6 438 8 441
rect 24 438 28 441
rect -38 430 -34 433
rect -8 430 8 433
rect 24 430 28 433
<< ndcontact >>
rect -34 460 -8 468
rect -22 447 -8 455
rect -34 434 -8 442
rect -34 421 -8 429
<< pdcontact >>
rect 8 450 24 458
rect 8 421 24 429
<< psubstratepcontact >>
rect -51 456 -43 464
<< nsubstratencontact >>
rect 8 459 24 467
<< polycontact >>
rect -4 459 4 467
rect -46 443 -38 451
rect -46 430 -38 438
<< metal1 >>
rect -21 468 -8 469
rect -34 464 -8 468
rect 8 467 21 469
rect -51 460 -8 464
rect -4 463 4 467
rect -51 456 -26 460
rect -46 443 -38 445
rect -34 442 -26 456
rect -22 453 -8 455
rect -22 447 4 453
rect 8 450 24 467
rect -34 434 -8 442
rect -46 430 -38 433
rect -4 429 4 447
rect -34 427 24 429
rect -34 421 -4 427
rect 4 421 24 427
<< m2contact >>
rect -21 469 -8 475
rect 8 469 21 475
rect -4 457 4 463
rect -46 445 -38 451
rect -46 433 -38 439
rect -4 421 4 427
<< metal2 >>
rect -6 457 6 463
rect -46 445 0 451
rect -46 433 0 439
rect -6 421 6 427
<< m3contact >>
rect -21 469 -3 475
rect 3 469 21 475
<< metal3 >>
rect -21 418 -3 478
rect 3 418 21 478
<< labels >>
rlabel polysilicon -35 444 -35 444 1 b
rlabel polysilicon -35 431 -35 431 1 a
rlabel polysilicon -35 457 -35 457 1 c
rlabel metal2 0 433 0 439 7 a
rlabel metal2 0 445 0 451 7 b
rlabel polysilicon 25 431 25 431 7 a
rlabel polysilicon 25 439 25 439 7 b
rlabel polysilicon 25 447 25 447 7 c
rlabel metal1 -12 451 -12 451 5 x
rlabel metal1 -12 425 -12 425 1 x
rlabel metal1 -12 438 -12 438 5 GND!
rlabel metal1 -12 464 -12 464 5 GND!
rlabel metal1 16 425 16 425 1 x
rlabel metal2 0 421 0 427 1 x
rlabel metal1 16 454 16 454 1 Vdd!
rlabel metal2 0 457 0 463 3 c
rlabel metal1 -47 460 -47 460 3 GND!
rlabel space -52 420 -22 469 7 ^n
rlabel space 24 421 29 467 3 ^p
rlabel metal2 -42 448 -42 448 1 b
rlabel metal2 -42 436 -42 436 1 a
<< end >>
