magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -24 71 -20 72
rect -24 65 -20 69
rect -24 59 -20 63
rect -24 53 -20 57
rect -24 47 -20 51
rect -24 41 -20 45
rect -24 38 -20 39
<< pdiffusion >>
rect 3 76 5 80
rect -5 75 5 76
rect -5 72 5 73
rect -5 68 1 72
rect -5 67 5 68
rect -5 64 5 65
rect 3 60 5 64
rect -5 59 5 60
rect -5 56 5 57
rect -5 52 1 56
rect -5 51 5 52
rect -5 48 5 49
rect 3 44 5 48
rect -5 43 5 44
rect -5 40 5 41
rect -5 36 1 40
rect -5 34 3 36
rect -5 31 3 32
rect -1 28 3 31
<< ntransistor >>
rect -24 69 -20 71
rect -24 63 -20 65
rect -24 57 -20 59
rect -24 51 -20 53
rect -24 45 -20 47
rect -24 39 -20 41
<< ptransistor >>
rect -5 73 5 75
rect -5 65 5 67
rect -5 57 5 59
rect -5 49 5 51
rect -5 41 5 43
rect -5 32 3 34
<< polysilicon >>
rect -18 73 -5 75
rect 5 73 8 75
rect -18 71 -16 73
rect -27 69 -24 71
rect -20 69 -16 71
rect -9 65 -5 67
rect 5 65 8 67
rect -27 63 -24 65
rect -20 63 -7 65
rect -27 57 -24 59
rect -20 57 -5 59
rect 5 57 8 59
rect -27 51 -24 53
rect -20 51 -7 53
rect -9 49 -5 51
rect 5 49 8 51
rect -27 45 -24 47
rect -20 45 -12 47
rect -14 43 -12 45
rect -14 41 -5 43
rect 5 41 8 43
rect -27 39 -24 41
rect -20 39 -17 41
rect -8 32 -5 34
rect 3 32 6 34
<< ndcontact >>
rect -24 72 -20 76
rect -24 34 -20 38
<< pdcontact >>
rect -5 76 3 80
rect 1 68 5 72
rect -5 60 3 64
rect 1 52 5 56
rect -5 44 3 48
rect 1 36 5 40
rect -5 27 -1 31
<< metal1 >>
rect -5 76 3 80
rect -24 72 -2 76
rect -5 64 -2 72
rect 1 68 5 72
rect -5 60 3 64
rect -5 48 -2 60
rect 1 52 5 56
rect -5 44 3 48
rect -24 34 -20 38
rect -5 31 -2 44
rect 1 36 5 40
rect -5 27 -1 31
<< labels >>
rlabel space 2 38 8 81 3 ^p
rlabel polysilicon 6 74 6 74 3 e
rlabel polysilicon 6 66 6 66 3 d
rlabel polysilicon 6 58 6 58 3 c
rlabel polysilicon 6 50 6 50 3 b
rlabel polysilicon 6 42 6 42 3 a
rlabel polysilicon -25 40 -25 40 3 _SReset!
rlabel space -27 34 -24 76 7 ^n
rlabel polysilicon -25 70 -25 70 3 e
rlabel polysilicon -25 46 -25 46 3 a
rlabel polysilicon -25 52 -25 52 3 b
rlabel polysilicon -25 58 -25 58 3 c
rlabel polysilicon -25 64 -25 64 3 d
rlabel polysilicon 4 33 4 33 8 _PReset!
rlabel pdcontact 3 54 3 54 1 Vdd!
rlabel pdcontact 3 70 3 70 5 Vdd!
rlabel pdcontact -1 62 -1 62 5 x
rlabel pdcontact -1 46 -1 46 5 x
rlabel pdcontact -1 78 -1 78 5 x
rlabel pdcontact 3 38 3 38 1 Vdd!
rlabel ndcontact -22 36 -22 36 5 GND!
rlabel ndcontact -22 74 -22 74 4 x
<< end >>
