magic
tech scmos
timestamp 965153727
<< ndiffusion >>
rect 401 536 427 537
rect 401 532 427 533
rect 401 524 413 532
rect 401 523 427 524
rect 401 519 427 520
rect 415 511 427 519
rect 401 510 427 511
rect 401 506 427 507
rect 401 498 413 506
rect 401 497 427 498
rect 401 493 427 494
<< pdiffusion >>
rect 443 536 469 537
rect 443 532 469 533
rect 457 524 469 532
rect 443 523 469 524
rect 443 519 469 520
rect 443 511 455 519
rect 443 510 469 511
rect 443 506 469 507
rect 457 498 469 506
rect 443 497 469 498
rect 443 493 469 494
<< ntransistor >>
rect 401 533 427 536
rect 401 520 427 523
rect 401 507 427 510
rect 401 494 427 497
<< ptransistor >>
rect 443 533 469 536
rect 443 520 469 523
rect 443 507 469 510
rect 443 494 469 497
<< polysilicon >>
rect 397 533 401 536
rect 427 533 443 536
rect 469 533 473 536
rect 431 523 439 533
rect 397 520 401 523
rect 427 520 443 523
rect 469 520 473 523
rect 431 512 439 520
rect 397 507 401 510
rect 427 507 431 510
rect 397 494 401 497
rect 427 494 431 497
rect 439 507 443 510
rect 469 507 473 510
rect 439 494 443 497
rect 469 494 473 497
<< ndcontact >>
rect 401 537 427 545
rect 413 524 427 532
rect 401 511 415 519
rect 413 498 427 506
rect 401 485 427 493
<< pdcontact >>
rect 443 537 469 545
rect 443 524 457 532
rect 455 511 469 519
rect 443 498 457 506
rect 443 485 469 493
<< polycontact >>
rect 431 494 439 512
<< metal1 >>
rect 401 537 427 545
rect 443 537 469 545
rect 401 519 409 537
rect 413 524 457 532
rect 401 511 415 519
rect 419 516 451 524
rect 461 519 469 537
rect 401 493 409 511
rect 419 506 427 516
rect 413 498 427 506
rect 431 494 439 512
rect 443 506 451 516
rect 455 511 469 519
rect 443 498 457 506
rect 461 493 469 511
rect 401 485 427 493
rect 443 485 469 493
<< labels >>
rlabel ndcontact 408 489 408 489 1 GND!
rlabel ndcontact 408 515 408 515 5 GND!
rlabel ndcontact 408 541 408 541 5 GND!
rlabel ndcontact 420 528 420 528 1 x
rlabel ndcontact 420 502 420 502 1 x
rlabel pdcontact 451 528 451 528 1 x
rlabel pdcontact 451 502 451 502 1 x
rlabel pdcontact 461 489 461 489 1 Vdd!
rlabel pdcontact 461 515 461 515 5 Vdd!
rlabel pdcontact 461 541 461 541 5 Vdd!
rlabel space 396 484 414 546 7 ^n
rlabel space 456 484 474 546 3 ^p
rlabel metal1 435 503 435 503 1 a
<< end >>
