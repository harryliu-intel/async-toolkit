///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Jon Bagge <jon.bagge.com> 
// -- Project Name : MBY 
// -- Description  : PPE shared table memory netlist. 
// ------------------------------------------------------------------- 

module ppe_stm_top (
input logic reset, 
//Input List
input                   cclk,                                     
input           [98:0]  i_ibus_ctrl,                              

//Interface List
egr_ppe_stm_if.stm                egr_ppe_stm_if0,  
egr_ppe_stm_if.stm                egr_ppe_stm_if1,  
egr_mc_table_if.mc_table          mc_table_if0_0,  
egr_mc_table_if.mc_table          mc_table_if0_1,  
egr_mc_table_if.mc_table          mc_table_if1_0,  
egr_mc_table_if.mc_table          mc_table_if1_1,  
rx_ppe_ppe_stm0_if.stm            rx_ppe_ppe_stm0_if0,  
rx_ppe_ppe_stm0_if.stm            rx_ppe_ppe_stm0_if1,  
rx_ppe_ppe_stm1_if.stm            rx_ppe_ppe_stm1_if0,  
rx_ppe_ppe_stm1_if.stm            rx_ppe_ppe_stm1_if1,  

//Output List
output          [66:0]  o_ibus_resp                               
);

logic [47:0][3:0][11:0] fwd_tbl0_addr;                  
logic [47:0][3:0][71:0] fwd_tbl0_rdata;                 
logic [15:0][3:0][10:0] fwd_tbl1_addr;                  
logic [15:0][3:0][71:0] fwd_tbl1_rdata;                 
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_0_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_0_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_100_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_100_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_101_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_101_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_102_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_102_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_103_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_103_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_104_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_104_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_105_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_105_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_106_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_106_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_107_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_107_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_108_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_108_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_109_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_109_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_10_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_10_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_110_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_110_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_111_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_111_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_112_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_112_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_113_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_113_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_114_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_114_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_115_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_115_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_116_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_116_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_117_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_117_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_118_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_118_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_119_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_119_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_11_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_11_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_120_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_120_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_121_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_121_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_122_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_122_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_123_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_123_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_124_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_124_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_125_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_125_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_126_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_126_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_127_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_127_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_128_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_128_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_129_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_129_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_12_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_12_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_130_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_130_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_131_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_131_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_132_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_132_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_133_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_133_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_134_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_134_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_135_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_135_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_136_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_136_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_137_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_137_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_138_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_138_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_139_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_139_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_13_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_13_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_140_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_140_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_141_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_141_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_142_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_142_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_143_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_143_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_144_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_144_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_145_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_145_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_146_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_146_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_147_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_147_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_148_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_148_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_149_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_149_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_14_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_14_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_150_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_150_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_151_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_151_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_152_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_152_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_153_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_153_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_154_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_154_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_155_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_155_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_156_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_156_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_157_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_157_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_158_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_158_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_159_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_159_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_15_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_15_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_160_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_160_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_161_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_161_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_162_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_162_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_163_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_163_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_164_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_164_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_165_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_165_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_166_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_166_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_167_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_167_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_168_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_168_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_169_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_169_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_16_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_16_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_170_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_170_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_171_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_171_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_172_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_172_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_173_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_173_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_174_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_174_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_175_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_175_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_176_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_176_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_177_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_177_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_178_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_178_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_179_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_179_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_17_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_17_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_180_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_180_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_181_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_181_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_182_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_182_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_183_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_183_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_184_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_184_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_185_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_185_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_186_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_186_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_187_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_187_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_188_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_188_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_189_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_189_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_18_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_18_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_190_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_190_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_191_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_191_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_19_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_19_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_1_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_1_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_20_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_20_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_21_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_21_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_22_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_22_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_23_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_23_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_24_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_24_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_25_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_25_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_26_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_26_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_27_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_27_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_28_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_28_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_29_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_29_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_2_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_2_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_30_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_30_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_31_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_31_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_32_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_32_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_33_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_33_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_34_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_34_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_35_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_35_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_36_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_36_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_37_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_37_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_38_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_38_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_39_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_39_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_3_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_3_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_40_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_40_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_41_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_41_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_42_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_42_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_43_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_43_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_44_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_44_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_45_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_45_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_46_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_46_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_47_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_47_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_48_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_48_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_49_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_49_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_4_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_4_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_50_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_50_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_51_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_51_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_52_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_52_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_53_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_53_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_54_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_54_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_55_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_55_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_56_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_56_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_57_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_57_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_58_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_58_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_59_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_59_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_5_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_5_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_60_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_60_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_61_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_61_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_62_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_62_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_63_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_63_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_64_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_64_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_65_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_65_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_66_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_66_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_67_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_67_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_68_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_68_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_69_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_69_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_6_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_6_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_70_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_70_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_71_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_71_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_72_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_72_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_73_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_73_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_74_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_74_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_75_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_75_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_76_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_76_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_77_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_77_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_78_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_78_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_79_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_79_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_7_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_7_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_80_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_80_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_81_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_81_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_82_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_82_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_83_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_83_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_84_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_84_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_85_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_85_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_86_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_86_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_87_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_87_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_88_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_88_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_89_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_89_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_8_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_8_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_90_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_90_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_91_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_91_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_92_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_92_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_93_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_93_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_94_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_94_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_95_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_95_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_96_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_96_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_97_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_97_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_98_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_98_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_99_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_99_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl0_9_from_mem;
logic            [92:0] ppe_stm_ppe_stm_fwd_tbl0_9_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_0_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_0_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_10_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_10_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_11_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_11_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_12_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_12_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_13_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_13_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_14_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_14_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_15_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_15_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_16_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_16_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_17_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_17_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_18_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_18_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_19_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_19_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_1_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_1_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_20_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_20_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_21_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_21_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_22_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_22_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_23_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_23_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_24_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_24_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_25_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_25_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_26_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_26_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_27_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_27_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_28_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_28_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_29_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_29_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_2_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_2_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_30_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_30_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_31_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_31_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_32_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_32_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_33_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_33_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_34_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_34_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_35_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_35_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_36_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_36_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_37_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_37_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_38_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_38_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_39_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_39_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_3_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_3_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_40_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_40_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_41_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_41_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_42_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_42_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_43_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_43_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_44_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_44_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_45_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_45_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_46_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_46_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_47_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_47_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_48_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_48_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_49_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_49_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_4_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_4_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_50_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_50_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_51_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_51_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_52_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_52_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_53_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_53_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_54_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_54_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_55_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_55_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_56_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_56_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_57_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_57_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_58_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_58_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_59_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_59_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_5_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_5_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_60_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_60_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_61_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_61_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_62_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_62_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_63_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_63_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_6_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_6_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_7_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_7_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_8_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_8_to_mem;
logic            [72:0] ppe_stm_ppe_stm_fwd_tbl1_9_from_mem;
logic            [91:0] ppe_stm_ppe_stm_fwd_tbl1_9_to_mem;
logic           [576:0] ppe_stm_ppe_stm_l3mc_tbl_from_mem;
logic           [596:0] ppe_stm_ppe_stm_l3mc_tbl_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_0_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_0_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_10_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_10_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_11_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_11_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_12_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_12_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_13_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_13_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_14_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_14_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_15_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_15_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_16_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_16_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_17_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_17_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_18_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_18_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_19_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_19_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_1_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_1_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_20_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_20_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_21_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_21_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_22_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_22_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_23_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_23_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_24_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_24_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_25_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_25_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_26_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_26_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_27_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_27_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_28_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_28_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_29_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_29_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_2_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_2_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_30_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_30_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_31_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_31_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_32_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_32_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_33_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_33_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_34_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_34_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_35_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_35_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_36_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_36_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_37_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_37_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_38_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_38_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_39_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_39_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_3_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_3_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_40_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_40_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_41_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_41_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_42_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_42_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_43_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_43_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_44_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_44_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_45_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_45_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_46_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_46_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_47_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_47_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_48_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_48_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_49_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_49_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_4_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_4_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_50_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_50_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_51_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_51_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_52_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_52_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_53_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_53_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_54_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_54_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_55_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_55_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_56_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_56_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_57_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_57_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_58_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_58_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_59_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_59_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_5_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_5_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_60_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_60_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_61_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_61_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_62_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_62_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_63_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_63_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_64_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_64_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_65_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_65_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_66_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_66_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_67_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_67_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_68_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_68_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_69_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_69_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_6_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_6_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_70_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_70_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_71_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_71_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_72_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_72_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_73_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_73_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_74_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_74_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_75_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_75_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_76_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_76_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_77_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_77_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_78_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_78_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_79_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_79_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_7_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_7_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_8_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_8_to_mem;
logic            [72:0] ppe_stm_ppe_stm_mod_tbl_9_from_mem;
logic            [91:0] ppe_stm_ppe_stm_mod_tbl_9_to_mem;
logic            [40:0] ppe_stm_ppe_stm_shcp_tbl_from_mem;
logic            [63:0] ppe_stm_ppe_stm_shcp_tbl_to_mem;
logic       [47:0][3:0] q_fwd_tbl0_ren;                 
logic       [3:0][71:0] q_fwd_tbl0_wdata;               
logic       [47:0][3:0] q_fwd_tbl0_wen;                 
logic       [15:0][3:0] q_fwd_tbl1_ren;                 
logic       [3:0][71:0] q_fwd_tbl1_wdata;               
logic       [15:0][3:0] q_fwd_tbl1_wen;                 
logic reset_n; 
assign reset_n = !reset;


// module ppe_stm_logic    from ppe_stm_logic using ppe_stm_logic.map 
ppe_stm_logic     #(.FWD_TBL0_BANKS(48),
                    .FWD_TBL0_CHUNKS(4),
                    .FWD_TBL0_RDATA_WIDTH(72),
                    .FWD_TBL0_MEM_SIZE(4096),
                    .LOG2_FWD_TBL0_MEM_SIZE(12),
                    .FWD_TBL0_RPORTS(6),
                    .FWD_TBL0_ADDR_WIDTH(20),
                    .FWD_TBL0_WDATA_WIDTH(72),
                    .FWD_TBL1_BANKS(16),
                    .FWD_TBL1_CHUNKS(4),
                    .FWD_TBL1_RDATA_WIDTH(72),
                    .FWD_TBL1_MEM_SIZE(2047),
                    .LOG2_FWD_TBL1_MEM_SIZE(11),
                    .FWD_TBL1_RPORTS(4),
                    .FWD_TBL1_ADDR_WIDTH(17),
                    .FWD_TBL1_WDATA_WIDTH(72)) ppe_stm_logic(
/* input  logic                          */ .cclk                (cclk),                                
/* input  logic  [48-1:0][4-1:0][72-1:0] */ .i_fwd_tbl0_rdata    (fwd_tbl0_rdata),                      
/* output logic          [48-1:0][4-1:0] */ .o_q_fwd_tbl0_ren    (q_fwd_tbl0_ren),                      
/* output logic          [48-1:0][4-1:0] */ .o_q_fwd_tbl0_wen    (q_fwd_tbl0_wen),                      
/* output logic  [48-1:0][4-1:0][12-1:0] */ .o_fwd_tbl0_addr     (fwd_tbl0_addr),                       
/* output logic          [4-1:0][72-1:0] */ .o_q_fwd_tbl0_wdata  (q_fwd_tbl0_wdata),                    
/* input  logic  [16-1:0][4-1:0][72-1:0] */ .i_fwd_tbl1_rdata    (fwd_tbl1_rdata),                      
/* output logic          [16-1:0][4-1:0] */ .o_q_fwd_tbl1_ren    (q_fwd_tbl1_ren),                      
/* output logic          [16-1:0][4-1:0] */ .o_q_fwd_tbl1_wen    (q_fwd_tbl1_wen),                      
/* output logic  [16-1:0][4-1:0][11-1:0] */ .o_fwd_tbl1_addr     (fwd_tbl1_addr),                       
/* output logic          [4-1:0][72-1:0] */ .o_q_fwd_tbl1_wdata  (q_fwd_tbl1_wdata),                    
/* input  logic                   [98:0] */ .i_ibus_ctrl         (i_ibus_ctrl),                         
/* output logic                   [66:0] */ .o_ibus_resp         (o_ibus_resp),                         
/* Interface rx_ppe_ppe_stm0_if.stm      */ .rx_ppe_ppe_stm0_if0 (rx_ppe_ppe_stm0_if0),                 
/* Interface rx_ppe_ppe_stm1_if.stm      */ .rx_ppe_ppe_stm1_if0 (rx_ppe_ppe_stm1_if0),                 
/* Interface rx_ppe_ppe_stm0_if.stm      */ .rx_ppe_ppe_stm0_if1 (rx_ppe_ppe_stm0_if1),                 
/* Interface rx_ppe_ppe_stm1_if.stm      */ .rx_ppe_ppe_stm1_if1 (rx_ppe_ppe_stm1_if1),                 
/* Interface egr_ppe_stm_if.stm          */ .egr_ppe_stm_if0     (egr_ppe_stm_if0),                     
/* Interface egr_ppe_stm_if.stm          */ .egr_ppe_stm_if1     (egr_ppe_stm_if1),                     
/* Interface egr_mc_table_if.mc_table    */ .mc_table_if0_0      (mc_table_if0_0),                      
/* Interface egr_mc_table_if.mc_table    */ .mc_table_if0_1      (mc_table_if0_1),                      
/* Interface egr_mc_table_if.mc_table    */ .mc_table_if1_0      (mc_table_if1_0),                      
/* Interface egr_mc_table_if.mc_table    */ .mc_table_if1_1      (mc_table_if1_1));                      
// End of module ppe_stm_logic from ppe_stm_logic


// module ppe_stm_shells_wrapper    from ppe_stm_shells_wrapper using ppe_stm_shells_wrapper.map 
ppe_stm_shells_wrapper    ppe_stm_shells_wrapper(
/* input  logic          */ .PPE_STM_FWD_TBL0_114_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_115_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_115_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_116_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_116_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_117_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_117_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_118_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_118_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_119_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_119_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_11_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_11_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_120_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_120_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_121_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_121_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_122_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_122_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_123_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_123_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_124_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_124_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_125_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_125_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_126_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_126_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_127_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_127_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_128_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_128_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_129_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_129_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_12_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_12_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_130_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_130_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_131_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_131_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_134_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_134_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_135_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_135_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_136_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_136_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_137_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_137_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_138_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_138_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_139_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_139_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_13_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_13_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_140_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_140_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_141_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_141_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_142_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_142_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_143_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_143_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_144_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_144_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_145_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_145_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_146_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_146_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_147_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_147_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_148_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_148_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_149_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_149_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_14_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_14_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_150_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_150_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_151_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_151_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_152_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_152_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_153_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_153_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_154_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_154_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_155_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_155_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_156_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_156_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_157_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_157_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_158_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_158_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_159_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_159_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_15_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_15_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_160_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_160_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_161_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_161_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_162_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_162_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_163_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_163_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_164_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_164_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_165_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_165_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_166_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_166_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_167_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_167_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_168_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_168_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_169_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_169_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_16_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_16_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_170_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_172_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_172_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_173_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_173_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_174_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_174_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_175_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_175_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_176_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_176_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_177_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_177_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_178_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_178_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_179_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_179_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_17_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_17_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_180_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_180_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_181_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_181_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_182_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_182_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_183_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_183_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_184_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_184_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_185_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_185_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_186_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_186_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_187_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_187_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_188_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_188_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_189_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_189_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_18_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_18_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_190_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_190_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_191_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_191_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_19_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_19_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_1_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_1_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_20_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_20_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_21_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_21_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_22_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_22_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_23_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_23_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_24_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_24_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_25_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_25_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_26_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_26_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_27_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_27_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_28_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_28_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_29_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_29_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_2_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_2_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_30_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_30_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_31_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_31_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_32_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_32_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_33_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_33_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_34_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_34_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_35_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_35_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_36_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_36_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_37_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_39_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_3_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_3_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_40_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_40_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_41_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_41_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_42_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_42_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_43_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_43_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_44_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_44_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_45_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_45_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_46_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_46_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_47_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_47_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_48_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_48_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_49_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_49_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_4_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_4_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_50_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_50_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_51_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_51_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_52_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_52_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_53_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_53_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_54_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_54_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_55_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_55_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_56_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_56_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_57_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_57_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_58_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_58_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_59_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_59_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_5_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_5_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_60_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_60_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_61_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_61_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_62_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_62_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_63_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_63_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_64_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_64_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_65_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_65_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_66_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_66_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_67_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_67_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_68_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_68_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_69_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_69_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_6_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_6_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_70_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_70_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_71_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_71_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_72_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_72_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_73_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_73_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_74_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_74_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_75_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_77_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_78_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_78_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_79_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_79_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_7_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_7_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_80_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_80_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_81_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_81_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_82_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_82_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_83_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_83_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_84_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_84_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_85_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_85_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_86_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_86_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_87_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_87_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_88_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_88_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_89_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_89_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_8_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_8_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_90_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_90_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_91_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_91_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_92_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_92_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_93_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_93_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_94_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_94_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_95_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_95_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_96_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_96_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_97_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_97_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_98_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_98_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_99_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_99_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_9_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_9_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_0_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_0_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_10_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_10_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_11_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_11_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_12_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_12_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_13_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_13_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_14_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_14_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_15_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_15_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_16_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_16_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_17_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_17_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_18_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_18_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_19_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_19_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_1_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_1_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_20_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_20_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_21_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_21_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_22_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_22_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_23_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_23_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_24_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_24_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_27_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_27_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_28_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_28_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_29_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_29_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_2_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_2_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_30_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_30_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_31_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_31_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_32_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_32_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_33_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_33_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_34_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_34_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_35_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_35_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_36_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_36_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_37_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_37_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_38_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_38_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_39_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_39_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_3_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_3_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_40_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_40_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_41_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_41_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_42_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_42_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_43_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_43_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_44_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_44_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_45_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_45_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_46_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_46_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_47_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_47_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_48_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_48_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_49_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_49_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_4_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_4_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_50_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_50_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_51_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_51_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_52_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_52_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_53_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_53_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_54_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_54_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_55_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_55_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_56_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_56_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_57_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_57_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_58_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_58_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_59_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_59_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_5_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_5_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_60_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_60_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_61_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_61_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_62_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_62_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_7_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_7_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_8_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_8_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_9_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_9_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_L3MC_TBL_CFG_reg_sel          (),                                                
/* input  logic          */ .PPE_STM_L3MC_TBL_STATUS_reg_sel       (),                                                
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_162_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_162_wr_en            (q_fwd_tbl0_wen[40][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_163_adr              (fwd_tbl0_addr[40][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_163_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_163_rd_en            (q_fwd_tbl0_ren[40][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_163_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_163_wr_en            (q_fwd_tbl0_wen[40][3]),                           
/* input  logic          */ .PPE_STM_MOD_TBL_0_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_0_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_10_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_10_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_11_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_11_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_12_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_12_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_13_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_13_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_14_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_14_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_15_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_15_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_16_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_16_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_17_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_17_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_18_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_18_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_19_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_19_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_1_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_1_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_20_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_20_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_21_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_21_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_22_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_22_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_23_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_23_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_24_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_24_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_25_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_25_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_26_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_26_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_27_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_27_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_28_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_28_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_29_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_29_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_2_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_2_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_30_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_30_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_31_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_31_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_32_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_32_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_33_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_33_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_34_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_34_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_35_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_35_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_36_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_36_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_37_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_37_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_38_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_38_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_39_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_39_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_3_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_3_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_40_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_40_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_41_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_41_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_42_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_42_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_43_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_43_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_44_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_46_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_47_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_47_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_48_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_48_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_49_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_49_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_4_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_4_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_50_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_50_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_51_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_51_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_52_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_52_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_53_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_53_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_54_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_54_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_55_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_55_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_56_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_56_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_57_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_57_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_58_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_58_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_59_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_59_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_5_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_5_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_60_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_60_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_61_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_61_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_62_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_62_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_63_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_63_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_64_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_64_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_65_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_65_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_66_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_66_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_67_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_67_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_68_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_68_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_69_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_69_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_6_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_6_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_70_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_70_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_71_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_71_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_72_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_72_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_73_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_73_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_74_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_74_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_75_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_75_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_76_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_76_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_77_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_77_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_78_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_78_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_79_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_79_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_7_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_7_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_8_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_8_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_9_CFG_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_9_STATUS_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_SHCP_TBL_CFG_reg_sel          (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_0_rd_en              (q_fwd_tbl0_ren[0][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_0_wr_data            (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_0_wr_en              (q_fwd_tbl0_wen[0][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_100_adr              (fwd_tbl0_addr[25][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_100_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_100_rd_en            (q_fwd_tbl0_ren[25][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_100_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_100_wr_en            (q_fwd_tbl0_wen[25][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_101_adr              (fwd_tbl0_addr[25][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_101_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_101_rd_en            (q_fwd_tbl0_ren[25][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_101_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_101_wr_en            (q_fwd_tbl0_wen[25][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_102_adr              (fwd_tbl0_addr[25][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_102_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_102_rd_en            (q_fwd_tbl0_ren[25][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_102_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_102_wr_en            (q_fwd_tbl0_wen[25][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_103_adr              (fwd_tbl0_addr[25][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_103_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_103_rd_en            (q_fwd_tbl0_ren[25][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_103_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_103_wr_en            (q_fwd_tbl0_wen[25][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_104_adr              (fwd_tbl0_addr[26][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_104_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_104_rd_en            (q_fwd_tbl0_ren[26][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_104_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_104_wr_en            (q_fwd_tbl0_wen[26][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_105_adr              (fwd_tbl0_addr[26][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_105_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_105_rd_en            (q_fwd_tbl0_ren[26][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_105_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_105_wr_en            (q_fwd_tbl0_wen[26][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_106_adr              (fwd_tbl0_addr[26][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_106_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_106_rd_en            (q_fwd_tbl0_ren[26][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_106_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_106_wr_en            (q_fwd_tbl0_wen[26][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_107_adr              (fwd_tbl0_addr[26][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_107_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_107_rd_en            (q_fwd_tbl0_ren[26][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_107_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_107_wr_en            (q_fwd_tbl0_wen[26][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_108_adr              (fwd_tbl0_addr[27][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_108_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_108_rd_en            (q_fwd_tbl0_ren[27][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_108_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_108_wr_en            (q_fwd_tbl0_wen[27][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_109_adr              (fwd_tbl0_addr[27][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_109_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_109_rd_en            (q_fwd_tbl0_ren[27][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_109_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_109_wr_en            (q_fwd_tbl0_wen[27][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_10_adr               (fwd_tbl0_addr[2][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_10_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_10_rd_en             (q_fwd_tbl0_ren[2][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_10_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_10_wr_en             (q_fwd_tbl0_wen[2][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_110_adr              (fwd_tbl0_addr[27][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_110_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_110_rd_en            (q_fwd_tbl0_ren[27][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_110_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_110_wr_en            (q_fwd_tbl0_wen[27][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_111_adr              (fwd_tbl0_addr[27][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_111_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_111_rd_en            (q_fwd_tbl0_ren[27][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_111_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_111_wr_en            (q_fwd_tbl0_wen[27][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_112_adr              (fwd_tbl0_addr[28][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_112_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_112_rd_en            (q_fwd_tbl0_ren[28][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_112_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_112_wr_en            (q_fwd_tbl0_wen[28][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_113_adr              (fwd_tbl0_addr[28][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_113_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_113_rd_en            (q_fwd_tbl0_ren[28][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_113_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_113_wr_en            (q_fwd_tbl0_wen[28][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_114_adr              (fwd_tbl0_addr[28][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_114_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_114_rd_en            (q_fwd_tbl0_ren[28][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_114_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_114_wr_en            (q_fwd_tbl0_wen[28][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_115_adr              (fwd_tbl0_addr[28][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_115_mem_ls_enter     (),                                                
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_116_adr              (fwd_tbl0_addr[29][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_116_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_116_rd_en            (q_fwd_tbl0_ren[29][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_116_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_116_wr_en            (q_fwd_tbl0_wen[29][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_117_adr              (fwd_tbl0_addr[29][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_117_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_117_rd_en            (q_fwd_tbl0_ren[29][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_117_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_117_wr_en            (q_fwd_tbl0_wen[29][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_118_adr              (fwd_tbl0_addr[29][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_118_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_118_rd_en            (q_fwd_tbl0_ren[29][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_118_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_118_wr_en            (q_fwd_tbl0_wen[29][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_119_adr              (fwd_tbl0_addr[29][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_119_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_119_rd_en            (q_fwd_tbl0_ren[29][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_119_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_119_wr_en            (q_fwd_tbl0_wen[29][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_11_adr               (fwd_tbl0_addr[2][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_11_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_11_rd_en             (q_fwd_tbl0_ren[2][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_11_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_11_wr_en             (q_fwd_tbl0_wen[2][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_120_adr              (fwd_tbl0_addr[30][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_120_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_120_rd_en            (q_fwd_tbl0_ren[30][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_120_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_120_wr_en            (q_fwd_tbl0_wen[30][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_121_adr              (fwd_tbl0_addr[30][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_121_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_121_rd_en            (q_fwd_tbl0_ren[30][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_121_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_121_wr_en            (q_fwd_tbl0_wen[30][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_122_adr              (fwd_tbl0_addr[30][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_122_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_122_rd_en            (q_fwd_tbl0_ren[30][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_122_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_122_wr_en            (q_fwd_tbl0_wen[30][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_123_adr              (fwd_tbl0_addr[30][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_123_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_123_rd_en            (q_fwd_tbl0_ren[30][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_123_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_123_wr_en            (q_fwd_tbl0_wen[30][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_124_adr              (fwd_tbl0_addr[31][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_124_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_124_rd_en            (q_fwd_tbl0_ren[31][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_124_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_124_wr_en            (q_fwd_tbl0_wen[31][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_125_adr              (fwd_tbl0_addr[31][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_125_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_125_rd_en            (q_fwd_tbl0_ren[31][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_125_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_125_wr_en            (q_fwd_tbl0_wen[31][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_126_adr              (fwd_tbl0_addr[31][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_126_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_126_rd_en            (q_fwd_tbl0_ren[31][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_126_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_126_wr_en            (q_fwd_tbl0_wen[31][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_127_adr              (fwd_tbl0_addr[31][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_127_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_127_rd_en            (q_fwd_tbl0_ren[31][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_127_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_127_wr_en            (q_fwd_tbl0_wen[31][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_128_adr              (fwd_tbl0_addr[32][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_128_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_128_rd_en            (q_fwd_tbl0_ren[32][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_128_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_128_wr_en            (q_fwd_tbl0_wen[32][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_129_adr              (fwd_tbl0_addr[32][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_129_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_129_rd_en            (q_fwd_tbl0_ren[32][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_129_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_129_wr_en            (q_fwd_tbl0_wen[32][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_12_adr               (fwd_tbl0_addr[3][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_12_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_12_rd_en             (q_fwd_tbl0_ren[3][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_12_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_12_wr_en             (q_fwd_tbl0_wen[3][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_130_adr              (fwd_tbl0_addr[32][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_131_adr              (fwd_tbl0_addr[32][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_131_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_131_rd_en            (q_fwd_tbl0_ren[32][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_131_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_131_wr_en            (q_fwd_tbl0_wen[32][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_132_adr              (fwd_tbl0_addr[33][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_132_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_132_rd_en            (q_fwd_tbl0_ren[33][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_132_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_132_wr_en            (q_fwd_tbl0_wen[33][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_133_adr              (fwd_tbl0_addr[33][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_133_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_133_rd_en            (q_fwd_tbl0_ren[33][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_133_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_133_wr_en            (q_fwd_tbl0_wen[33][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_134_adr              (fwd_tbl0_addr[33][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_134_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_134_rd_en            (q_fwd_tbl0_ren[33][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_134_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_134_wr_en            (q_fwd_tbl0_wen[33][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_135_adr              (fwd_tbl0_addr[33][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_135_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_135_rd_en            (q_fwd_tbl0_ren[33][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_135_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_135_wr_en            (q_fwd_tbl0_wen[33][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_136_adr              (fwd_tbl0_addr[34][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_136_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_136_rd_en            (q_fwd_tbl0_ren[34][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_136_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_136_wr_en            (q_fwd_tbl0_wen[34][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_137_adr              (fwd_tbl0_addr[34][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_137_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_137_rd_en            (q_fwd_tbl0_ren[34][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_137_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_137_wr_en            (q_fwd_tbl0_wen[34][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_138_adr              (fwd_tbl0_addr[34][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_138_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_138_rd_en            (q_fwd_tbl0_ren[34][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_138_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_138_wr_en            (q_fwd_tbl0_wen[34][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_139_adr              (fwd_tbl0_addr[34][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_139_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_139_rd_en            (q_fwd_tbl0_ren[34][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_139_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_139_wr_en            (q_fwd_tbl0_wen[34][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_13_adr               (fwd_tbl0_addr[3][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_13_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_13_rd_en             (q_fwd_tbl0_ren[3][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_13_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_13_wr_en             (q_fwd_tbl0_wen[3][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_140_adr              (fwd_tbl0_addr[35][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_140_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_140_rd_en            (q_fwd_tbl0_ren[35][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_140_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_140_wr_en            (q_fwd_tbl0_wen[35][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_141_adr              (fwd_tbl0_addr[35][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_141_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_141_rd_en            (q_fwd_tbl0_ren[35][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_141_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_141_wr_en            (q_fwd_tbl0_wen[35][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_142_adr              (fwd_tbl0_addr[35][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_142_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_142_rd_en            (q_fwd_tbl0_ren[35][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_142_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_142_wr_en            (q_fwd_tbl0_wen[35][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_143_adr              (fwd_tbl0_addr[35][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_143_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_143_rd_en            (q_fwd_tbl0_ren[35][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_143_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_143_wr_en            (q_fwd_tbl0_wen[35][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_144_adr              (fwd_tbl0_addr[36][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_144_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_144_rd_en            (q_fwd_tbl0_ren[36][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_144_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_144_wr_en            (q_fwd_tbl0_wen[36][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_145_adr              (fwd_tbl0_addr[36][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_145_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_145_rd_en            (q_fwd_tbl0_ren[36][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_145_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_145_wr_en            (q_fwd_tbl0_wen[36][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_146_adr              (fwd_tbl0_addr[36][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_146_wr_en            (q_fwd_tbl0_wen[36][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_147_adr              (fwd_tbl0_addr[36][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_147_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_147_rd_en            (q_fwd_tbl0_ren[36][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_147_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_147_wr_en            (q_fwd_tbl0_wen[36][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_148_adr              (fwd_tbl0_addr[37][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_148_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_148_rd_en            (q_fwd_tbl0_ren[37][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_148_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_148_wr_en            (q_fwd_tbl0_wen[37][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_149_adr              (fwd_tbl0_addr[37][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_149_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_149_rd_en            (q_fwd_tbl0_ren[37][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_149_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_149_wr_en            (q_fwd_tbl0_wen[37][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_14_adr               (fwd_tbl0_addr[3][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_14_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_14_rd_en             (q_fwd_tbl0_ren[3][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_14_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_14_wr_en             (q_fwd_tbl0_wen[3][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_150_adr              (fwd_tbl0_addr[37][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_150_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_150_rd_en            (q_fwd_tbl0_ren[37][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_150_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_150_wr_en            (q_fwd_tbl0_wen[37][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_151_adr              (fwd_tbl0_addr[37][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_151_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_151_rd_en            (q_fwd_tbl0_ren[37][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_151_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_151_wr_en            (q_fwd_tbl0_wen[37][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_152_adr              (fwd_tbl0_addr[38][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_152_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_152_rd_en            (q_fwd_tbl0_ren[38][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_152_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_152_wr_en            (q_fwd_tbl0_wen[38][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_153_adr              (fwd_tbl0_addr[38][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_153_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_153_rd_en            (q_fwd_tbl0_ren[38][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_153_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_153_wr_en            (q_fwd_tbl0_wen[38][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_154_adr              (fwd_tbl0_addr[38][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_154_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_154_rd_en            (q_fwd_tbl0_ren[38][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_154_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_154_wr_en            (q_fwd_tbl0_wen[38][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_155_adr              (fwd_tbl0_addr[38][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_155_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_155_rd_en            (q_fwd_tbl0_ren[38][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_155_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_155_wr_en            (q_fwd_tbl0_wen[38][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_156_adr              (fwd_tbl0_addr[39][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_156_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_156_rd_en            (q_fwd_tbl0_ren[39][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_156_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_156_wr_en            (q_fwd_tbl0_wen[39][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_157_adr              (fwd_tbl0_addr[39][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_157_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_157_rd_en            (q_fwd_tbl0_ren[39][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_157_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_157_wr_en            (q_fwd_tbl0_wen[39][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_158_adr              (fwd_tbl0_addr[39][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_158_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_158_rd_en            (q_fwd_tbl0_ren[39][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_158_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_158_wr_en            (q_fwd_tbl0_wen[39][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_159_adr              (fwd_tbl0_addr[39][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_159_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_159_rd_en            (q_fwd_tbl0_ren[39][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_159_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_159_wr_en            (q_fwd_tbl0_wen[39][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_15_adr               (fwd_tbl0_addr[3][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_15_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_15_rd_en             (q_fwd_tbl0_ren[3][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_15_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_15_wr_en             (q_fwd_tbl0_wen[3][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_160_adr              (fwd_tbl0_addr[40][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_160_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_160_rd_en            (q_fwd_tbl0_ren[40][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_160_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_160_wr_en            (q_fwd_tbl0_wen[40][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_161_adr              (fwd_tbl0_addr[40][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_161_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_161_rd_en            (q_fwd_tbl0_ren[40][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_161_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_mod_tbl_24_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_24_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_24_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_24_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_25_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_25_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_25_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_25_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_25_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_26_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_26_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_26_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_26_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_26_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_27_adr                (),                                                
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_164_adr              (fwd_tbl0_addr[41][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_164_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_164_rd_en            (q_fwd_tbl0_ren[41][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_164_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_164_wr_en            (q_fwd_tbl0_wen[41][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_165_adr              (fwd_tbl0_addr[41][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_165_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_165_rd_en            (q_fwd_tbl0_ren[41][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_165_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_165_wr_en            (q_fwd_tbl0_wen[41][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_166_adr              (fwd_tbl0_addr[41][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_166_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_166_rd_en            (q_fwd_tbl0_ren[41][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_166_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_166_wr_en            (q_fwd_tbl0_wen[41][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_167_adr              (fwd_tbl0_addr[41][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_167_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_167_rd_en            (q_fwd_tbl0_ren[41][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_167_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_167_wr_en            (q_fwd_tbl0_wen[41][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_168_adr              (fwd_tbl0_addr[42][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_168_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_168_rd_en            (q_fwd_tbl0_ren[42][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_168_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_168_wr_en            (q_fwd_tbl0_wen[42][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_169_adr              (fwd_tbl0_addr[42][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_169_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_169_rd_en            (q_fwd_tbl0_ren[42][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_169_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_169_wr_en            (q_fwd_tbl0_wen[42][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_16_adr               (fwd_tbl0_addr[4][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_16_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_16_rd_en             (q_fwd_tbl0_ren[4][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_16_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_16_wr_en             (q_fwd_tbl0_wen[4][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_170_adr              (fwd_tbl0_addr[42][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_170_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_170_rd_en            (q_fwd_tbl0_ren[42][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_170_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_170_wr_en            (q_fwd_tbl0_wen[42][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_171_adr              (fwd_tbl0_addr[42][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_171_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_171_rd_en            (q_fwd_tbl0_ren[42][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_171_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_171_wr_en            (q_fwd_tbl0_wen[42][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_172_adr              (fwd_tbl0_addr[43][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_172_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_172_rd_en            (q_fwd_tbl0_ren[43][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_172_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_172_wr_en            (q_fwd_tbl0_wen[43][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_173_adr              (fwd_tbl0_addr[43][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_173_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_173_rd_en            (q_fwd_tbl0_ren[43][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_173_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_173_wr_en            (q_fwd_tbl0_wen[43][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_174_adr              (fwd_tbl0_addr[43][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_174_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_174_rd_en            (q_fwd_tbl0_ren[43][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_174_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_174_wr_en            (q_fwd_tbl0_wen[43][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_175_adr              (fwd_tbl0_addr[43][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_175_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_175_rd_en            (q_fwd_tbl0_ren[43][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_175_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_175_wr_en            (q_fwd_tbl0_wen[43][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_176_adr              (fwd_tbl0_addr[44][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_176_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_176_rd_en            (q_fwd_tbl0_ren[44][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_176_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_176_wr_en            (q_fwd_tbl0_wen[44][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_177_adr              (fwd_tbl0_addr[44][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_177_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_177_rd_en            (q_fwd_tbl0_ren[44][1]),                           
/* input  logic          */ .ppe_stm_fwd_tbl0_178_rd_en            (q_fwd_tbl0_ren[44][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_178_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_178_wr_en            (q_fwd_tbl0_wen[44][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_179_adr              (fwd_tbl0_addr[44][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_179_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_179_rd_en            (q_fwd_tbl0_ren[44][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_179_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_179_wr_en            (q_fwd_tbl0_wen[44][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_17_adr               (fwd_tbl0_addr[4][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_17_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_17_rd_en             (q_fwd_tbl0_ren[4][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_17_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_17_wr_en             (q_fwd_tbl0_wen[4][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_180_adr              (fwd_tbl0_addr[45][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_180_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_180_rd_en            (q_fwd_tbl0_ren[45][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_180_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_180_wr_en            (q_fwd_tbl0_wen[45][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_181_adr              (fwd_tbl0_addr[45][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_181_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_181_rd_en            (q_fwd_tbl0_ren[45][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_181_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_181_wr_en            (q_fwd_tbl0_wen[45][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_182_adr              (fwd_tbl0_addr[45][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_182_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_182_rd_en            (q_fwd_tbl0_ren[45][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_182_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_182_wr_en            (q_fwd_tbl0_wen[45][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_183_adr              (fwd_tbl0_addr[45][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_183_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_183_rd_en            (q_fwd_tbl0_ren[45][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_183_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_183_wr_en            (q_fwd_tbl0_wen[45][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_184_adr              (fwd_tbl0_addr[46][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_184_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_184_rd_en            (q_fwd_tbl0_ren[46][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_184_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_184_wr_en            (q_fwd_tbl0_wen[46][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_185_adr              (fwd_tbl0_addr[46][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_185_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_185_rd_en            (q_fwd_tbl0_ren[46][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_185_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_185_wr_en            (q_fwd_tbl0_wen[46][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_186_adr              (fwd_tbl0_addr[46][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_186_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_186_rd_en            (q_fwd_tbl0_ren[46][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_186_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_186_wr_en            (q_fwd_tbl0_wen[46][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_187_adr              (fwd_tbl0_addr[46][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_187_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_187_rd_en            (q_fwd_tbl0_ren[46][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_187_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_187_wr_en            (q_fwd_tbl0_wen[46][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_188_adr              (fwd_tbl0_addr[47][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_188_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_188_rd_en            (q_fwd_tbl0_ren[47][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_188_wr_data          (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_188_wr_en            (q_fwd_tbl0_wen[47][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_189_adr              (fwd_tbl0_addr[47][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_189_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_189_rd_en            (q_fwd_tbl0_ren[47][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_189_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_189_wr_en            (q_fwd_tbl0_wen[47][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_18_adr               (fwd_tbl0_addr[4][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_18_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_18_rd_en             (q_fwd_tbl0_ren[4][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_18_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_18_wr_en             (q_fwd_tbl0_wen[4][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_190_adr              (fwd_tbl0_addr[47][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_190_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_190_rd_en            (q_fwd_tbl0_ren[47][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_190_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_190_wr_en            (q_fwd_tbl0_wen[47][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_191_adr              (fwd_tbl0_addr[47][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_191_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_191_rd_en            (q_fwd_tbl0_ren[47][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_191_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_191_wr_en            (q_fwd_tbl0_wen[47][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_19_adr               (fwd_tbl0_addr[4][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_19_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_19_rd_en             (q_fwd_tbl0_ren[4][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_19_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_19_wr_en             (q_fwd_tbl0_wen[4][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_1_adr                (fwd_tbl0_addr[0][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_1_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_1_rd_en              (q_fwd_tbl0_ren[0][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_1_wr_data            (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_1_wr_en              (q_fwd_tbl0_wen[0][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_20_adr               (fwd_tbl0_addr[5][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_20_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_20_rd_en             (q_fwd_tbl0_ren[5][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_20_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_20_wr_en             (q_fwd_tbl0_wen[5][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_21_adr               (fwd_tbl0_addr[5][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_21_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_21_rd_en             (q_fwd_tbl0_ren[5][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_21_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_21_wr_en             (q_fwd_tbl0_wen[5][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_22_adr               (fwd_tbl0_addr[5][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_22_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_22_rd_en             (q_fwd_tbl0_ren[5][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_22_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_22_wr_en             (q_fwd_tbl0_wen[5][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_23_adr               (fwd_tbl0_addr[5][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_23_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_23_rd_en             (q_fwd_tbl0_ren[5][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_23_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_23_wr_en             (q_fwd_tbl0_wen[5][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_24_adr               (fwd_tbl0_addr[6][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_24_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_24_rd_en             (q_fwd_tbl0_ren[6][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_24_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_24_wr_en             (q_fwd_tbl0_wen[6][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_25_adr               (fwd_tbl0_addr[6][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_25_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_25_rd_en             (q_fwd_tbl0_ren[6][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_25_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_25_wr_en             (q_fwd_tbl0_wen[6][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_26_adr               (fwd_tbl0_addr[6][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_26_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_26_rd_en             (q_fwd_tbl0_ren[6][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_26_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_26_wr_en             (q_fwd_tbl0_wen[6][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_27_adr               (fwd_tbl0_addr[6][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_27_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_27_rd_en             (q_fwd_tbl0_ren[6][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_27_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_27_wr_en             (q_fwd_tbl0_wen[6][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_28_adr               (fwd_tbl0_addr[7][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_28_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_28_rd_en             (q_fwd_tbl0_ren[7][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_28_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_28_wr_en             (q_fwd_tbl0_wen[7][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_29_adr               (fwd_tbl0_addr[7][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_29_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_29_rd_en             (q_fwd_tbl0_ren[7][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_29_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_29_wr_en             (q_fwd_tbl0_wen[7][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_2_adr                (fwd_tbl0_addr[0][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_2_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_2_rd_en              (q_fwd_tbl0_ren[0][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_2_wr_data            (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_2_wr_en              (q_fwd_tbl0_wen[0][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_30_adr               (fwd_tbl0_addr[7][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_30_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_30_rd_en             (q_fwd_tbl0_ren[7][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_30_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_30_wr_en             (q_fwd_tbl0_wen[7][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_31_adr               (fwd_tbl0_addr[7][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_31_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_31_rd_en             (q_fwd_tbl0_ren[7][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_31_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_31_wr_en             (q_fwd_tbl0_wen[7][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_32_adr               (fwd_tbl0_addr[8][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_32_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_32_rd_en             (q_fwd_tbl0_ren[8][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_32_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_32_wr_en             (q_fwd_tbl0_wen[8][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_33_adr               (fwd_tbl0_addr[8][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_33_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_33_rd_en             (q_fwd_tbl0_ren[8][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_33_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_33_wr_en             (q_fwd_tbl0_wen[8][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_34_adr               (fwd_tbl0_addr[8][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_34_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_34_rd_en             (q_fwd_tbl0_ren[8][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_34_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_34_wr_en             (q_fwd_tbl0_wen[8][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_35_adr               (fwd_tbl0_addr[8][3]),                             
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_36_adr               (fwd_tbl0_addr[9][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_36_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_36_rd_en             (q_fwd_tbl0_ren[9][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_36_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_36_wr_en             (q_fwd_tbl0_wen[9][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_37_adr               (fwd_tbl0_addr[9][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_37_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_37_rd_en             (q_fwd_tbl0_ren[9][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_37_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_37_wr_en             (q_fwd_tbl0_wen[9][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_38_adr               (fwd_tbl0_addr[9][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_38_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_38_rd_en             (q_fwd_tbl0_ren[9][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_38_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_38_wr_en             (q_fwd_tbl0_wen[9][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_39_adr               (fwd_tbl0_addr[9][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_39_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_39_rd_en             (q_fwd_tbl0_ren[9][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_39_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_39_wr_en             (q_fwd_tbl0_wen[9][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_3_adr                (fwd_tbl0_addr[0][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_3_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_3_rd_en              (q_fwd_tbl0_ren[0][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_3_wr_data            (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_3_wr_en              (q_fwd_tbl0_wen[0][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_40_adr               (fwd_tbl0_addr[10][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_40_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_40_rd_en             (q_fwd_tbl0_ren[10][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_40_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_40_wr_en             (q_fwd_tbl0_wen[10][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_41_adr               (fwd_tbl0_addr[10][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_41_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_41_rd_en             (q_fwd_tbl0_ren[10][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_41_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_41_wr_en             (q_fwd_tbl0_wen[10][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_42_adr               (fwd_tbl0_addr[10][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_42_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_42_rd_en             (q_fwd_tbl0_ren[10][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_42_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_42_wr_en             (q_fwd_tbl0_wen[10][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_43_adr               (fwd_tbl0_addr[10][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_43_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_43_rd_en             (q_fwd_tbl0_ren[10][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_43_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_43_wr_en             (q_fwd_tbl0_wen[10][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_44_adr               (fwd_tbl0_addr[11][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_44_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_44_rd_en             (q_fwd_tbl0_ren[11][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_44_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_44_wr_en             (q_fwd_tbl0_wen[11][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_45_adr               (fwd_tbl0_addr[11][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_45_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_45_rd_en             (q_fwd_tbl0_ren[11][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_45_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_45_wr_en             (q_fwd_tbl0_wen[11][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_46_adr               (fwd_tbl0_addr[11][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_46_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_46_rd_en             (q_fwd_tbl0_ren[11][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_46_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_46_wr_en             (q_fwd_tbl0_wen[11][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_47_adr               (fwd_tbl0_addr[11][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_47_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_47_rd_en             (q_fwd_tbl0_ren[11][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_47_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_47_wr_en             (q_fwd_tbl0_wen[11][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_48_adr               (fwd_tbl0_addr[12][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_48_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_48_rd_en             (q_fwd_tbl0_ren[12][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_48_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_48_wr_en             (q_fwd_tbl0_wen[12][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_49_adr               (fwd_tbl0_addr[12][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_49_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_49_rd_en             (q_fwd_tbl0_ren[12][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_49_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_49_wr_en             (q_fwd_tbl0_wen[12][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_4_adr                (fwd_tbl0_addr[1][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_4_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_4_rd_en              (q_fwd_tbl0_ren[1][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_4_wr_data            (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_4_wr_en              (q_fwd_tbl0_wen[1][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_50_adr               (fwd_tbl0_addr[12][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_50_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_50_rd_en             (q_fwd_tbl0_ren[12][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_50_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_50_wr_en             (q_fwd_tbl0_wen[12][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_51_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_51_wr_en             (q_fwd_tbl0_wen[12][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_52_adr               (fwd_tbl0_addr[13][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_52_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_52_rd_en             (q_fwd_tbl0_ren[13][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_52_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_52_wr_en             (q_fwd_tbl0_wen[13][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_53_adr               (fwd_tbl0_addr[13][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_53_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_53_rd_en             (q_fwd_tbl0_ren[13][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_53_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_53_wr_en             (q_fwd_tbl0_wen[13][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_54_adr               (fwd_tbl0_addr[13][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_54_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_54_rd_en             (q_fwd_tbl0_ren[13][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_54_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_54_wr_en             (q_fwd_tbl0_wen[13][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_55_adr               (fwd_tbl0_addr[13][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_55_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_55_rd_en             (q_fwd_tbl0_ren[13][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_55_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_55_wr_en             (q_fwd_tbl0_wen[13][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_56_adr               (fwd_tbl0_addr[14][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_56_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_56_rd_en             (q_fwd_tbl0_ren[14][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_56_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_56_wr_en             (q_fwd_tbl0_wen[14][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_57_adr               (fwd_tbl0_addr[14][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_57_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_57_rd_en             (q_fwd_tbl0_ren[14][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_57_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_57_wr_en             (q_fwd_tbl0_wen[14][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_58_adr               (fwd_tbl0_addr[14][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_58_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_58_rd_en             (q_fwd_tbl0_ren[14][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_58_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_58_wr_en             (q_fwd_tbl0_wen[14][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_59_adr               (fwd_tbl0_addr[14][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_59_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_59_rd_en             (q_fwd_tbl0_ren[14][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_59_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_59_wr_en             (q_fwd_tbl0_wen[14][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_5_adr                (fwd_tbl0_addr[1][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_5_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_5_rd_en              (q_fwd_tbl0_ren[1][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_5_wr_data            (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_5_wr_en              (q_fwd_tbl0_wen[1][1]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_60_adr               (fwd_tbl0_addr[15][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_60_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_60_rd_en             (q_fwd_tbl0_ren[15][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_60_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_60_wr_en             (q_fwd_tbl0_wen[15][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_61_adr               (fwd_tbl0_addr[15][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_61_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_61_rd_en             (q_fwd_tbl0_ren[15][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_61_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_61_wr_en             (q_fwd_tbl0_wen[15][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_62_adr               (fwd_tbl0_addr[15][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_62_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_62_rd_en             (q_fwd_tbl0_ren[15][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_62_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_62_wr_en             (q_fwd_tbl0_wen[15][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_63_adr               (fwd_tbl0_addr[15][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_63_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_63_rd_en             (q_fwd_tbl0_ren[15][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_63_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_63_wr_en             (q_fwd_tbl0_wen[15][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_64_adr               (fwd_tbl0_addr[16][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_64_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_64_rd_en             (q_fwd_tbl0_ren[16][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_64_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_64_wr_en             (q_fwd_tbl0_wen[16][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_65_adr               (fwd_tbl0_addr[16][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_65_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_65_rd_en             (q_fwd_tbl0_ren[16][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_65_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_65_wr_en             (q_fwd_tbl0_wen[16][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_66_adr               (fwd_tbl0_addr[16][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_66_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_66_rd_en             (q_fwd_tbl0_ren[16][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_66_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_67_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_67_wr_en             (q_fwd_tbl0_wen[16][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_68_adr               (fwd_tbl0_addr[17][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_68_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_68_rd_en             (q_fwd_tbl0_ren[17][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_68_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_68_wr_en             (q_fwd_tbl0_wen[17][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_69_adr               (fwd_tbl0_addr[17][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_69_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_69_rd_en             (q_fwd_tbl0_ren[17][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_69_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_69_wr_en             (q_fwd_tbl0_wen[17][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_6_adr                (fwd_tbl0_addr[1][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_6_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_6_rd_en              (q_fwd_tbl0_ren[1][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_6_wr_data            (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_6_wr_en              (q_fwd_tbl0_wen[1][2]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_70_adr               (fwd_tbl0_addr[17][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_70_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_70_rd_en             (q_fwd_tbl0_ren[17][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_70_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_70_wr_en             (q_fwd_tbl0_wen[17][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_71_adr               (fwd_tbl0_addr[17][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_71_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_71_rd_en             (q_fwd_tbl0_ren[17][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_71_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_71_wr_en             (q_fwd_tbl0_wen[17][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_72_adr               (fwd_tbl0_addr[18][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_72_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_72_rd_en             (q_fwd_tbl0_ren[18][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_72_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_72_wr_en             (q_fwd_tbl0_wen[18][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_73_adr               (fwd_tbl0_addr[18][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_73_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_73_rd_en             (q_fwd_tbl0_ren[18][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_73_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_73_wr_en             (q_fwd_tbl0_wen[18][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_74_adr               (fwd_tbl0_addr[18][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_74_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_74_rd_en             (q_fwd_tbl0_ren[18][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_74_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_74_wr_en             (q_fwd_tbl0_wen[18][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_75_adr               (fwd_tbl0_addr[18][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_75_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_75_rd_en             (q_fwd_tbl0_ren[18][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_75_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_75_wr_en             (q_fwd_tbl0_wen[18][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_76_adr               (fwd_tbl0_addr[19][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_76_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_76_rd_en             (q_fwd_tbl0_ren[19][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_76_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_76_wr_en             (q_fwd_tbl0_wen[19][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_77_adr               (fwd_tbl0_addr[19][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_77_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_77_rd_en             (q_fwd_tbl0_ren[19][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_77_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_77_wr_en             (q_fwd_tbl0_wen[19][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_78_adr               (fwd_tbl0_addr[19][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_78_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_78_rd_en             (q_fwd_tbl0_ren[19][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_78_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_78_wr_en             (q_fwd_tbl0_wen[19][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_79_adr               (fwd_tbl0_addr[19][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_79_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_79_rd_en             (q_fwd_tbl0_ren[19][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_79_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_79_wr_en             (q_fwd_tbl0_wen[19][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_7_adr                (fwd_tbl0_addr[1][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_7_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_7_rd_en              (q_fwd_tbl0_ren[1][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_7_wr_data            (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_7_wr_en              (q_fwd_tbl0_wen[1][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_80_adr               (fwd_tbl0_addr[20][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_80_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_80_rd_en             (q_fwd_tbl0_ren[20][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_80_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_80_wr_en             (q_fwd_tbl0_wen[20][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_81_adr               (fwd_tbl0_addr[20][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_81_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_81_rd_en             (q_fwd_tbl0_ren[20][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_81_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_81_wr_en             (q_fwd_tbl0_wen[20][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_82_adr               (fwd_tbl0_addr[20][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_82_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_83_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_83_rd_en             (q_fwd_tbl0_ren[20][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_83_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_83_wr_en             (q_fwd_tbl0_wen[20][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_84_adr               (fwd_tbl0_addr[21][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_84_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_84_rd_en             (q_fwd_tbl0_ren[21][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_84_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_84_wr_en             (q_fwd_tbl0_wen[21][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_85_adr               (fwd_tbl0_addr[21][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_85_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_85_rd_en             (q_fwd_tbl0_ren[21][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_85_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_85_wr_en             (q_fwd_tbl0_wen[21][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_86_adr               (fwd_tbl0_addr[21][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_86_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_86_rd_en             (q_fwd_tbl0_ren[21][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_86_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_86_wr_en             (q_fwd_tbl0_wen[21][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_87_adr               (fwd_tbl0_addr[21][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_87_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_87_rd_en             (q_fwd_tbl0_ren[21][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_87_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_87_wr_en             (q_fwd_tbl0_wen[21][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_88_adr               (fwd_tbl0_addr[22][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_88_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_88_rd_en             (q_fwd_tbl0_ren[22][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_88_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_88_wr_en             (q_fwd_tbl0_wen[22][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_89_adr               (fwd_tbl0_addr[22][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_89_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_89_rd_en             (q_fwd_tbl0_ren[22][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_89_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_89_wr_en             (q_fwd_tbl0_wen[22][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_8_adr                (fwd_tbl0_addr[2][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_8_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_8_rd_en              (q_fwd_tbl0_ren[2][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_8_wr_data            (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_8_wr_en              (q_fwd_tbl0_wen[2][0]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_90_adr               (fwd_tbl0_addr[22][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_90_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_90_rd_en             (q_fwd_tbl0_ren[22][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_90_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_90_wr_en             (q_fwd_tbl0_wen[22][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_91_adr               (fwd_tbl0_addr[22][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_91_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_91_rd_en             (q_fwd_tbl0_ren[22][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_91_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_91_wr_en             (q_fwd_tbl0_wen[22][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_92_adr               (fwd_tbl0_addr[23][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_92_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_92_rd_en             (q_fwd_tbl0_ren[23][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_92_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_92_wr_en             (q_fwd_tbl0_wen[23][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_93_adr               (fwd_tbl0_addr[23][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_93_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_93_rd_en             (q_fwd_tbl0_ren[23][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_93_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_93_wr_en             (q_fwd_tbl0_wen[23][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_94_adr               (fwd_tbl0_addr[23][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_94_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_94_rd_en             (q_fwd_tbl0_ren[23][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_94_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_94_wr_en             (q_fwd_tbl0_wen[23][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_95_adr               (fwd_tbl0_addr[23][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_95_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_95_rd_en             (q_fwd_tbl0_ren[23][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_95_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_95_wr_en             (q_fwd_tbl0_wen[23][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_96_adr               (fwd_tbl0_addr[24][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_96_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_96_rd_en             (q_fwd_tbl0_ren[24][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_96_wr_data           (q_fwd_tbl0_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_96_wr_en             (q_fwd_tbl0_wen[24][0]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_97_adr               (fwd_tbl0_addr[24][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_97_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_97_rd_en             (q_fwd_tbl0_ren[24][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_97_wr_data           (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_97_wr_en             (q_fwd_tbl0_wen[24][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_98_adr               (fwd_tbl0_addr[24][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_98_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_99_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_99_rd_en             (q_fwd_tbl0_ren[24][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_99_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_99_wr_en             (q_fwd_tbl0_wen[24][3]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_9_adr                (fwd_tbl0_addr[2][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_9_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_9_rd_en              (q_fwd_tbl0_ren[2][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_9_wr_data            (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_9_wr_en              (q_fwd_tbl0_wen[2][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_0_adr                (fwd_tbl1_addr[0][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_0_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_0_rd_en              (q_fwd_tbl1_ren[0][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_0_wr_data            (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_0_wr_en              (q_fwd_tbl1_wen[0][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_10_adr               (fwd_tbl1_addr[2][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_10_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_10_rd_en             (q_fwd_tbl1_ren[2][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_10_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_10_wr_en             (q_fwd_tbl1_wen[2][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_11_adr               (fwd_tbl1_addr[2][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_11_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_11_rd_en             (q_fwd_tbl1_ren[2][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_11_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_11_wr_en             (q_fwd_tbl1_wen[2][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_12_adr               (fwd_tbl1_addr[3][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_12_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_12_rd_en             (q_fwd_tbl1_ren[3][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_12_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_12_wr_en             (q_fwd_tbl1_wen[3][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_13_adr               (fwd_tbl1_addr[3][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_13_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_13_rd_en             (q_fwd_tbl1_ren[3][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_13_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_13_wr_en             (q_fwd_tbl1_wen[3][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_14_adr               (fwd_tbl1_addr[3][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_14_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_14_rd_en             (q_fwd_tbl1_ren[3][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_14_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_14_wr_en             (q_fwd_tbl1_wen[3][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_15_adr               (fwd_tbl1_addr[3][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_15_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_15_rd_en             (q_fwd_tbl1_ren[3][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_15_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_15_wr_en             (q_fwd_tbl1_wen[3][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_16_adr               (fwd_tbl1_addr[4][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_16_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_16_rd_en             (q_fwd_tbl1_ren[4][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_16_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_16_wr_en             (q_fwd_tbl1_wen[4][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_17_adr               (fwd_tbl1_addr[4][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_17_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_17_rd_en             (q_fwd_tbl1_ren[4][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_17_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_17_wr_en             (q_fwd_tbl1_wen[4][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_18_adr               (fwd_tbl1_addr[4][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_18_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_18_rd_en             (q_fwd_tbl1_ren[4][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_18_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_18_wr_en             (q_fwd_tbl1_wen[4][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_19_adr               (fwd_tbl1_addr[4][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_19_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_19_rd_en             (q_fwd_tbl1_ren[4][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_19_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_19_wr_en             (q_fwd_tbl1_wen[4][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_1_adr                (fwd_tbl1_addr[0][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_1_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_1_rd_en              (q_fwd_tbl1_ren[0][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_1_wr_data            (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_1_wr_en              (q_fwd_tbl1_wen[0][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_20_adr               (fwd_tbl1_addr[5][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_20_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_20_rd_en             (q_fwd_tbl1_ren[5][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_20_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_20_wr_en             (q_fwd_tbl1_wen[5][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_21_adr               (fwd_tbl1_addr[5][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_21_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_21_rd_en             (q_fwd_tbl1_ren[5][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_21_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_21_wr_en             (q_fwd_tbl1_wen[5][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_22_adr               (fwd_tbl1_addr[5][2]),                             
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_23_adr               (fwd_tbl1_addr[5][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_23_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_23_rd_en             (q_fwd_tbl1_ren[5][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_23_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_23_wr_en             (q_fwd_tbl1_wen[5][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_24_adr               (fwd_tbl1_addr[6][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_24_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_24_rd_en             (q_fwd_tbl1_ren[6][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_24_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_24_wr_en             (q_fwd_tbl1_wen[6][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_25_adr               (fwd_tbl1_addr[6][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_25_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_25_rd_en             (q_fwd_tbl1_ren[6][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_25_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_25_wr_en             (q_fwd_tbl1_wen[6][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_26_adr               (fwd_tbl1_addr[6][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_26_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_26_rd_en             (q_fwd_tbl1_ren[6][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_26_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_26_wr_en             (q_fwd_tbl1_wen[6][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_27_adr               (fwd_tbl1_addr[6][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_27_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_27_rd_en             (q_fwd_tbl1_ren[6][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_27_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_27_wr_en             (q_fwd_tbl1_wen[6][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_28_adr               (fwd_tbl1_addr[7][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_28_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_28_rd_en             (q_fwd_tbl1_ren[7][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_28_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_28_wr_en             (q_fwd_tbl1_wen[7][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_29_adr               (fwd_tbl1_addr[7][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_29_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_29_rd_en             (q_fwd_tbl1_ren[7][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_29_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_29_wr_en             (q_fwd_tbl1_wen[7][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_2_adr                (fwd_tbl1_addr[0][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_2_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_2_rd_en              (q_fwd_tbl1_ren[0][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_2_wr_data            (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_2_wr_en              (q_fwd_tbl1_wen[0][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_30_adr               (fwd_tbl1_addr[7][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_30_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_30_rd_en             (q_fwd_tbl1_ren[7][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_30_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_30_wr_en             (q_fwd_tbl1_wen[7][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_31_adr               (fwd_tbl1_addr[7][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_31_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_31_rd_en             (q_fwd_tbl1_ren[7][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_31_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_31_wr_en             (q_fwd_tbl1_wen[7][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_32_adr               (fwd_tbl1_addr[8][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_32_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_32_rd_en             (q_fwd_tbl1_ren[8][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_32_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_32_wr_en             (q_fwd_tbl1_wen[8][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_33_adr               (fwd_tbl1_addr[8][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_33_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_33_rd_en             (q_fwd_tbl1_ren[8][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_33_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_33_wr_en             (q_fwd_tbl1_wen[8][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_34_adr               (fwd_tbl1_addr[8][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_34_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_34_rd_en             (q_fwd_tbl1_ren[8][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_34_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_34_wr_en             (q_fwd_tbl1_wen[8][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_35_adr               (fwd_tbl1_addr[8][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_35_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_35_rd_en             (q_fwd_tbl1_ren[8][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_35_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_35_wr_en             (q_fwd_tbl1_wen[8][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_36_adr               (fwd_tbl1_addr[9][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_36_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_36_rd_en             (q_fwd_tbl1_ren[9][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_36_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_36_wr_en             (q_fwd_tbl1_wen[9][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_37_adr               (fwd_tbl1_addr[9][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_37_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_37_rd_en             (q_fwd_tbl1_ren[9][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_37_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_37_wr_en             (q_fwd_tbl1_wen[9][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_38_adr               (fwd_tbl1_addr[9][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_38_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_38_rd_en             (q_fwd_tbl1_ren[9][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_38_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_38_wr_en             (q_fwd_tbl1_wen[9][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_39_wr_en             (q_fwd_tbl1_wen[9][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_3_adr                (fwd_tbl1_addr[0][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_3_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_3_rd_en              (q_fwd_tbl1_ren[0][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_3_wr_data            (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_3_wr_en              (q_fwd_tbl1_wen[0][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_40_adr               (fwd_tbl1_addr[10][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_40_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_40_rd_en             (q_fwd_tbl1_ren[10][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_40_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_40_wr_en             (q_fwd_tbl1_wen[10][0]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_41_adr               (fwd_tbl1_addr[10][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_41_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_41_rd_en             (q_fwd_tbl1_ren[10][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_41_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_41_wr_en             (q_fwd_tbl1_wen[10][1]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_42_adr               (fwd_tbl1_addr[10][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_42_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_42_rd_en             (q_fwd_tbl1_ren[10][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_42_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_42_wr_en             (q_fwd_tbl1_wen[10][2]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_43_adr               (fwd_tbl1_addr[10][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_43_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_43_rd_en             (q_fwd_tbl1_ren[10][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_43_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_43_wr_en             (q_fwd_tbl1_wen[10][3]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_44_adr               (fwd_tbl1_addr[11][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_44_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_44_rd_en             (q_fwd_tbl1_ren[11][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_44_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_44_wr_en             (q_fwd_tbl1_wen[11][0]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_45_adr               (fwd_tbl1_addr[11][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_45_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_45_rd_en             (q_fwd_tbl1_ren[11][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_45_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_45_wr_en             (q_fwd_tbl1_wen[11][1]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_46_adr               (fwd_tbl1_addr[11][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_46_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_46_rd_en             (q_fwd_tbl1_ren[11][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_46_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_46_wr_en             (q_fwd_tbl1_wen[11][2]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_47_adr               (fwd_tbl1_addr[11][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_49_rd_en             (q_fwd_tbl1_ren[12][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_49_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_49_wr_en             (q_fwd_tbl1_wen[12][1]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_4_adr                (fwd_tbl1_addr[1][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_4_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_4_rd_en              (q_fwd_tbl1_ren[1][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_4_wr_data            (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_4_wr_en              (q_fwd_tbl1_wen[1][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_50_adr               (fwd_tbl1_addr[12][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_50_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_50_rd_en             (q_fwd_tbl1_ren[12][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_50_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_50_wr_en             (q_fwd_tbl1_wen[12][2]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_51_adr               (fwd_tbl1_addr[12][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_51_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_51_rd_en             (q_fwd_tbl1_ren[12][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_51_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_51_wr_en             (q_fwd_tbl1_wen[12][3]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_52_adr               (fwd_tbl1_addr[13][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_52_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_52_rd_en             (q_fwd_tbl1_ren[13][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_52_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_52_wr_en             (q_fwd_tbl1_wen[13][0]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_53_adr               (fwd_tbl1_addr[13][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_53_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_53_rd_en             (q_fwd_tbl1_ren[13][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_53_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_54_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_54_wr_en             (q_fwd_tbl1_wen[13][2]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_55_adr               (fwd_tbl1_addr[13][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_55_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_55_rd_en             (q_fwd_tbl1_ren[13][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_55_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_55_wr_en             (q_fwd_tbl1_wen[13][3]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_56_adr               (fwd_tbl1_addr[14][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_56_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_56_rd_en             (q_fwd_tbl1_ren[14][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_56_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_56_wr_en             (q_fwd_tbl1_wen[14][0]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_57_adr               (fwd_tbl1_addr[14][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_57_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_57_rd_en             (q_fwd_tbl1_ren[14][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_57_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_57_wr_en             (q_fwd_tbl1_wen[14][1]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_58_adr               (fwd_tbl1_addr[14][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_58_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_58_rd_en             (q_fwd_tbl1_ren[14][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_58_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_58_wr_en             (q_fwd_tbl1_wen[14][2]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_59_adr               (fwd_tbl1_addr[14][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_59_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_59_rd_en             (q_fwd_tbl1_ren[14][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_59_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_59_wr_en             (q_fwd_tbl1_wen[14][3]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_5_adr                (fwd_tbl1_addr[1][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_5_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_5_rd_en              (q_fwd_tbl1_ren[1][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_5_wr_data            (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_5_wr_en              (q_fwd_tbl1_wen[1][1]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_60_adr               (fwd_tbl1_addr[15][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_60_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_60_rd_en             (q_fwd_tbl1_ren[15][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_60_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_60_wr_en             (q_fwd_tbl1_wen[15][0]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_61_adr               (fwd_tbl1_addr[15][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_61_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_61_rd_en             (q_fwd_tbl1_ren[15][1]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_61_wr_data           (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_61_wr_en             (q_fwd_tbl1_wen[15][1]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_62_adr               (fwd_tbl1_addr[15][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_62_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_62_rd_en             (q_fwd_tbl1_ren[15][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_62_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_62_wr_en             (q_fwd_tbl1_wen[15][2]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_63_adr               (fwd_tbl1_addr[15][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_63_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_63_rd_en             (q_fwd_tbl1_ren[15][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_63_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_63_wr_en             (q_fwd_tbl1_wen[15][3]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_6_adr                (fwd_tbl1_addr[1][2]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_6_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_6_rd_en              (q_fwd_tbl1_ren[1][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_6_wr_data            (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_6_wr_en              (q_fwd_tbl1_wen[1][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_7_adr                (fwd_tbl1_addr[1][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_7_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_7_rd_en              (q_fwd_tbl1_ren[1][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_7_wr_data            (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_7_wr_en              (q_fwd_tbl1_wen[1][3]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_8_adr                (fwd_tbl1_addr[2][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_8_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_8_rd_en              (q_fwd_tbl1_ren[2][0]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_8_wr_data            (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_8_wr_en              (q_fwd_tbl1_wen[2][0]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_9_adr                (fwd_tbl1_addr[2][1]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_9_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_9_rd_en              (q_fwd_tbl1_ren[2][1]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_9_wr_data            (q_fwd_tbl1_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_9_wr_en              (q_fwd_tbl1_wen[2][1]),                            
/* input  logic   [11:0] */ .ppe_stm_l3mc_tbl_adr                  (),                                                
/* input  logic          */ .ppe_stm_l3mc_tbl_mem_ls_enter         (),                                                
/* input  logic          */ .ppe_stm_l3mc_tbl_rd_en                (),                                                
/* input  logic  [511:0] */ .ppe_stm_l3mc_tbl_wr_data              (),                                                
/* input  logic          */ .ppe_stm_l3mc_tbl_wr_en                (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_0_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_0_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_0_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_0_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_0_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_10_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_10_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_10_rd_en              (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_11_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_11_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_11_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_11_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_12_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_12_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_12_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_12_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_12_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_13_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_13_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_13_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_13_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_13_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_14_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_14_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_14_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_14_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_14_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_15_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_15_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_15_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_15_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_15_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_16_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_16_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_16_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_16_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_16_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_17_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_17_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_17_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_17_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_17_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_18_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_18_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_18_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_18_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_18_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_19_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_19_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_19_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_19_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_19_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_1_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_1_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_1_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_1_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_1_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_20_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_20_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_20_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_20_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_20_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_21_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_21_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_21_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_21_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_21_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_22_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_22_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_22_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_22_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_22_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_23_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_23_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_23_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_23_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_23_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_24_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_28_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_29_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_29_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_29_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_29_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_29_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_2_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_2_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_2_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_2_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_2_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_30_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_30_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_30_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_30_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_30_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_31_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_31_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_31_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_31_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_31_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_32_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_32_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_32_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_32_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_32_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_33_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_33_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_33_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_33_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_33_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_34_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_34_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_34_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_34_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_34_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_35_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_35_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_35_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_35_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_35_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_36_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_36_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_36_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_36_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_36_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_37_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_37_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_37_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_37_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_37_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_38_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_38_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_38_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_38_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_38_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_39_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_39_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_39_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_39_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_39_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_3_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_3_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_3_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_3_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_3_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_40_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_40_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_40_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_40_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_40_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_41_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_41_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_41_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_41_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_41_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_42_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_42_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_42_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_42_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_42_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_43_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_43_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_43_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_43_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_43_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_44_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_44_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_44_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_44_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_44_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_45_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_45_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_45_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_45_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_45_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_46_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_46_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_46_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_46_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_46_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_47_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_47_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_47_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_47_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_47_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_48_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_48_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_48_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_48_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_48_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_49_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_49_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_49_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_49_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_49_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_4_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_4_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_4_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_4_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_4_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_50_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_50_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_50_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_50_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_50_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_51_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_51_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_51_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_51_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_51_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_52_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_52_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_52_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_52_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_52_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_53_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_53_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_53_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_53_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_53_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_54_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_54_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_54_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_54_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_54_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_55_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_55_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_55_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_55_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_55_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_56_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_56_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_56_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_56_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_56_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_57_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_57_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_57_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_57_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_57_wr_en              (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_58_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_59_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_59_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_59_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_59_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_59_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_5_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_5_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_5_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_5_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_5_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_60_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_60_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_60_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_60_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_60_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_61_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_61_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_61_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_61_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_61_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_62_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_62_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_62_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_62_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_62_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_63_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_63_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_63_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_63_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_63_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_64_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_64_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_64_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_64_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_64_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_65_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_65_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_65_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_65_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_65_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_66_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_66_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_66_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_66_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_66_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_67_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_67_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_67_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_67_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_67_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_68_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_68_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_68_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_68_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_68_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_69_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_69_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_69_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_69_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_69_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_6_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_6_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_6_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_6_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_6_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_70_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_70_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_70_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_70_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_70_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_71_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_71_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_71_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_71_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_71_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_72_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_72_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_72_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_72_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_72_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_73_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_73_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_73_rd_en              (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_74_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_74_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_74_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_75_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_75_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_75_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_75_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_75_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_76_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_76_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_76_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_76_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_76_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_77_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_77_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_77_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_77_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_77_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_78_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_78_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_78_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_78_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_78_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_79_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_79_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_79_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_79_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_79_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_7_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_7_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_7_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_7_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_7_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_8_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_8_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_8_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_8_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_8_wr_en               (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_9_adr                 (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_9_mem_ls_enter        (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_9_rd_en               (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_9_wr_data             (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_9_wr_en               (),                                                
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_0_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_0_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_100_from_mem (ppe_stm_ppe_stm_fwd_tbl0_100_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_101_from_mem (ppe_stm_ppe_stm_fwd_tbl0_101_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_102_from_mem (ppe_stm_ppe_stm_fwd_tbl0_102_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_103_from_mem (ppe_stm_ppe_stm_fwd_tbl0_103_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_104_from_mem (ppe_stm_ppe_stm_fwd_tbl0_104_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_105_from_mem (ppe_stm_ppe_stm_fwd_tbl0_105_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_106_from_mem (ppe_stm_ppe_stm_fwd_tbl0_106_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_107_from_mem (ppe_stm_ppe_stm_fwd_tbl0_107_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_108_from_mem (ppe_stm_ppe_stm_fwd_tbl0_108_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_109_from_mem (ppe_stm_ppe_stm_fwd_tbl0_109_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_10_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_10_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_110_from_mem (ppe_stm_ppe_stm_fwd_tbl0_110_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_111_from_mem (ppe_stm_ppe_stm_fwd_tbl0_111_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_112_from_mem (ppe_stm_ppe_stm_fwd_tbl0_112_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_113_from_mem (ppe_stm_ppe_stm_fwd_tbl0_113_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_114_from_mem (ppe_stm_ppe_stm_fwd_tbl0_114_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_115_from_mem (ppe_stm_ppe_stm_fwd_tbl0_115_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_116_from_mem (ppe_stm_ppe_stm_fwd_tbl0_116_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_117_from_mem (ppe_stm_ppe_stm_fwd_tbl0_117_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_118_from_mem (ppe_stm_ppe_stm_fwd_tbl0_118_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_119_from_mem (ppe_stm_ppe_stm_fwd_tbl0_119_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_11_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_11_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_120_from_mem (ppe_stm_ppe_stm_fwd_tbl0_120_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_121_from_mem (ppe_stm_ppe_stm_fwd_tbl0_121_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_122_from_mem (ppe_stm_ppe_stm_fwd_tbl0_122_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_123_from_mem (ppe_stm_ppe_stm_fwd_tbl0_123_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_124_from_mem (ppe_stm_ppe_stm_fwd_tbl0_124_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_125_from_mem (ppe_stm_ppe_stm_fwd_tbl0_125_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_126_from_mem (ppe_stm_ppe_stm_fwd_tbl0_126_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_127_from_mem (ppe_stm_ppe_stm_fwd_tbl0_127_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_128_from_mem (ppe_stm_ppe_stm_fwd_tbl0_128_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_129_from_mem (ppe_stm_ppe_stm_fwd_tbl0_129_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_12_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_12_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_130_from_mem (ppe_stm_ppe_stm_fwd_tbl0_130_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_131_from_mem (ppe_stm_ppe_stm_fwd_tbl0_131_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_132_from_mem (ppe_stm_ppe_stm_fwd_tbl0_132_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_133_from_mem (ppe_stm_ppe_stm_fwd_tbl0_133_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_134_from_mem (ppe_stm_ppe_stm_fwd_tbl0_134_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_135_from_mem (ppe_stm_ppe_stm_fwd_tbl0_135_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_136_from_mem (ppe_stm_ppe_stm_fwd_tbl0_136_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_137_from_mem (ppe_stm_ppe_stm_fwd_tbl0_137_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_138_from_mem (ppe_stm_ppe_stm_fwd_tbl0_138_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_139_from_mem (ppe_stm_ppe_stm_fwd_tbl0_139_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_13_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_13_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_140_from_mem (ppe_stm_ppe_stm_fwd_tbl0_140_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_141_from_mem (ppe_stm_ppe_stm_fwd_tbl0_141_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_142_from_mem (ppe_stm_ppe_stm_fwd_tbl0_142_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_143_from_mem (ppe_stm_ppe_stm_fwd_tbl0_143_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_144_from_mem (ppe_stm_ppe_stm_fwd_tbl0_144_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_145_from_mem (ppe_stm_ppe_stm_fwd_tbl0_145_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_146_from_mem (ppe_stm_ppe_stm_fwd_tbl0_146_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_147_from_mem (ppe_stm_ppe_stm_fwd_tbl0_147_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_148_from_mem (ppe_stm_ppe_stm_fwd_tbl0_148_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_149_from_mem (ppe_stm_ppe_stm_fwd_tbl0_149_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_14_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_14_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_150_from_mem (ppe_stm_ppe_stm_fwd_tbl0_150_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_155_from_mem (ppe_stm_ppe_stm_fwd_tbl0_155_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_156_from_mem (ppe_stm_ppe_stm_fwd_tbl0_156_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_157_from_mem (ppe_stm_ppe_stm_fwd_tbl0_157_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_158_from_mem (ppe_stm_ppe_stm_fwd_tbl0_158_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_159_from_mem (ppe_stm_ppe_stm_fwd_tbl0_159_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_15_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_15_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_160_from_mem (ppe_stm_ppe_stm_fwd_tbl0_160_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_161_from_mem (ppe_stm_ppe_stm_fwd_tbl0_161_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_162_from_mem (ppe_stm_ppe_stm_fwd_tbl0_162_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_163_from_mem (ppe_stm_ppe_stm_fwd_tbl0_163_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_164_from_mem (ppe_stm_ppe_stm_fwd_tbl0_164_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_165_from_mem (ppe_stm_ppe_stm_fwd_tbl0_165_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_166_from_mem (ppe_stm_ppe_stm_fwd_tbl0_166_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_167_from_mem (ppe_stm_ppe_stm_fwd_tbl0_167_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_168_from_mem (ppe_stm_ppe_stm_fwd_tbl0_168_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_169_from_mem (ppe_stm_ppe_stm_fwd_tbl0_169_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_16_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_16_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_170_from_mem (ppe_stm_ppe_stm_fwd_tbl0_170_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_171_from_mem (ppe_stm_ppe_stm_fwd_tbl0_171_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_172_from_mem (ppe_stm_ppe_stm_fwd_tbl0_172_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_173_from_mem (ppe_stm_ppe_stm_fwd_tbl0_173_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_174_from_mem (ppe_stm_ppe_stm_fwd_tbl0_174_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_175_from_mem (ppe_stm_ppe_stm_fwd_tbl0_175_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_176_from_mem (ppe_stm_ppe_stm_fwd_tbl0_176_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_177_from_mem (ppe_stm_ppe_stm_fwd_tbl0_177_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_178_from_mem (ppe_stm_ppe_stm_fwd_tbl0_178_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_179_from_mem (ppe_stm_ppe_stm_fwd_tbl0_179_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_17_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_17_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_180_from_mem (ppe_stm_ppe_stm_fwd_tbl0_180_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_181_from_mem (ppe_stm_ppe_stm_fwd_tbl0_181_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_182_from_mem (ppe_stm_ppe_stm_fwd_tbl0_182_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_183_from_mem (ppe_stm_ppe_stm_fwd_tbl0_183_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_184_from_mem (ppe_stm_ppe_stm_fwd_tbl0_184_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_185_from_mem (ppe_stm_ppe_stm_fwd_tbl0_185_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_186_from_mem (ppe_stm_ppe_stm_fwd_tbl0_186_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_187_from_mem (ppe_stm_ppe_stm_fwd_tbl0_187_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_188_from_mem (ppe_stm_ppe_stm_fwd_tbl0_188_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_189_from_mem (ppe_stm_ppe_stm_fwd_tbl0_189_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_18_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_18_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_190_from_mem (ppe_stm_ppe_stm_fwd_tbl0_190_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_191_from_mem (ppe_stm_ppe_stm_fwd_tbl0_191_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_19_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_19_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_1_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_1_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_20_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_20_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_21_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_21_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_22_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_22_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_23_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_23_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_24_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_24_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_25_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_25_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_26_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_26_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_27_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_27_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_28_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_28_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_29_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_29_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_2_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_2_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_30_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_30_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_31_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_31_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_32_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_32_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_33_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_33_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_34_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_34_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_35_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_35_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_36_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_36_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_37_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_37_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_38_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_38_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_39_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_39_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_3_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_3_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_40_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_40_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_41_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_41_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_42_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_42_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_43_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_43_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_44_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_44_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_45_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_45_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_46_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_46_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_47_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_47_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_48_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_48_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_49_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_49_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_4_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_4_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_50_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_50_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_51_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_51_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_52_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_52_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_53_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_53_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_54_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_54_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_55_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_55_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_56_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_56_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_57_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_57_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_58_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_58_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_59_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_59_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_5_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_5_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_60_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_60_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_61_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_61_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_62_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_62_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_63_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_63_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_64_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_64_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_65_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_65_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_66_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_66_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_67_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_67_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_68_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_68_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_69_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_69_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_6_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_6_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_70_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_70_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_71_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_71_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_72_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_72_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_73_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_73_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_74_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_74_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_75_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_75_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_76_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_76_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_77_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_77_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_78_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_78_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_79_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_79_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_7_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_7_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_80_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_80_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_81_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_81_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_82_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_82_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_83_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_83_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_84_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_84_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_85_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_85_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_86_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_86_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_87_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_87_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_88_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_88_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_89_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_89_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_8_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_8_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_90_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_90_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_91_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_91_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_92_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_92_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_97_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_97_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_98_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_98_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_99_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_99_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_9_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_9_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_0_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_0_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_10_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_10_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_11_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_11_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_12_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_12_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_13_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_13_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_14_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_14_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_15_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_15_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_16_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_16_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_17_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_17_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_18_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_18_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_19_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_19_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_1_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_1_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_20_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_20_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_21_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_21_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_22_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_22_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_23_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_23_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_24_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_24_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_25_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_25_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_26_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_26_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_27_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_27_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_28_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_28_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_29_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_29_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_2_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_2_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_30_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_30_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_31_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_31_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_32_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_32_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_33_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_33_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_34_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_34_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_35_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_35_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_36_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_36_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_37_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_37_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_38_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_38_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_39_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_39_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_3_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_3_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_40_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_40_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_41_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_41_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_42_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_42_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_43_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_43_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_44_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_44_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_45_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_45_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_46_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_46_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_47_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_47_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_48_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_48_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_49_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_49_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_4_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_4_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_50_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_50_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_51_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_51_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_52_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_52_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_53_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_53_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_54_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_54_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_55_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_55_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_56_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_56_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_57_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_57_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_58_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_58_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_59_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_59_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_5_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_5_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_60_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_60_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_61_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_61_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_62_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_62_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_63_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_63_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_6_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_6_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_7_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_7_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_8_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_8_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_9_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_9_from_mem),             
/* input  logic  [576:0] */ .ppe_stm_ppe_stm_l3mc_tbl_from_mem     (ppe_stm_ppe_stm_l3mc_tbl_from_mem),               
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_0_from_mem    (ppe_stm_ppe_stm_mod_tbl_0_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_10_from_mem   (ppe_stm_ppe_stm_mod_tbl_10_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_11_from_mem   (ppe_stm_ppe_stm_mod_tbl_11_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_12_from_mem   (ppe_stm_ppe_stm_mod_tbl_12_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_13_from_mem   (ppe_stm_ppe_stm_mod_tbl_13_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_14_from_mem   (ppe_stm_ppe_stm_mod_tbl_14_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_15_from_mem   (ppe_stm_ppe_stm_mod_tbl_15_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_16_from_mem   (ppe_stm_ppe_stm_mod_tbl_16_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_17_from_mem   (ppe_stm_ppe_stm_mod_tbl_17_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_18_from_mem   (ppe_stm_ppe_stm_mod_tbl_18_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_19_from_mem   (ppe_stm_ppe_stm_mod_tbl_19_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_1_from_mem    (ppe_stm_ppe_stm_mod_tbl_1_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_20_from_mem   (ppe_stm_ppe_stm_mod_tbl_20_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_21_from_mem   (ppe_stm_ppe_stm_mod_tbl_21_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_22_from_mem   (ppe_stm_ppe_stm_mod_tbl_22_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_23_from_mem   (ppe_stm_ppe_stm_mod_tbl_23_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_24_from_mem   (ppe_stm_ppe_stm_mod_tbl_24_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_25_from_mem   (ppe_stm_ppe_stm_mod_tbl_25_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_26_from_mem   (ppe_stm_ppe_stm_mod_tbl_26_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_27_from_mem   (ppe_stm_ppe_stm_mod_tbl_27_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_28_from_mem   (ppe_stm_ppe_stm_mod_tbl_28_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_29_from_mem   (ppe_stm_ppe_stm_mod_tbl_29_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_2_from_mem    (ppe_stm_ppe_stm_mod_tbl_2_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_30_from_mem   (ppe_stm_ppe_stm_mod_tbl_30_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_31_from_mem   (ppe_stm_ppe_stm_mod_tbl_31_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_32_from_mem   (ppe_stm_ppe_stm_mod_tbl_32_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_33_from_mem   (ppe_stm_ppe_stm_mod_tbl_33_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_34_from_mem   (ppe_stm_ppe_stm_mod_tbl_34_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_35_from_mem   (ppe_stm_ppe_stm_mod_tbl_35_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_36_from_mem   (ppe_stm_ppe_stm_mod_tbl_36_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_37_from_mem   (ppe_stm_ppe_stm_mod_tbl_37_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_38_from_mem   (ppe_stm_ppe_stm_mod_tbl_38_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_39_from_mem   (ppe_stm_ppe_stm_mod_tbl_39_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_3_from_mem    (ppe_stm_ppe_stm_mod_tbl_3_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_40_from_mem   (ppe_stm_ppe_stm_mod_tbl_40_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_41_from_mem   (ppe_stm_ppe_stm_mod_tbl_41_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_42_from_mem   (ppe_stm_ppe_stm_mod_tbl_42_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_43_from_mem   (ppe_stm_ppe_stm_mod_tbl_43_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_44_from_mem   (ppe_stm_ppe_stm_mod_tbl_44_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_45_from_mem   (ppe_stm_ppe_stm_mod_tbl_45_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_46_from_mem   (ppe_stm_ppe_stm_mod_tbl_46_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_47_from_mem   (ppe_stm_ppe_stm_mod_tbl_47_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_48_from_mem   (ppe_stm_ppe_stm_mod_tbl_48_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_49_from_mem   (ppe_stm_ppe_stm_mod_tbl_49_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_4_from_mem    (ppe_stm_ppe_stm_mod_tbl_4_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_50_from_mem   (ppe_stm_ppe_stm_mod_tbl_50_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_51_from_mem   (ppe_stm_ppe_stm_mod_tbl_51_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_52_from_mem   (ppe_stm_ppe_stm_mod_tbl_52_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_53_from_mem   (ppe_stm_ppe_stm_mod_tbl_53_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_54_from_mem   (ppe_stm_ppe_stm_mod_tbl_54_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_55_from_mem   (ppe_stm_ppe_stm_mod_tbl_55_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_56_from_mem   (ppe_stm_ppe_stm_mod_tbl_56_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_57_from_mem   (ppe_stm_ppe_stm_mod_tbl_57_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_61_from_mem   (ppe_stm_ppe_stm_mod_tbl_61_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_62_from_mem   (ppe_stm_ppe_stm_mod_tbl_62_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_63_from_mem   (ppe_stm_ppe_stm_mod_tbl_63_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_64_from_mem   (ppe_stm_ppe_stm_mod_tbl_64_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_65_from_mem   (ppe_stm_ppe_stm_mod_tbl_65_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_66_from_mem   (ppe_stm_ppe_stm_mod_tbl_66_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_67_from_mem   (ppe_stm_ppe_stm_mod_tbl_67_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_68_from_mem   (ppe_stm_ppe_stm_mod_tbl_68_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_69_from_mem   (ppe_stm_ppe_stm_mod_tbl_69_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_6_from_mem    (ppe_stm_ppe_stm_mod_tbl_6_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_70_from_mem   (ppe_stm_ppe_stm_mod_tbl_70_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_71_from_mem   (ppe_stm_ppe_stm_mod_tbl_71_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_72_from_mem   (ppe_stm_ppe_stm_mod_tbl_72_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_73_from_mem   (ppe_stm_ppe_stm_mod_tbl_73_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_74_from_mem   (ppe_stm_ppe_stm_mod_tbl_74_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_75_from_mem   (ppe_stm_ppe_stm_mod_tbl_75_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_76_from_mem   (ppe_stm_ppe_stm_mod_tbl_76_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_77_from_mem   (ppe_stm_ppe_stm_mod_tbl_77_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_78_from_mem   (ppe_stm_ppe_stm_mod_tbl_78_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_79_from_mem   (ppe_stm_ppe_stm_mod_tbl_79_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_7_from_mem    (ppe_stm_ppe_stm_mod_tbl_7_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_8_from_mem    (ppe_stm_ppe_stm_mod_tbl_8_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_9_from_mem    (ppe_stm_ppe_stm_mod_tbl_9_from_mem),              
/* input  logic   [40:0] */ .ppe_stm_ppe_stm_shcp_tbl_from_mem     (ppe_stm_ppe_stm_shcp_tbl_from_mem),               
/* input  logic   [14:0] */ .ppe_stm_shcp_tbl_adr                  (),                                                
/* input  logic          */ .ppe_stm_shcp_tbl_mem_ls_enter         (),                                                
/* input  logic          */ .ppe_stm_shcp_tbl_rd_en                (),                                                
/* input  logic   [32:0] */ .ppe_stm_shcp_tbl_wr_data              (),                                                
/* input  logic          */ .ppe_stm_shcp_tbl_wr_en                (),                                                
/* input  logic          */ .reset_n                               (reset_n),                                         
/* input  logic          */ .unified_regs_rd                       (),                                                
/* input  logic   [31:0] */ .unified_regs_wr_data                  (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_47_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_47_rd_en             (q_fwd_tbl1_ren[11][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_47_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_47_wr_en             (q_fwd_tbl1_wen[11][3]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_48_adr               (fwd_tbl1_addr[12][0]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_48_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_48_rd_en             (q_fwd_tbl1_ren[12][0]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_48_wr_data           (q_fwd_tbl1_wdata[0][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_48_wr_en             (q_fwd_tbl1_wen[12][0]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_49_adr               (fwd_tbl1_addr[12][1]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_49_mem_ls_enter      (),                                                
/* input  logic          */ .PPE_STM_ECC_COR_ERR_reg_sel           (),                                                
/* input  logic          */ .PPE_STM_ECC_UNCOR_ERR_reg_sel         (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_0_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_0_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_100_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_100_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_101_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_101_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_102_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_SHCP_TBL_STATUS_reg_sel       (),                                                
/* input  logic          */ .clk                                   (cclk),                                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_0_adr                (fwd_tbl0_addr[0][0]),                             
/* input  logic          */ .ppe_stm_fwd_tbl0_0_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_115_rd_en            (q_fwd_tbl0_ren[28][3]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_115_wr_data          (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_115_wr_en            (q_fwd_tbl0_wen[28][3]),                           
/* input  logic          */ .PPE_STM_FWD_TBL0_170_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_171_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_171_STATUS_reg_sel   (),                                                
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_177_wr_data          (q_fwd_tbl0_wdata[1][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_177_wr_en            (q_fwd_tbl0_wen[44][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_178_adr              (fwd_tbl0_addr[44][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_178_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_22_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_22_rd_en             (q_fwd_tbl1_ren[5][2]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_22_wr_data           (q_fwd_tbl1_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl1_22_wr_en             (q_fwd_tbl1_wen[5][2]),                            
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_39_adr               (fwd_tbl1_addr[9][3]),                             
/* input  logic          */ .ppe_stm_fwd_tbl1_39_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_39_rd_en             (q_fwd_tbl1_ren[9][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl1_39_wr_data           (q_fwd_tbl1_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_mod_tbl_27_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_27_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_27_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_27_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_28_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_28_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_28_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_28_wr_data            (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_98_rd_en             (q_fwd_tbl0_ren[24][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_98_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_98_wr_en             (q_fwd_tbl0_wen[24][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_99_adr               (fwd_tbl0_addr[24][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_53_wr_en             (q_fwd_tbl1_wen[13][1]),                           
/* input  logic   [10:0] */ .ppe_stm_fwd_tbl1_54_adr               (fwd_tbl1_addr[13][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl1_54_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl1_54_rd_en             (q_fwd_tbl1_ren[13][2]),                           
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_10_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_10_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_11_adr                (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_58_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_58_mem_ls_enter       (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_58_rd_en              (),                                                
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_58_wr_data            (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_104_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_105_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_105_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_106_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_106_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_107_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_107_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_108_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_108_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_109_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_109_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_10_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_10_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_110_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_110_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_37_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_38_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_38_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_39_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_75_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_76_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_76_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_77_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_25_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_25_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_26_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_26_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_63_CFG_reg_sel       (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_63_STATUS_reg_sel    (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_6_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL1_6_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_44_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_45_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_45_STATUS_reg_sel     (),                                                
/* input  logic          */ .PPE_STM_MOD_TBL_46_CFG_reg_sel        (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_102_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_103_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_103_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_104_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_132_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_132_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_133_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_133_STATUS_reg_sel   (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_35_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_35_rd_en             (q_fwd_tbl0_ren[8][3]),                            
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_35_wr_data           (q_fwd_tbl0_wdata[3][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_35_wr_en             (q_fwd_tbl0_wen[8][3]),                            
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_51_adr               (fwd_tbl0_addr[12][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_51_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_51_rd_en             (q_fwd_tbl0_ren[12][3]),                           
/* input  logic          */ .ppe_stm_fwd_tbl0_146_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_146_rd_en            (q_fwd_tbl0_ren[36][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_146_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_161_wr_en            (q_fwd_tbl0_wen[40][1]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_162_adr              (fwd_tbl0_addr[40][2]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_162_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_162_rd_en            (q_fwd_tbl0_ren[40][2]),                           
/* input  logic          */ .ppe_stm_fwd_tbl0_130_mem_ls_enter     (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_130_rd_en            (q_fwd_tbl0_ren[32][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_130_wr_data          (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_130_wr_en            (q_fwd_tbl0_wen[32][2]),                           
/* input  logic   [63:0] */ .ppe_stm_mod_tbl_73_wr_data            (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_73_wr_en              (),                                                
/* input  logic   [10:0] */ .ppe_stm_mod_tbl_74_adr                (),                                                
/* input  logic          */ .ppe_stm_mod_tbl_74_mem_ls_enter       (),                                                
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_151_from_mem (ppe_stm_ppe_stm_fwd_tbl0_151_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_152_from_mem (ppe_stm_ppe_stm_fwd_tbl0_152_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_153_from_mem (ppe_stm_ppe_stm_fwd_tbl0_153_from_mem),           
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_154_from_mem (ppe_stm_ppe_stm_fwd_tbl0_154_from_mem),           
/* input  logic          */ .ppe_stm_fwd_tbl0_66_wr_en             (q_fwd_tbl0_wen[16][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_67_adr               (fwd_tbl0_addr[16][3]),                            
/* input  logic          */ .ppe_stm_fwd_tbl0_67_mem_ls_enter      (),                                                
/* input  logic          */ .ppe_stm_fwd_tbl0_67_rd_en             (q_fwd_tbl0_ren[16][3]),                           
/* input  logic          */ .ppe_stm_fwd_tbl0_82_rd_en             (q_fwd_tbl0_ren[20][2]),                           
/* input  logic   [71:0] */ .ppe_stm_fwd_tbl0_82_wr_data           (q_fwd_tbl0_wdata[2][71:0]),                       
/* input  logic          */ .ppe_stm_fwd_tbl0_82_wr_en             (q_fwd_tbl0_wen[20][2]),                           
/* input  logic   [11:0] */ .ppe_stm_fwd_tbl0_83_adr               (fwd_tbl0_addr[20][3]),                            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_93_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_93_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_94_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_94_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_95_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_95_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_96_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_96_from_mem),            
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_58_from_mem   (ppe_stm_ppe_stm_mod_tbl_58_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_59_from_mem   (ppe_stm_ppe_stm_mod_tbl_59_from_mem),             
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_5_from_mem    (ppe_stm_ppe_stm_mod_tbl_5_from_mem),              
/* input  logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_60_from_mem   (ppe_stm_ppe_stm_mod_tbl_60_from_mem),             
/* input  logic          */ .PPE_STM_FWD_TBL0_111_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_111_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_112_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_112_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_113_CFG_reg_sel      (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_113_STATUS_reg_sel   (),                                                
/* input  logic          */ .PPE_STM_FWD_TBL0_114_CFG_reg_sel      (),                                                
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_132_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_132_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_133_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_133_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_134_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_134_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_135_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_135_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_136_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_136_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_137_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_137_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_138_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_138_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_139_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_139_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_13_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_13_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_140_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_140_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_141_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_141_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_142_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_142_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_143_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_143_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_144_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_144_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_145_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_145_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_146_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_146_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_147_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_147_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_148_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_148_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_149_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_149_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_14_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_14_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_150_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_150_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_151_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_151_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_152_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_152_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_153_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_153_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_154_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_154_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_155_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_155_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_156_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_156_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_157_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_157_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_158_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_158_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_159_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_159_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_15_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_15_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_160_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_160_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_161_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_161_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_162_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_162_to_mem),             
/* output logic          */ .ppe_stm_ecc_int                       (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_0_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_0_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_0_rd_data            (fwd_tbl0_rdata[0][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_0_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_100_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_100_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_100_rd_data          (fwd_tbl0_rdata[25][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_100_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_101_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_101_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_101_rd_data          (fwd_tbl0_rdata[25][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_101_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_102_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_102_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_102_rd_data          (fwd_tbl0_rdata[25][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_102_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_103_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_103_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_103_rd_data          (fwd_tbl0_rdata[25][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_103_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_104_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_104_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_104_rd_data          (fwd_tbl0_rdata[26][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_104_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_105_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_105_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_105_rd_data          (fwd_tbl0_rdata[26][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_105_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_106_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_106_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_106_rd_data          (fwd_tbl0_rdata[26][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_106_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_107_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_107_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_107_rd_data          (fwd_tbl0_rdata[26][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_107_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_108_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_108_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_108_rd_data          (fwd_tbl0_rdata[27][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_108_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_109_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_109_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_109_rd_data          (fwd_tbl0_rdata[27][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_109_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_10_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_10_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_10_rd_data           (fwd_tbl0_rdata[2][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_10_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_110_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_110_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_110_rd_data          (fwd_tbl0_rdata[27][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_110_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_111_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_111_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_111_rd_data          (fwd_tbl0_rdata[27][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_111_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_112_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_112_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_112_rd_data          (fwd_tbl0_rdata[28][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_113_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_114_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_114_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_114_rd_data          (fwd_tbl0_rdata[28][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_114_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_115_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_115_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_115_rd_data          (fwd_tbl0_rdata[28][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_115_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_116_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_116_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_116_rd_data          (fwd_tbl0_rdata[29][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_116_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_117_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_117_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_117_rd_data          (fwd_tbl0_rdata[29][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_117_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_118_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_118_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_118_rd_data          (fwd_tbl0_rdata[29][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_118_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_119_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_119_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_119_rd_data          (fwd_tbl0_rdata[29][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_119_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_11_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_11_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_11_rd_data           (fwd_tbl0_rdata[2][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_11_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_120_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_120_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_120_rd_data          (fwd_tbl0_rdata[30][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_120_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_121_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_121_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_121_rd_data          (fwd_tbl0_rdata[30][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_121_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_122_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_122_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_122_rd_data          (fwd_tbl0_rdata[30][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_122_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_123_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_123_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_123_rd_data          (fwd_tbl0_rdata[30][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_123_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_124_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_124_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_124_rd_data          (fwd_tbl0_rdata[31][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_124_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_125_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_125_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_125_rd_data          (fwd_tbl0_rdata[31][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_125_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_126_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_126_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_126_rd_data          (fwd_tbl0_rdata[31][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_126_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_127_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_127_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_127_rd_data          (fwd_tbl0_rdata[31][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_127_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_128_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_128_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_128_rd_data          (fwd_tbl0_rdata[32][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_128_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_129_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_129_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_129_rd_data          (fwd_tbl0_rdata[32][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_129_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_12_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_12_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_12_rd_data           (fwd_tbl0_rdata[3][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_12_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_130_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_130_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_130_rd_data          (fwd_tbl0_rdata[32][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_130_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_131_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_131_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_131_rd_data          (fwd_tbl0_rdata[32][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_131_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_132_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_132_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_132_rd_data          (fwd_tbl0_rdata[33][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_132_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_134_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_134_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_134_rd_data          (fwd_tbl0_rdata[33][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_134_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_135_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_135_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_135_rd_data          (fwd_tbl0_rdata[33][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_135_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_136_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_136_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_136_rd_data          (fwd_tbl0_rdata[34][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_136_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_137_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_137_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_137_rd_data          (fwd_tbl0_rdata[34][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_137_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_138_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_138_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_138_rd_data          (fwd_tbl0_rdata[34][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_138_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_139_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_139_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_139_rd_data          (fwd_tbl0_rdata[34][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_139_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_13_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_13_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_13_rd_data           (fwd_tbl0_rdata[3][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_13_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_140_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_140_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_140_rd_data          (fwd_tbl0_rdata[35][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_140_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_141_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_141_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_141_rd_data          (fwd_tbl0_rdata[35][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_141_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_142_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_142_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_142_rd_data          (fwd_tbl0_rdata[35][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_142_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_143_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_143_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_143_rd_data          (fwd_tbl0_rdata[35][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_143_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_144_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_144_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_144_rd_data          (fwd_tbl0_rdata[36][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_144_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_145_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_145_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_145_rd_data          (fwd_tbl0_rdata[36][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_145_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_146_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_146_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_146_rd_data          (fwd_tbl0_rdata[36][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_146_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_147_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_147_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_147_rd_data          (fwd_tbl0_rdata[36][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_147_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_148_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_148_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_148_rd_data          (fwd_tbl0_rdata[37][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_148_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_149_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_149_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_149_rd_data          (fwd_tbl0_rdata[37][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_149_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_14_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_14_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_14_rd_data           (fwd_tbl0_rdata[3][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_14_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_150_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_150_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_150_rd_data          (fwd_tbl0_rdata[37][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_150_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_151_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_151_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_151_rd_data          (fwd_tbl0_rdata[37][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_151_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_153_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_153_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_153_rd_data          (fwd_tbl0_rdata[38][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_153_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_154_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_154_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_154_rd_data          (fwd_tbl0_rdata[38][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_154_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_155_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_155_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_155_rd_data          (fwd_tbl0_rdata[38][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_155_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_156_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_156_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_156_rd_data          (fwd_tbl0_rdata[39][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_156_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_157_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_157_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_157_rd_data          (fwd_tbl0_rdata[39][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_157_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_158_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_158_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_158_rd_data          (fwd_tbl0_rdata[39][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_158_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_159_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_159_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_159_rd_data          (fwd_tbl0_rdata[39][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_159_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_15_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_15_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_15_rd_data           (fwd_tbl0_rdata[3][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_15_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_160_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_160_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_160_rd_data          (fwd_tbl0_rdata[40][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_160_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_161_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_161_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_161_rd_data          (fwd_tbl0_rdata[40][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_161_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_162_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_162_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_162_rd_data          (fwd_tbl0_rdata[40][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_162_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_163_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_163_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_163_rd_data          (fwd_tbl0_rdata[40][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_163_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_164_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_164_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_164_rd_data          (fwd_tbl0_rdata[41][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_164_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_165_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_165_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_165_rd_data          (fwd_tbl0_rdata[41][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_165_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_166_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_166_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_166_rd_data          (fwd_tbl0_rdata[41][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_166_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_167_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_167_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_167_rd_data          (fwd_tbl0_rdata[41][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_167_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_168_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_168_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_168_rd_data          (fwd_tbl0_rdata[42][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_168_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_169_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_169_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_169_rd_data          (fwd_tbl0_rdata[42][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_169_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_16_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_16_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_16_rd_data           (fwd_tbl0_rdata[4][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_16_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_170_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_170_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_170_rd_data          (fwd_tbl0_rdata[42][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_170_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_171_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_171_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_171_rd_data          (fwd_tbl0_rdata[42][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_171_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_172_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_173_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_173_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_173_rd_data          (fwd_tbl0_rdata[43][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_173_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_174_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_174_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_174_rd_data          (fwd_tbl0_rdata[43][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_174_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_175_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_175_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_175_rd_data          (fwd_tbl0_rdata[43][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_175_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_176_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_176_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_176_rd_data          (fwd_tbl0_rdata[44][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_176_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_177_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_177_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_177_rd_data          (fwd_tbl0_rdata[44][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_177_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_178_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_178_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_178_rd_data          (fwd_tbl0_rdata[44][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_178_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_179_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_179_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_179_rd_data          (fwd_tbl0_rdata[44][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_179_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_17_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_17_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_17_rd_data           (fwd_tbl0_rdata[4][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_17_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_180_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_180_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_180_rd_data          (fwd_tbl0_rdata[45][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_180_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_181_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_181_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_181_rd_data          (fwd_tbl0_rdata[45][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_181_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_182_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_182_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_182_rd_data          (fwd_tbl0_rdata[45][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_182_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_183_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_183_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_183_rd_data          (fwd_tbl0_rdata[45][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_183_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_184_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_184_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_184_rd_data          (fwd_tbl0_rdata[46][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_184_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_185_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_185_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_185_rd_data          (fwd_tbl0_rdata[46][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_185_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_186_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_186_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_186_rd_data          (fwd_tbl0_rdata[46][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_186_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_187_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_187_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_187_rd_data          (fwd_tbl0_rdata[46][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_187_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_188_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_188_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_188_rd_data          (fwd_tbl0_rdata[47][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_188_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_189_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_189_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_189_rd_data          (fwd_tbl0_rdata[47][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_189_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_18_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_18_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_18_rd_data           (fwd_tbl0_rdata[4][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_18_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_190_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_190_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_190_rd_data          (fwd_tbl0_rdata[47][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_190_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_191_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_19_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_19_rd_data           (fwd_tbl0_rdata[4][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_19_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_1_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_1_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_1_rd_data            (fwd_tbl0_rdata[0][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_1_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_20_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_20_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_20_rd_data           (fwd_tbl0_rdata[5][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_20_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_21_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_21_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_21_rd_data           (fwd_tbl0_rdata[5][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_21_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_22_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_22_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_22_rd_data           (fwd_tbl0_rdata[5][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_22_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_23_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_23_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_23_rd_data           (fwd_tbl0_rdata[5][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_23_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_24_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_24_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_24_rd_data           (fwd_tbl0_rdata[6][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_24_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_25_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_25_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_25_rd_data           (fwd_tbl0_rdata[6][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_25_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_26_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_26_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_26_rd_data           (fwd_tbl0_rdata[6][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_26_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_27_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_27_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_27_rd_data           (fwd_tbl0_rdata[6][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_27_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_28_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_28_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_28_rd_data           (fwd_tbl0_rdata[7][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_28_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_29_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_29_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_29_rd_data           (fwd_tbl0_rdata[7][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_29_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_2_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_2_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_2_rd_data            (fwd_tbl0_rdata[0][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_2_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_30_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_30_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_30_rd_data           (fwd_tbl0_rdata[7][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_30_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_31_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_31_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_31_rd_data           (fwd_tbl0_rdata[7][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_31_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_32_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_32_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_32_rd_data           (fwd_tbl0_rdata[8][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_32_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_33_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_33_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_33_rd_data           (fwd_tbl0_rdata[8][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_33_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_34_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_34_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_34_rd_data           (fwd_tbl0_rdata[8][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_34_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_35_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_35_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_35_rd_data           (fwd_tbl0_rdata[8][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_35_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_36_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_36_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_36_rd_data           (fwd_tbl0_rdata[9][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_36_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_37_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_37_init_done         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_38_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_38_rd_data           (fwd_tbl0_rdata[9][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_38_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_39_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_39_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_39_rd_data           (fwd_tbl0_rdata[9][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_39_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_3_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_3_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_3_rd_data            (fwd_tbl0_rdata[0][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_3_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_40_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_40_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_40_rd_data           (fwd_tbl0_rdata[10][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_40_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_41_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_41_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_41_rd_data           (fwd_tbl0_rdata[10][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_41_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_42_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_42_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_42_rd_data           (fwd_tbl0_rdata[10][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_42_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_43_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_43_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_43_rd_data           (fwd_tbl0_rdata[10][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_43_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_44_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_44_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_44_rd_data           (fwd_tbl0_rdata[11][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_44_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_45_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_45_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_45_rd_data           (fwd_tbl0_rdata[11][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_45_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_46_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_46_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_46_rd_data           (fwd_tbl0_rdata[11][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_46_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_47_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_47_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_47_rd_data           (fwd_tbl0_rdata[11][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_47_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_48_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_48_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_48_rd_data           (fwd_tbl0_rdata[12][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_48_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_49_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_49_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_49_rd_data           (fwd_tbl0_rdata[12][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_49_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_4_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_4_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_4_rd_data            (fwd_tbl0_rdata[1][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_4_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_50_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_50_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_50_rd_data           (fwd_tbl0_rdata[12][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_50_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_51_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_51_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_51_rd_data           (fwd_tbl0_rdata[12][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_51_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_52_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_52_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_52_rd_data           (fwd_tbl0_rdata[13][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_52_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_53_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_53_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_53_rd_data           (fwd_tbl0_rdata[13][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_53_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_54_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_54_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_54_rd_data           (fwd_tbl0_rdata[13][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_54_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_55_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_55_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_55_rd_data           (fwd_tbl0_rdata[13][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_55_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_56_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_56_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_56_rd_data           (fwd_tbl0_rdata[14][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_56_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_57_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_57_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_58_rd_data           (fwd_tbl0_rdata[14][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_58_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_59_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_59_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_59_rd_data           (fwd_tbl0_rdata[14][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_59_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_5_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_5_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_5_rd_data            (fwd_tbl0_rdata[1][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_5_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_60_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_60_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_60_rd_data           (fwd_tbl0_rdata[15][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_60_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_61_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_61_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_61_rd_data           (fwd_tbl0_rdata[15][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_61_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_62_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_62_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_62_rd_data           (fwd_tbl0_rdata[15][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_62_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_63_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_63_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_63_rd_data           (fwd_tbl0_rdata[15][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_63_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_64_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_64_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_64_rd_data           (fwd_tbl0_rdata[16][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_64_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_65_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_65_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_65_rd_data           (fwd_tbl0_rdata[16][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_65_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_66_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_66_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_66_rd_data           (fwd_tbl0_rdata[16][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_66_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_67_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_67_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_67_rd_data           (fwd_tbl0_rdata[16][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_67_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_68_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_68_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_68_rd_data           (fwd_tbl0_rdata[17][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_68_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_69_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_69_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_69_rd_data           (fwd_tbl0_rdata[17][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_69_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_6_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_6_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_6_rd_data            (fwd_tbl0_rdata[1][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_6_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_70_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_70_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_70_rd_data           (fwd_tbl0_rdata[17][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_70_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_71_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_71_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_71_rd_data           (fwd_tbl0_rdata[17][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_71_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_72_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_72_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_72_rd_data           (fwd_tbl0_rdata[18][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_72_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_73_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_73_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_73_rd_data           (fwd_tbl0_rdata[18][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_73_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_74_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_74_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_74_rd_data           (fwd_tbl0_rdata[18][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_74_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_75_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_75_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_75_rd_data           (fwd_tbl0_rdata[18][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_75_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_76_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_76_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_77_rd_data           (fwd_tbl0_rdata[19][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_77_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_78_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_78_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_78_rd_data           (fwd_tbl0_rdata[19][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_78_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_79_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_79_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_79_rd_data           (fwd_tbl0_rdata[19][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_79_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_7_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_7_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_7_rd_data            (fwd_tbl0_rdata[1][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_7_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_80_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_80_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_80_rd_data           (fwd_tbl0_rdata[20][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_80_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_81_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_81_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_81_rd_data           (fwd_tbl0_rdata[20][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_81_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_82_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_82_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_82_rd_data           (fwd_tbl0_rdata[20][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_82_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_83_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_83_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_83_rd_data           (fwd_tbl0_rdata[20][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_83_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_84_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_84_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_84_rd_data           (fwd_tbl0_rdata[21][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_84_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_85_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_85_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_85_rd_data           (fwd_tbl0_rdata[21][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_85_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_86_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_86_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_86_rd_data           (fwd_tbl0_rdata[21][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_86_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_87_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_87_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_87_rd_data           (fwd_tbl0_rdata[21][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_87_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_88_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_88_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_88_rd_data           (fwd_tbl0_rdata[22][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_88_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_89_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_89_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_89_rd_data           (fwd_tbl0_rdata[22][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_89_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_8_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_8_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_8_rd_data            (fwd_tbl0_rdata[2][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_8_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_90_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_90_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_90_rd_data           (fwd_tbl0_rdata[22][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_90_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_91_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_91_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_91_rd_data           (fwd_tbl0_rdata[22][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_91_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_92_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_92_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_92_rd_data           (fwd_tbl0_rdata[23][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_92_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_93_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_93_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_93_rd_data           (fwd_tbl0_rdata[23][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_93_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_94_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_94_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_94_rd_data           (fwd_tbl0_rdata[23][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_94_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_95_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_95_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_95_rd_data           (fwd_tbl0_rdata[23][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_95_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_96_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_96_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_96_rd_data           (fwd_tbl0_rdata[24][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_97_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_98_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_98_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_98_rd_data           (fwd_tbl0_rdata[24][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_98_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_99_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_99_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_99_rd_data           (fwd_tbl0_rdata[24][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_99_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_9_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_9_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_9_rd_data            (fwd_tbl0_rdata[2][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_9_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_0_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_0_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_0_rd_data            (fwd_tbl1_rdata[0][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_0_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_10_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_10_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_10_rd_data           (fwd_tbl1_rdata[2][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_10_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_11_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_11_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_11_rd_data           (fwd_tbl1_rdata[2][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_11_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_12_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_12_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_12_rd_data           (fwd_tbl1_rdata[3][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_12_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_13_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_13_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_13_rd_data           (fwd_tbl1_rdata[3][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_13_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_14_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_14_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_14_rd_data           (fwd_tbl1_rdata[3][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_14_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_15_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_15_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_15_rd_data           (fwd_tbl1_rdata[3][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_15_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_16_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_16_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_16_rd_data           (fwd_tbl1_rdata[4][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_16_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_17_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_17_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_17_rd_data           (fwd_tbl1_rdata[4][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_17_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_18_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_18_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_18_rd_data           (fwd_tbl1_rdata[4][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_18_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_19_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_19_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_19_rd_data           (fwd_tbl1_rdata[4][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_19_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_1_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_1_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_1_rd_data            (fwd_tbl1_rdata[0][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_1_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_20_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_20_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_20_rd_data           (fwd_tbl1_rdata[5][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_20_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_21_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_21_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_21_rd_data           (fwd_tbl1_rdata[5][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_21_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_22_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_22_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_22_rd_data           (fwd_tbl1_rdata[5][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_22_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_23_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_23_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_23_rd_data           (fwd_tbl1_rdata[5][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_23_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_24_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_24_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_24_rd_data           (fwd_tbl1_rdata[6][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_25_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_26_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_26_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_26_rd_data           (fwd_tbl1_rdata[6][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_26_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_27_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_27_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_27_rd_data           (fwd_tbl1_rdata[6][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_27_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_28_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_28_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_28_rd_data           (fwd_tbl1_rdata[7][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_28_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_29_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_29_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_29_rd_data           (fwd_tbl1_rdata[7][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_29_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_2_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_2_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_2_rd_data            (fwd_tbl1_rdata[0][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_2_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_30_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_30_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_30_rd_data           (fwd_tbl1_rdata[7][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_30_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_31_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_31_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_31_rd_data           (fwd_tbl1_rdata[7][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_31_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_32_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_32_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_32_rd_data           (fwd_tbl1_rdata[8][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_32_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_33_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_33_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_33_rd_data           (fwd_tbl1_rdata[8][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_33_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_34_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_34_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_34_rd_data           (fwd_tbl1_rdata[8][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_34_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_35_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_35_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_35_rd_data           (fwd_tbl1_rdata[8][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_35_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_36_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_36_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_36_rd_data           (fwd_tbl1_rdata[9][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_36_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_37_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_37_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_37_rd_data           (fwd_tbl1_rdata[9][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_37_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_38_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_38_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_38_rd_data           (fwd_tbl1_rdata[9][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_38_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_39_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_39_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_39_rd_data           (fwd_tbl1_rdata[9][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_39_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_3_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_3_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_3_rd_data            (fwd_tbl1_rdata[0][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_3_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_40_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_40_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_40_rd_data           (fwd_tbl1_rdata[10][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_40_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_41_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_41_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_41_rd_data           (fwd_tbl1_rdata[10][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_41_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_42_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_42_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_42_rd_data           (fwd_tbl1_rdata[10][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_42_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_43_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_43_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_43_rd_data           (fwd_tbl1_rdata[10][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_43_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_44_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_44_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_44_rd_data           (fwd_tbl1_rdata[11][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_44_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_46_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_46_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_46_rd_data           (fwd_tbl1_rdata[11][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_46_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_47_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_47_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_47_rd_data           (fwd_tbl1_rdata[11][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_47_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_48_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_48_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_48_rd_data           (fwd_tbl1_rdata[12][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_48_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_49_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_49_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_49_rd_data           (fwd_tbl1_rdata[12][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_49_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_4_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_4_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_4_rd_data            (fwd_tbl1_rdata[1][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_4_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_50_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_50_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_50_rd_data           (fwd_tbl1_rdata[12][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_50_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_51_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_51_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_51_rd_data           (fwd_tbl1_rdata[12][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_51_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_52_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_52_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_52_rd_data           (fwd_tbl1_rdata[13][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_52_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_53_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_53_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_53_rd_data           (fwd_tbl1_rdata[13][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_53_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_54_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_54_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_54_rd_data           (fwd_tbl1_rdata[13][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_54_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_55_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_55_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_55_rd_data           (fwd_tbl1_rdata[13][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_55_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_56_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_56_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_56_rd_data           (fwd_tbl1_rdata[14][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_56_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_57_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_57_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_57_rd_data           (fwd_tbl1_rdata[14][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_57_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_58_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_58_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_58_rd_data           (fwd_tbl1_rdata[14][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_58_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_59_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_59_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_59_rd_data           (fwd_tbl1_rdata[14][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_59_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_5_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_5_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_5_rd_data            (fwd_tbl1_rdata[1][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_5_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_60_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_60_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_60_rd_data           (fwd_tbl1_rdata[15][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_60_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_61_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_61_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_61_rd_data           (fwd_tbl1_rdata[15][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_61_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_62_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_62_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_62_rd_data           (fwd_tbl1_rdata[15][2][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_62_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_63_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_63_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_63_rd_data           (fwd_tbl1_rdata[15][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_63_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_7_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_7_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_7_rd_data            (fwd_tbl1_rdata[1][3][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_7_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_8_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_8_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_8_rd_data            (fwd_tbl1_rdata[2][0][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_8_rd_valid           (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_9_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_9_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_9_rd_data            (fwd_tbl1_rdata[2][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_9_rd_valid           (),                                                
/* output logic          */ .ppe_stm_init_done                     (),                                                
/* output logic          */ .ppe_stm_l3mc_tbl_ecc_uncor_err        (),                                                
/* output logic          */ .ppe_stm_l3mc_tbl_init_done            (),                                                
/* output logic  [511:0] */ .ppe_stm_l3mc_tbl_rd_data              (),                                                
/* output logic          */ .ppe_stm_l3mc_tbl_rd_valid             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_0_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_0_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_0_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_0_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_10_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_10_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_10_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_10_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_11_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_11_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_11_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_11_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_12_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_12_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_12_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_12_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_13_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_13_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_13_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_13_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_14_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_14_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_14_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_14_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_15_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_15_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_15_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_15_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_16_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_16_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_16_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_16_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_17_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_17_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_17_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_17_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_18_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_18_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_18_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_18_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_19_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_19_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_19_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_19_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_1_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_1_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_1_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_1_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_20_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_20_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_20_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_20_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_21_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_21_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_21_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_21_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_22_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_22_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_22_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_22_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_23_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_23_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_23_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_23_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_24_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_24_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_24_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_24_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_25_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_26_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_26_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_26_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_26_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_27_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_27_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_27_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_27_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_28_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_28_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_28_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_28_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_29_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_29_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_29_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_29_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_2_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_2_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_2_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_2_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_30_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_30_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_30_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_30_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_31_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_31_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_31_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_31_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_32_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_32_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_32_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_32_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_33_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_33_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_33_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_33_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_34_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_34_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_34_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_34_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_35_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_35_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_35_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_35_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_36_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_36_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_36_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_36_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_37_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_37_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_37_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_37_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_38_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_38_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_38_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_38_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_39_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_39_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_39_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_39_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_3_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_3_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_3_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_3_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_40_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_40_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_40_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_40_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_41_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_41_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_41_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_41_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_42_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_42_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_42_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_42_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_43_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_43_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_43_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_43_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_45_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_45_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_45_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_45_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_46_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_46_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_46_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_46_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_47_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_47_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_47_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_47_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_48_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_48_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_48_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_48_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_49_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_49_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_49_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_49_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_4_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_4_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_4_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_4_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_50_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_50_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_50_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_50_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_51_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_51_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_51_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_51_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_52_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_52_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_52_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_52_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_53_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_53_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_53_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_53_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_54_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_54_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_54_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_54_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_55_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_55_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_55_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_55_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_56_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_56_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_56_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_56_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_57_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_57_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_57_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_57_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_58_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_58_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_58_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_58_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_59_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_59_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_59_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_59_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_5_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_5_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_5_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_5_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_60_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_60_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_60_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_60_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_61_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_61_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_61_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_61_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_62_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_62_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_62_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_62_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_63_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_63_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_63_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_63_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_64_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_64_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_64_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_64_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_65_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_65_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_65_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_65_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_66_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_66_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_66_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_66_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_67_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_67_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_67_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_67_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_68_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_68_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_68_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_68_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_69_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_69_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_69_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_69_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_6_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_6_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_6_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_6_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_70_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_70_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_70_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_70_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_71_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_71_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_71_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_71_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_72_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_72_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_72_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_72_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_73_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_73_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_73_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_73_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_74_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_74_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_74_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_74_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_75_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_75_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_75_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_75_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_76_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_76_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_76_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_76_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_77_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_77_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_77_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_77_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_78_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_78_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_78_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_78_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_79_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_79_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_79_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_79_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_7_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_7_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_7_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_7_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_8_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_8_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_8_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_8_rd_valid            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_9_ecc_uncor_err       (),                                                
/* output logic          */ .ppe_stm_mod_tbl_9_init_done           (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_9_rd_data             (),                                                
/* output logic          */ .ppe_stm_mod_tbl_9_rd_valid            (),                                                
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_0_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_0_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_100_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_100_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_101_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_101_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_102_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_102_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_103_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_103_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_108_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_108_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_109_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_109_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_10_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_10_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_110_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_110_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_111_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_111_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_112_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_112_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_113_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_113_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_114_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_114_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_115_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_115_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_116_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_116_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_117_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_117_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_118_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_118_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_119_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_119_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_11_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_11_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_120_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_120_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_121_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_121_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_122_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_122_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_123_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_123_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_124_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_124_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_125_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_125_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_126_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_126_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_127_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_127_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_128_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_128_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_129_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_129_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_12_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_12_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_130_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_130_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_131_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_131_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_163_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_163_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_164_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_164_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_165_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_165_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_166_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_166_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_167_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_167_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_168_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_168_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_169_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_169_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_16_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_16_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_170_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_170_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_171_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_171_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_172_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_172_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_173_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_173_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_174_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_174_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_175_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_175_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_176_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_176_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_177_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_177_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_178_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_178_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_179_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_179_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_17_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_17_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_180_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_180_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_181_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_181_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_182_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_182_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_183_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_183_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_184_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_184_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_185_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_185_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_186_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_186_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_187_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_187_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_188_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_188_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_189_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_189_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_18_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_18_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_190_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_190_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_191_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_191_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_19_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_19_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_1_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_1_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_20_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_20_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_21_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_21_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_22_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_22_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_23_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_23_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_24_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_24_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_25_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_25_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_26_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_26_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_27_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_27_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_28_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_28_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_29_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_29_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_2_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_2_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_30_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_30_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_31_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_31_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_32_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_32_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_33_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_33_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_34_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_34_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_35_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_35_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_36_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_36_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_37_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_37_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_38_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_38_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_39_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_39_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_3_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_3_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_40_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_40_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_41_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_41_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_46_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_46_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_47_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_47_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_48_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_48_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_49_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_49_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_4_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_4_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_50_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_50_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_51_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_51_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_52_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_52_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_53_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_53_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_54_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_54_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_55_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_55_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_56_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_56_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_57_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_57_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_58_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_58_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_59_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_59_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_5_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_5_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_60_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_60_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_61_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_61_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_62_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_62_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_63_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_63_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_64_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_64_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_65_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_65_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_66_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_66_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_67_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_67_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_68_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_68_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_69_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_69_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_6_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_6_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_70_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_70_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_71_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_71_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_72_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_72_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_73_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_73_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_74_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_74_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_75_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_75_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_76_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_76_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_77_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_77_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_78_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_78_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_79_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_79_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_7_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_7_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_80_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_80_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_81_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_81_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_82_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_82_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_83_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_83_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_84_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_84_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_85_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_85_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_86_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_86_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_87_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_87_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_88_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_88_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_89_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_89_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_8_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_8_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_90_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_90_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_91_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_91_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_92_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_92_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_93_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_93_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_94_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_94_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_95_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_95_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_96_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_96_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_97_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_97_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_98_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_98_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_99_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_99_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_9_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_9_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_0_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_0_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_10_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_10_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_11_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_11_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_12_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_12_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_13_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_13_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_14_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_14_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_15_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_15_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_16_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_16_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_17_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_17_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_18_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_18_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_19_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_19_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_1_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_1_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_20_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_20_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_21_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_21_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_22_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_22_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_23_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_23_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_24_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_24_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_25_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_25_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_26_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_26_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_27_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_27_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_28_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_28_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_29_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_29_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_2_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_2_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_30_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_30_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_31_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_31_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_32_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_32_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_33_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_33_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_34_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_34_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_35_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_35_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_36_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_36_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_37_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_37_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_38_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_38_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_39_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_39_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_3_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_3_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_40_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_40_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_41_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_41_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_42_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_42_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_43_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_43_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_44_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_44_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_45_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_45_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_46_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_46_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_47_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_47_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_48_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_48_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_49_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_49_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_4_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_4_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_50_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_50_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_51_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_51_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_52_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_52_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_53_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_53_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_54_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_54_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_55_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_55_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_56_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_56_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_57_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_57_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_58_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_58_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_59_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_59_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_5_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_5_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_60_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_60_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_61_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_61_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_62_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_62_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_9_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_9_to_mem),               
/* output logic  [596:0] */ .ppe_stm_ppe_stm_l3mc_tbl_to_mem       (ppe_stm_ppe_stm_l3mc_tbl_to_mem),                 
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_0_to_mem      (ppe_stm_ppe_stm_mod_tbl_0_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_10_to_mem     (ppe_stm_ppe_stm_mod_tbl_10_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_11_to_mem     (ppe_stm_ppe_stm_mod_tbl_11_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_12_to_mem     (ppe_stm_ppe_stm_mod_tbl_12_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_13_to_mem     (ppe_stm_ppe_stm_mod_tbl_13_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_14_to_mem     (ppe_stm_ppe_stm_mod_tbl_14_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_15_to_mem     (ppe_stm_ppe_stm_mod_tbl_15_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_16_to_mem     (ppe_stm_ppe_stm_mod_tbl_16_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_17_to_mem     (ppe_stm_ppe_stm_mod_tbl_17_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_18_to_mem     (ppe_stm_ppe_stm_mod_tbl_18_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_19_to_mem     (ppe_stm_ppe_stm_mod_tbl_19_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_1_to_mem      (ppe_stm_ppe_stm_mod_tbl_1_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_20_to_mem     (ppe_stm_ppe_stm_mod_tbl_20_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_21_to_mem     (ppe_stm_ppe_stm_mod_tbl_21_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_22_to_mem     (ppe_stm_ppe_stm_mod_tbl_22_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_23_to_mem     (ppe_stm_ppe_stm_mod_tbl_23_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_24_to_mem     (ppe_stm_ppe_stm_mod_tbl_24_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_25_to_mem     (ppe_stm_ppe_stm_mod_tbl_25_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_26_to_mem     (ppe_stm_ppe_stm_mod_tbl_26_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_27_to_mem     (ppe_stm_ppe_stm_mod_tbl_27_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_28_to_mem     (ppe_stm_ppe_stm_mod_tbl_28_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_29_to_mem     (ppe_stm_ppe_stm_mod_tbl_29_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_2_to_mem      (ppe_stm_ppe_stm_mod_tbl_2_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_30_to_mem     (ppe_stm_ppe_stm_mod_tbl_30_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_31_to_mem     (ppe_stm_ppe_stm_mod_tbl_31_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_32_to_mem     (ppe_stm_ppe_stm_mod_tbl_32_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_33_to_mem     (ppe_stm_ppe_stm_mod_tbl_33_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_34_to_mem     (ppe_stm_ppe_stm_mod_tbl_34_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_35_to_mem     (ppe_stm_ppe_stm_mod_tbl_35_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_36_to_mem     (ppe_stm_ppe_stm_mod_tbl_36_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_37_to_mem     (ppe_stm_ppe_stm_mod_tbl_37_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_38_to_mem     (ppe_stm_ppe_stm_mod_tbl_38_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_39_to_mem     (ppe_stm_ppe_stm_mod_tbl_39_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_3_to_mem      (ppe_stm_ppe_stm_mod_tbl_3_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_40_to_mem     (ppe_stm_ppe_stm_mod_tbl_40_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_41_to_mem     (ppe_stm_ppe_stm_mod_tbl_41_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_42_to_mem     (ppe_stm_ppe_stm_mod_tbl_42_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_43_to_mem     (ppe_stm_ppe_stm_mod_tbl_43_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_44_to_mem     (ppe_stm_ppe_stm_mod_tbl_44_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_45_to_mem     (ppe_stm_ppe_stm_mod_tbl_45_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_46_to_mem     (ppe_stm_ppe_stm_mod_tbl_46_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_47_to_mem     (ppe_stm_ppe_stm_mod_tbl_47_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_48_to_mem     (ppe_stm_ppe_stm_mod_tbl_48_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_49_to_mem     (ppe_stm_ppe_stm_mod_tbl_49_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_4_to_mem      (ppe_stm_ppe_stm_mod_tbl_4_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_50_to_mem     (ppe_stm_ppe_stm_mod_tbl_50_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_51_to_mem     (ppe_stm_ppe_stm_mod_tbl_51_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_52_to_mem     (ppe_stm_ppe_stm_mod_tbl_52_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_53_to_mem     (ppe_stm_ppe_stm_mod_tbl_53_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_54_to_mem     (ppe_stm_ppe_stm_mod_tbl_54_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_55_to_mem     (ppe_stm_ppe_stm_mod_tbl_55_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_56_to_mem     (ppe_stm_ppe_stm_mod_tbl_56_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_57_to_mem     (ppe_stm_ppe_stm_mod_tbl_57_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_58_to_mem     (ppe_stm_ppe_stm_mod_tbl_58_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_59_to_mem     (ppe_stm_ppe_stm_mod_tbl_59_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_5_to_mem      (ppe_stm_ppe_stm_mod_tbl_5_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_60_to_mem     (ppe_stm_ppe_stm_mod_tbl_60_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_61_to_mem     (ppe_stm_ppe_stm_mod_tbl_61_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_62_to_mem     (ppe_stm_ppe_stm_mod_tbl_62_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_63_to_mem     (ppe_stm_ppe_stm_mod_tbl_63_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_64_to_mem     (ppe_stm_ppe_stm_mod_tbl_64_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_65_to_mem     (ppe_stm_ppe_stm_mod_tbl_65_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_66_to_mem     (ppe_stm_ppe_stm_mod_tbl_66_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_67_to_mem     (ppe_stm_ppe_stm_mod_tbl_67_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_68_to_mem     (ppe_stm_ppe_stm_mod_tbl_68_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_69_to_mem     (ppe_stm_ppe_stm_mod_tbl_69_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_6_to_mem      (ppe_stm_ppe_stm_mod_tbl_6_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_70_to_mem     (ppe_stm_ppe_stm_mod_tbl_70_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_71_to_mem     (ppe_stm_ppe_stm_mod_tbl_71_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_72_to_mem     (ppe_stm_ppe_stm_mod_tbl_72_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_73_to_mem     (ppe_stm_ppe_stm_mod_tbl_73_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_74_to_mem     (ppe_stm_ppe_stm_mod_tbl_74_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_75_to_mem     (ppe_stm_ppe_stm_mod_tbl_75_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_76_to_mem     (ppe_stm_ppe_stm_mod_tbl_76_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_77_to_mem     (ppe_stm_ppe_stm_mod_tbl_77_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_78_to_mem     (ppe_stm_ppe_stm_mod_tbl_78_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_79_to_mem     (ppe_stm_ppe_stm_mod_tbl_79_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_7_to_mem      (ppe_stm_ppe_stm_mod_tbl_7_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_8_to_mem      (ppe_stm_ppe_stm_mod_tbl_8_to_mem),                
/* output logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_9_to_mem      (ppe_stm_ppe_stm_mod_tbl_9_to_mem),                
/* output logic   [63:0] */ .ppe_stm_ppe_stm_shcp_tbl_to_mem       (ppe_stm_ppe_stm_shcp_tbl_to_mem),                 
/* output logic          */ .ppe_stm_shcp_tbl_ecc_uncor_err        (),                                                
/* output logic          */ .ppe_stm_shcp_tbl_init_done            (),                                                
/* output logic   [32:0] */ .ppe_stm_shcp_tbl_rd_data              (),                                                
/* output logic          */ .ppe_stm_shcp_tbl_rd_valid             (),                                                
/* output logic          */ .unified_regs_ack                      (),                                                
/* output logic   [31:0] */ .unified_regs_rd_data                  (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_133_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_133_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_133_rd_data          (fwd_tbl0_rdata[33][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_133_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_152_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_152_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_152_rd_data          (fwd_tbl0_rdata[38][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_152_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_24_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_25_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_25_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_25_rd_data           (fwd_tbl1_rdata[6][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_45_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_45_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_45_rd_data           (fwd_tbl1_rdata[11][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl1_45_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_112_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_113_ecc_uncor_err    (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_113_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_113_rd_data          (fwd_tbl0_rdata[28][1][71:0]),                     
/* output logic          */ .ppe_stm_mod_tbl_44_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_44_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_44_rd_data            (),                                                
/* output logic          */ .ppe_stm_mod_tbl_44_rd_valid           (),                                                
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_42_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_42_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_43_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_43_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_44_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_44_to_mem),              
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_45_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_45_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_63_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_63_to_mem),              
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_6_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_6_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_7_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_7_to_mem),               
/* output logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_8_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_8_to_mem),               
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_104_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_104_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_105_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_105_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_106_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_106_to_mem),             
/* output logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_107_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_107_to_mem),             
/* output logic          */ .ppe_stm_fwd_tbl0_172_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_172_rd_data          (fwd_tbl0_rdata[43][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_172_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_191_init_done        (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_191_rd_data          (fwd_tbl0_rdata[47][3][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_191_rd_valid         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_19_ecc_uncor_err     (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_37_rd_data           (fwd_tbl0_rdata[9][1][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl0_37_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_38_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_6_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_fwd_tbl1_6_init_done          (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl1_6_rd_data            (fwd_tbl1_rdata[1][2][71:0]),                      
/* output logic          */ .ppe_stm_fwd_tbl1_6_rd_valid           (),                                                
/* output logic          */ .ppe_stm_mod_tbl_25_ecc_uncor_err      (),                                                
/* output logic          */ .ppe_stm_mod_tbl_25_init_done          (),                                                
/* output logic   [63:0] */ .ppe_stm_mod_tbl_25_rd_data            (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_76_rd_data           (fwd_tbl0_rdata[19][0][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_76_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_77_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_77_init_done         (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_96_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_97_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_97_init_done         (),                                                
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_97_rd_data           (fwd_tbl0_rdata[24][1][71:0]),                     
/* output logic   [71:0] */ .ppe_stm_fwd_tbl0_57_rd_data           (fwd_tbl0_rdata[14][1][71:0]),                     
/* output logic          */ .ppe_stm_fwd_tbl0_57_rd_valid          (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_58_ecc_uncor_err     (),                                                
/* output logic          */ .ppe_stm_fwd_tbl0_58_init_done         ());                                                
// End of module ppe_stm_shells_wrapper from ppe_stm_shells_wrapper


// module ppe_stm_sram_mems    from ppe_stm_sram_mems using ppe_stm_sram_mems.map 
ppe_stm_sram_mems    ppe_stm_sram_mems(
/* input  logic          */ .fscan_ram_init_en                     (),                                                
/* input  logic          */ .fscan_ram_init_val                    (),                                                
/* input  logic  [337:0] */ .fscan_ram_odis_b                      (),                                                
/* input  logic          */ .fscan_ram_rddis_b                     (),                                                
/* input  logic          */ .fscan_ram_wrdis_b                     (),                                                
/* input  logic          */ .fscan_rstbypen                        (),                                                
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_0_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_0_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_100_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_100_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_101_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_101_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_102_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_102_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_103_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_103_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_104_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_104_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_105_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_105_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_106_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_106_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_107_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_107_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_108_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_108_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_109_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_109_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_10_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_10_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_110_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_110_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_111_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_111_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_112_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_112_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_113_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_113_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_114_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_114_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_115_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_115_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_116_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_116_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_117_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_117_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_118_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_118_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_119_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_119_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_11_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_11_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_120_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_120_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_121_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_121_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_122_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_122_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_123_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_123_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_124_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_124_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_125_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_125_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_126_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_126_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_127_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_127_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_128_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_128_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_129_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_129_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_12_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_12_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_130_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_130_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_131_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_131_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_132_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_132_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_133_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_133_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_134_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_134_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_135_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_135_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_136_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_136_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_137_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_137_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_138_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_138_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_139_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_139_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_13_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_13_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_140_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_140_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_141_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_141_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_142_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_142_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_143_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_143_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_144_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_144_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_145_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_145_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_146_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_146_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_147_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_147_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_148_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_148_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_149_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_149_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_14_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_14_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_150_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_150_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_151_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_151_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_152_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_152_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_153_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_153_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_154_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_154_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_155_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_155_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_156_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_156_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_157_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_157_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_158_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_158_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_159_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_159_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_15_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_15_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_160_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_160_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_161_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_161_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_162_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_162_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_163_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_163_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_168_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_168_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_169_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_169_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_16_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_16_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_170_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_170_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_171_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_171_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_172_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_172_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_173_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_173_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_174_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_174_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_175_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_175_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_176_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_176_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_177_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_177_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_178_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_178_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_179_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_179_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_17_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_17_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_180_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_180_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_181_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_181_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_182_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_182_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_183_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_183_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_184_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_184_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_185_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_185_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_186_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_186_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_187_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_187_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_188_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_188_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_189_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_189_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_18_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_18_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_190_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_190_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_191_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_191_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_19_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_19_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_1_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_1_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_20_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_20_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_21_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_21_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_22_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_22_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_23_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_23_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_24_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_24_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_25_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_25_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_26_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_26_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_27_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_27_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_28_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_28_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_29_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_29_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_2_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_2_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_30_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_30_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_31_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_31_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_32_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_32_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_33_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_33_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_34_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_34_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_35_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_35_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_36_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_36_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_37_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_37_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_38_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_38_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_39_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_39_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_3_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_3_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_40_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_40_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_41_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_41_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_42_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_42_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_43_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_43_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_44_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_44_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_45_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_45_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_46_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_46_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_47_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_47_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_48_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_48_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_49_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_49_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_4_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_4_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_50_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_50_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_51_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_51_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_52_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_52_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_53_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_53_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_54_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_54_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_55_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_55_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_56_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_56_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_57_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_57_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_58_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_58_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_59_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_59_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_5_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_5_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_60_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_60_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_61_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_61_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_62_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_62_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_63_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_63_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_64_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_64_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_65_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_65_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_66_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_66_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_67_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_67_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_68_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_68_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_69_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_69_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_6_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_6_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_70_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_70_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_71_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_71_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_72_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_72_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_73_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_73_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_74_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_74_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_75_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_75_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_76_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_76_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_77_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_77_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_78_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_78_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_79_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_79_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_7_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_7_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_80_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_80_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_81_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_81_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_82_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_82_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_83_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_83_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_84_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_84_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_85_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_85_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_86_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_86_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_87_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_87_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_88_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_88_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_89_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_89_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_8_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_8_to_mem),               
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_90_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_90_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_91_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_91_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_92_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_92_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_93_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_93_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_94_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_94_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_95_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_95_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_96_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_96_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_97_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_97_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_98_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_98_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_99_to_mem    (ppe_stm_ppe_stm_fwd_tbl0_99_to_mem),              
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_9_to_mem     (ppe_stm_ppe_stm_fwd_tbl0_9_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_0_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_0_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_10_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_10_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_15_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_15_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_16_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_16_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_17_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_17_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_18_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_18_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_19_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_19_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_1_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_1_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_20_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_20_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_21_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_21_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_22_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_22_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_23_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_23_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_24_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_24_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_25_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_25_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_26_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_26_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_27_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_27_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_28_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_28_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_29_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_29_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_2_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_2_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_30_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_30_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_31_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_31_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_32_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_32_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_33_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_33_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_34_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_34_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_35_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_35_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_36_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_36_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_37_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_37_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_38_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_38_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_39_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_39_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_3_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_3_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_40_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_40_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_41_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_41_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_42_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_42_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_43_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_43_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_44_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_44_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_45_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_45_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_46_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_46_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_47_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_47_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_48_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_48_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_49_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_49_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_4_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_4_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_50_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_50_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_51_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_51_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_52_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_52_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_53_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_53_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_54_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_54_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_55_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_55_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_56_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_56_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_57_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_57_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_58_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_58_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_59_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_59_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_5_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_5_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_60_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_60_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_61_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_61_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_62_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_62_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_63_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_63_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_6_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_6_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_7_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_7_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_8_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_8_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_9_to_mem     (ppe_stm_ppe_stm_fwd_tbl1_9_to_mem),               
/* input  logic  [596:0] */ .ppe_stm_ppe_stm_l3mc_tbl_to_mem       (ppe_stm_ppe_stm_l3mc_tbl_to_mem),                 
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_0_to_mem      (ppe_stm_ppe_stm_mod_tbl_0_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_10_to_mem     (ppe_stm_ppe_stm_mod_tbl_10_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_11_to_mem     (ppe_stm_ppe_stm_mod_tbl_11_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_12_to_mem     (ppe_stm_ppe_stm_mod_tbl_12_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_13_to_mem     (ppe_stm_ppe_stm_mod_tbl_13_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_14_to_mem     (ppe_stm_ppe_stm_mod_tbl_14_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_15_to_mem     (ppe_stm_ppe_stm_mod_tbl_15_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_16_to_mem     (ppe_stm_ppe_stm_mod_tbl_16_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_17_to_mem     (ppe_stm_ppe_stm_mod_tbl_17_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_18_to_mem     (ppe_stm_ppe_stm_mod_tbl_18_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_19_to_mem     (ppe_stm_ppe_stm_mod_tbl_19_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_1_to_mem      (ppe_stm_ppe_stm_mod_tbl_1_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_20_to_mem     (ppe_stm_ppe_stm_mod_tbl_20_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_21_to_mem     (ppe_stm_ppe_stm_mod_tbl_21_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_22_to_mem     (ppe_stm_ppe_stm_mod_tbl_22_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_23_to_mem     (ppe_stm_ppe_stm_mod_tbl_23_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_24_to_mem     (ppe_stm_ppe_stm_mod_tbl_24_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_25_to_mem     (ppe_stm_ppe_stm_mod_tbl_25_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_26_to_mem     (ppe_stm_ppe_stm_mod_tbl_26_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_27_to_mem     (ppe_stm_ppe_stm_mod_tbl_27_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_28_to_mem     (ppe_stm_ppe_stm_mod_tbl_28_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_29_to_mem     (ppe_stm_ppe_stm_mod_tbl_29_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_2_to_mem      (ppe_stm_ppe_stm_mod_tbl_2_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_30_to_mem     (ppe_stm_ppe_stm_mod_tbl_30_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_31_to_mem     (ppe_stm_ppe_stm_mod_tbl_31_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_32_to_mem     (ppe_stm_ppe_stm_mod_tbl_32_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_33_to_mem     (ppe_stm_ppe_stm_mod_tbl_33_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_34_to_mem     (ppe_stm_ppe_stm_mod_tbl_34_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_35_to_mem     (ppe_stm_ppe_stm_mod_tbl_35_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_36_to_mem     (ppe_stm_ppe_stm_mod_tbl_36_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_37_to_mem     (ppe_stm_ppe_stm_mod_tbl_37_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_38_to_mem     (ppe_stm_ppe_stm_mod_tbl_38_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_39_to_mem     (ppe_stm_ppe_stm_mod_tbl_39_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_3_to_mem      (ppe_stm_ppe_stm_mod_tbl_3_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_40_to_mem     (ppe_stm_ppe_stm_mod_tbl_40_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_41_to_mem     (ppe_stm_ppe_stm_mod_tbl_41_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_42_to_mem     (ppe_stm_ppe_stm_mod_tbl_42_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_43_to_mem     (ppe_stm_ppe_stm_mod_tbl_43_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_44_to_mem     (ppe_stm_ppe_stm_mod_tbl_44_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_45_to_mem     (ppe_stm_ppe_stm_mod_tbl_45_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_46_to_mem     (ppe_stm_ppe_stm_mod_tbl_46_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_47_to_mem     (ppe_stm_ppe_stm_mod_tbl_47_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_48_to_mem     (ppe_stm_ppe_stm_mod_tbl_48_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_49_to_mem     (ppe_stm_ppe_stm_mod_tbl_49_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_4_to_mem      (ppe_stm_ppe_stm_mod_tbl_4_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_50_to_mem     (ppe_stm_ppe_stm_mod_tbl_50_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_51_to_mem     (ppe_stm_ppe_stm_mod_tbl_51_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_52_to_mem     (ppe_stm_ppe_stm_mod_tbl_52_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_53_to_mem     (ppe_stm_ppe_stm_mod_tbl_53_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_54_to_mem     (ppe_stm_ppe_stm_mod_tbl_54_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_55_to_mem     (ppe_stm_ppe_stm_mod_tbl_55_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_56_to_mem     (ppe_stm_ppe_stm_mod_tbl_56_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_57_to_mem     (ppe_stm_ppe_stm_mod_tbl_57_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_58_to_mem     (ppe_stm_ppe_stm_mod_tbl_58_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_59_to_mem     (ppe_stm_ppe_stm_mod_tbl_59_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_5_to_mem      (ppe_stm_ppe_stm_mod_tbl_5_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_60_to_mem     (ppe_stm_ppe_stm_mod_tbl_60_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_61_to_mem     (ppe_stm_ppe_stm_mod_tbl_61_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_62_to_mem     (ppe_stm_ppe_stm_mod_tbl_62_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_63_to_mem     (ppe_stm_ppe_stm_mod_tbl_63_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_67_to_mem     (ppe_stm_ppe_stm_mod_tbl_67_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_68_to_mem     (ppe_stm_ppe_stm_mod_tbl_68_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_69_to_mem     (ppe_stm_ppe_stm_mod_tbl_69_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_6_to_mem      (ppe_stm_ppe_stm_mod_tbl_6_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_70_to_mem     (ppe_stm_ppe_stm_mod_tbl_70_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_71_to_mem     (ppe_stm_ppe_stm_mod_tbl_71_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_72_to_mem     (ppe_stm_ppe_stm_mod_tbl_72_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_73_to_mem     (ppe_stm_ppe_stm_mod_tbl_73_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_74_to_mem     (ppe_stm_ppe_stm_mod_tbl_74_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_75_to_mem     (ppe_stm_ppe_stm_mod_tbl_75_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_76_to_mem     (ppe_stm_ppe_stm_mod_tbl_76_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_77_to_mem     (ppe_stm_ppe_stm_mod_tbl_77_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_78_to_mem     (ppe_stm_ppe_stm_mod_tbl_78_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_79_to_mem     (ppe_stm_ppe_stm_mod_tbl_79_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_7_to_mem      (ppe_stm_ppe_stm_mod_tbl_7_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_8_to_mem      (ppe_stm_ppe_stm_mod_tbl_8_to_mem),                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_9_to_mem      (ppe_stm_ppe_stm_mod_tbl_9_to_mem),                
/* input  logic   [63:0] */ .ppe_stm_ppe_stm_shcp_tbl_to_mem       (ppe_stm_ppe_stm_shcp_tbl_to_mem),                 
/* input  logic          */ .cclk                                  (cclk),                                            
/* input  logic          */ .fary_enblfloat_sram                   (),                                                
/* input  logic          */ .fary_ensleep_sram                     (),                                                
/* input  logic          */ .car_raw_lan_power_good_with_byprst    (),                                                
/* input  logic   [19:0] */ .fary_ffuse_data_misc_sram             (),                                                
/* input  logic    [1:0] */ .fary_fwen_sram                        (),                                                
/* input  logic          */ .fary_pwren_b_sram                     (),                                                
/* input  logic          */ .fary_stm_enable                       (),                                                
/* input  logic          */ .fary_stm_hilo                         (),                                                
/* input  logic          */ .fary_wakeup_sram                      (),                                                
/* input  logic          */ .fdfx_lbist_test_mode                  (),                                                
/* input  logic          */ .fscan_byprst_b                        (),                                                
/* input  logic          */ .fscan_mode                            (),                                                
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_164_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_164_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_165_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_165_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_166_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_166_to_mem),             
/* input  logic   [92:0] */ .ppe_stm_ppe_stm_fwd_tbl0_167_to_mem   (ppe_stm_ppe_stm_fwd_tbl0_167_to_mem),             
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_64_to_mem     (ppe_stm_ppe_stm_mod_tbl_64_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_65_to_mem     (ppe_stm_ppe_stm_mod_tbl_65_to_mem),               
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_mod_tbl_66_to_mem     (ppe_stm_ppe_stm_mod_tbl_66_to_mem),               
/* input  logic  [337:0] */ .fscan_ram_awt_mode                    (),                                                
/* input  logic  [337:0] */ .fscan_ram_awt_ren                     (),                                                
/* input  logic  [337:0] */ .fscan_ram_awt_wen                     (),                                                
/* input  logic  [337:0] */ .fscan_ram_bypsel                      (),                                                
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_11_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_11_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_12_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_12_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_13_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_13_to_mem),              
/* input  logic   [91:0] */ .ppe_stm_ppe_stm_fwd_tbl1_14_to_mem    (ppe_stm_ppe_stm_fwd_tbl1_14_to_mem),              
/* output logic          */ .aary_pwren_b_sram                     (),                                                
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_0_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_0_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_100_from_mem (ppe_stm_ppe_stm_fwd_tbl0_100_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_101_from_mem (ppe_stm_ppe_stm_fwd_tbl0_101_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_102_from_mem (ppe_stm_ppe_stm_fwd_tbl0_102_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_103_from_mem (ppe_stm_ppe_stm_fwd_tbl0_103_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_104_from_mem (ppe_stm_ppe_stm_fwd_tbl0_104_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_105_from_mem (ppe_stm_ppe_stm_fwd_tbl0_105_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_106_from_mem (ppe_stm_ppe_stm_fwd_tbl0_106_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_107_from_mem (ppe_stm_ppe_stm_fwd_tbl0_107_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_108_from_mem (ppe_stm_ppe_stm_fwd_tbl0_108_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_109_from_mem (ppe_stm_ppe_stm_fwd_tbl0_109_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_10_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_10_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_110_from_mem (ppe_stm_ppe_stm_fwd_tbl0_110_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_111_from_mem (ppe_stm_ppe_stm_fwd_tbl0_111_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_112_from_mem (ppe_stm_ppe_stm_fwd_tbl0_112_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_113_from_mem (ppe_stm_ppe_stm_fwd_tbl0_113_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_114_from_mem (ppe_stm_ppe_stm_fwd_tbl0_114_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_115_from_mem (ppe_stm_ppe_stm_fwd_tbl0_115_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_116_from_mem (ppe_stm_ppe_stm_fwd_tbl0_116_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_117_from_mem (ppe_stm_ppe_stm_fwd_tbl0_117_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_118_from_mem (ppe_stm_ppe_stm_fwd_tbl0_118_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_119_from_mem (ppe_stm_ppe_stm_fwd_tbl0_119_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_11_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_11_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_120_from_mem (ppe_stm_ppe_stm_fwd_tbl0_120_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_121_from_mem (ppe_stm_ppe_stm_fwd_tbl0_121_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_122_from_mem (ppe_stm_ppe_stm_fwd_tbl0_122_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_123_from_mem (ppe_stm_ppe_stm_fwd_tbl0_123_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_124_from_mem (ppe_stm_ppe_stm_fwd_tbl0_124_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_125_from_mem (ppe_stm_ppe_stm_fwd_tbl0_125_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_126_from_mem (ppe_stm_ppe_stm_fwd_tbl0_126_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_127_from_mem (ppe_stm_ppe_stm_fwd_tbl0_127_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_128_from_mem (ppe_stm_ppe_stm_fwd_tbl0_128_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_129_from_mem (ppe_stm_ppe_stm_fwd_tbl0_129_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_12_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_12_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_130_from_mem (ppe_stm_ppe_stm_fwd_tbl0_130_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_131_from_mem (ppe_stm_ppe_stm_fwd_tbl0_131_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_132_from_mem (ppe_stm_ppe_stm_fwd_tbl0_132_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_133_from_mem (ppe_stm_ppe_stm_fwd_tbl0_133_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_134_from_mem (ppe_stm_ppe_stm_fwd_tbl0_134_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_135_from_mem (ppe_stm_ppe_stm_fwd_tbl0_135_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_136_from_mem (ppe_stm_ppe_stm_fwd_tbl0_136_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_137_from_mem (ppe_stm_ppe_stm_fwd_tbl0_137_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_138_from_mem (ppe_stm_ppe_stm_fwd_tbl0_138_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_139_from_mem (ppe_stm_ppe_stm_fwd_tbl0_139_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_13_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_13_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_140_from_mem (ppe_stm_ppe_stm_fwd_tbl0_140_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_141_from_mem (ppe_stm_ppe_stm_fwd_tbl0_141_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_142_from_mem (ppe_stm_ppe_stm_fwd_tbl0_142_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_143_from_mem (ppe_stm_ppe_stm_fwd_tbl0_143_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_144_from_mem (ppe_stm_ppe_stm_fwd_tbl0_144_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_145_from_mem (ppe_stm_ppe_stm_fwd_tbl0_145_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_146_from_mem (ppe_stm_ppe_stm_fwd_tbl0_146_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_147_from_mem (ppe_stm_ppe_stm_fwd_tbl0_147_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_148_from_mem (ppe_stm_ppe_stm_fwd_tbl0_148_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_149_from_mem (ppe_stm_ppe_stm_fwd_tbl0_149_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_14_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_14_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_150_from_mem (ppe_stm_ppe_stm_fwd_tbl0_150_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_151_from_mem (ppe_stm_ppe_stm_fwd_tbl0_151_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_152_from_mem (ppe_stm_ppe_stm_fwd_tbl0_152_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_153_from_mem (ppe_stm_ppe_stm_fwd_tbl0_153_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_154_from_mem (ppe_stm_ppe_stm_fwd_tbl0_154_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_155_from_mem (ppe_stm_ppe_stm_fwd_tbl0_155_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_156_from_mem (ppe_stm_ppe_stm_fwd_tbl0_156_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_157_from_mem (ppe_stm_ppe_stm_fwd_tbl0_157_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_158_from_mem (ppe_stm_ppe_stm_fwd_tbl0_158_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_159_from_mem (ppe_stm_ppe_stm_fwd_tbl0_159_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_15_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_15_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_160_from_mem (ppe_stm_ppe_stm_fwd_tbl0_160_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_161_from_mem (ppe_stm_ppe_stm_fwd_tbl0_161_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_162_from_mem (ppe_stm_ppe_stm_fwd_tbl0_162_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_163_from_mem (ppe_stm_ppe_stm_fwd_tbl0_163_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_164_from_mem (ppe_stm_ppe_stm_fwd_tbl0_164_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_165_from_mem (ppe_stm_ppe_stm_fwd_tbl0_165_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_166_from_mem (ppe_stm_ppe_stm_fwd_tbl0_166_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_167_from_mem (ppe_stm_ppe_stm_fwd_tbl0_167_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_168_from_mem (ppe_stm_ppe_stm_fwd_tbl0_168_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_169_from_mem (ppe_stm_ppe_stm_fwd_tbl0_169_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_16_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_16_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_170_from_mem (ppe_stm_ppe_stm_fwd_tbl0_170_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_171_from_mem (ppe_stm_ppe_stm_fwd_tbl0_171_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_172_from_mem (ppe_stm_ppe_stm_fwd_tbl0_172_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_173_from_mem (ppe_stm_ppe_stm_fwd_tbl0_173_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_174_from_mem (ppe_stm_ppe_stm_fwd_tbl0_174_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_175_from_mem (ppe_stm_ppe_stm_fwd_tbl0_175_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_176_from_mem (ppe_stm_ppe_stm_fwd_tbl0_176_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_177_from_mem (ppe_stm_ppe_stm_fwd_tbl0_177_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_178_from_mem (ppe_stm_ppe_stm_fwd_tbl0_178_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_179_from_mem (ppe_stm_ppe_stm_fwd_tbl0_179_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_17_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_17_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_180_from_mem (ppe_stm_ppe_stm_fwd_tbl0_180_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_181_from_mem (ppe_stm_ppe_stm_fwd_tbl0_181_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_182_from_mem (ppe_stm_ppe_stm_fwd_tbl0_182_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_183_from_mem (ppe_stm_ppe_stm_fwd_tbl0_183_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_184_from_mem (ppe_stm_ppe_stm_fwd_tbl0_184_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_185_from_mem (ppe_stm_ppe_stm_fwd_tbl0_185_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_186_from_mem (ppe_stm_ppe_stm_fwd_tbl0_186_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_187_from_mem (ppe_stm_ppe_stm_fwd_tbl0_187_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_188_from_mem (ppe_stm_ppe_stm_fwd_tbl0_188_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_189_from_mem (ppe_stm_ppe_stm_fwd_tbl0_189_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_18_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_18_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_190_from_mem (ppe_stm_ppe_stm_fwd_tbl0_190_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_20_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_20_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_21_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_21_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_22_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_22_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_23_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_23_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_24_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_24_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_25_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_25_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_26_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_26_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_27_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_27_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_28_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_28_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_29_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_29_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_2_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_2_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_30_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_30_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_31_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_31_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_32_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_32_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_33_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_33_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_34_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_34_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_35_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_35_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_36_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_36_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_37_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_37_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_38_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_38_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_39_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_39_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_3_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_3_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_40_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_40_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_41_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_41_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_42_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_42_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_43_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_43_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_44_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_44_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_45_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_45_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_46_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_46_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_47_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_47_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_48_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_48_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_49_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_49_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_4_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_4_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_50_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_50_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_51_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_51_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_52_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_52_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_53_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_53_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_54_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_54_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_55_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_55_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_56_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_56_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_57_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_57_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_58_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_58_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_59_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_59_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_5_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_5_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_60_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_60_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_61_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_61_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_62_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_62_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_63_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_63_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_64_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_64_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_65_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_65_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_66_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_66_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_67_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_67_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_68_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_68_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_69_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_69_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_6_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_6_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_70_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_70_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_71_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_71_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_72_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_72_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_73_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_73_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_74_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_74_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_75_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_75_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_76_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_76_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_77_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_77_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_78_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_78_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_79_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_79_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_7_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_7_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_80_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_80_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_81_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_81_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_82_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_82_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_83_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_83_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_84_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_84_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_85_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_85_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_86_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_86_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_87_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_87_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_88_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_88_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_89_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_89_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_8_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_8_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_90_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_90_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_91_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_91_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_92_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_92_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_93_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_93_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_94_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_94_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_95_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_95_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_96_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_96_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_97_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_97_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_98_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_98_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_99_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_99_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_9_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_9_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_0_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_0_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_10_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_10_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_11_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_11_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_12_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_12_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_13_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_13_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_14_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_14_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_15_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_15_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_16_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_16_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_17_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_17_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_18_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_18_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_19_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_19_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_1_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_1_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_20_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_20_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_21_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_21_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_22_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_22_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_23_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_23_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_24_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_24_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_25_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_25_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_26_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_26_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_27_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_27_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_28_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_28_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_29_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_29_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_2_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_2_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_30_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_30_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_31_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_31_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_32_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_32_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_33_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_33_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_34_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_34_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_35_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_35_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_36_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_36_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_37_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_37_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_38_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_38_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_39_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_39_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_3_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_3_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_40_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_40_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_41_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_41_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_42_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_42_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_43_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_43_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_44_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_44_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_49_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_49_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_4_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_4_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_50_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_50_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_51_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_51_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_52_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_52_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_53_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_53_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_54_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_54_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_55_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_55_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_56_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_56_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_57_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_57_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_58_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_58_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_59_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_59_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_5_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_5_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_60_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_60_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_61_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_61_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_62_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_62_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_63_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_63_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_6_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_6_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_7_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_7_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_8_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_8_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_9_from_mem   (ppe_stm_ppe_stm_fwd_tbl1_9_from_mem),             
/* output logic  [576:0] */ .ppe_stm_ppe_stm_l3mc_tbl_from_mem     (ppe_stm_ppe_stm_l3mc_tbl_from_mem),               
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_0_from_mem    (ppe_stm_ppe_stm_mod_tbl_0_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_10_from_mem   (ppe_stm_ppe_stm_mod_tbl_10_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_11_from_mem   (ppe_stm_ppe_stm_mod_tbl_11_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_12_from_mem   (ppe_stm_ppe_stm_mod_tbl_12_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_13_from_mem   (ppe_stm_ppe_stm_mod_tbl_13_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_14_from_mem   (ppe_stm_ppe_stm_mod_tbl_14_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_15_from_mem   (ppe_stm_ppe_stm_mod_tbl_15_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_16_from_mem   (ppe_stm_ppe_stm_mod_tbl_16_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_17_from_mem   (ppe_stm_ppe_stm_mod_tbl_17_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_18_from_mem   (ppe_stm_ppe_stm_mod_tbl_18_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_19_from_mem   (ppe_stm_ppe_stm_mod_tbl_19_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_1_from_mem    (ppe_stm_ppe_stm_mod_tbl_1_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_20_from_mem   (ppe_stm_ppe_stm_mod_tbl_20_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_21_from_mem   (ppe_stm_ppe_stm_mod_tbl_21_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_22_from_mem   (ppe_stm_ppe_stm_mod_tbl_22_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_23_from_mem   (ppe_stm_ppe_stm_mod_tbl_23_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_24_from_mem   (ppe_stm_ppe_stm_mod_tbl_24_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_25_from_mem   (ppe_stm_ppe_stm_mod_tbl_25_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_26_from_mem   (ppe_stm_ppe_stm_mod_tbl_26_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_27_from_mem   (ppe_stm_ppe_stm_mod_tbl_27_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_28_from_mem   (ppe_stm_ppe_stm_mod_tbl_28_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_29_from_mem   (ppe_stm_ppe_stm_mod_tbl_29_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_2_from_mem    (ppe_stm_ppe_stm_mod_tbl_2_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_30_from_mem   (ppe_stm_ppe_stm_mod_tbl_30_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_31_from_mem   (ppe_stm_ppe_stm_mod_tbl_31_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_32_from_mem   (ppe_stm_ppe_stm_mod_tbl_32_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_33_from_mem   (ppe_stm_ppe_stm_mod_tbl_33_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_34_from_mem   (ppe_stm_ppe_stm_mod_tbl_34_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_35_from_mem   (ppe_stm_ppe_stm_mod_tbl_35_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_36_from_mem   (ppe_stm_ppe_stm_mod_tbl_36_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_37_from_mem   (ppe_stm_ppe_stm_mod_tbl_37_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_38_from_mem   (ppe_stm_ppe_stm_mod_tbl_38_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_39_from_mem   (ppe_stm_ppe_stm_mod_tbl_39_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_3_from_mem    (ppe_stm_ppe_stm_mod_tbl_3_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_40_from_mem   (ppe_stm_ppe_stm_mod_tbl_40_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_41_from_mem   (ppe_stm_ppe_stm_mod_tbl_41_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_42_from_mem   (ppe_stm_ppe_stm_mod_tbl_42_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_43_from_mem   (ppe_stm_ppe_stm_mod_tbl_43_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_44_from_mem   (ppe_stm_ppe_stm_mod_tbl_44_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_45_from_mem   (ppe_stm_ppe_stm_mod_tbl_45_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_46_from_mem   (ppe_stm_ppe_stm_mod_tbl_46_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_47_from_mem   (ppe_stm_ppe_stm_mod_tbl_47_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_48_from_mem   (ppe_stm_ppe_stm_mod_tbl_48_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_49_from_mem   (ppe_stm_ppe_stm_mod_tbl_49_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_4_from_mem    (ppe_stm_ppe_stm_mod_tbl_4_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_50_from_mem   (ppe_stm_ppe_stm_mod_tbl_50_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_51_from_mem   (ppe_stm_ppe_stm_mod_tbl_51_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_52_from_mem   (ppe_stm_ppe_stm_mod_tbl_52_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_53_from_mem   (ppe_stm_ppe_stm_mod_tbl_53_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_54_from_mem   (ppe_stm_ppe_stm_mod_tbl_54_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_55_from_mem   (ppe_stm_ppe_stm_mod_tbl_55_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_56_from_mem   (ppe_stm_ppe_stm_mod_tbl_56_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_57_from_mem   (ppe_stm_ppe_stm_mod_tbl_57_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_58_from_mem   (ppe_stm_ppe_stm_mod_tbl_58_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_59_from_mem   (ppe_stm_ppe_stm_mod_tbl_59_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_5_from_mem    (ppe_stm_ppe_stm_mod_tbl_5_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_60_from_mem   (ppe_stm_ppe_stm_mod_tbl_60_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_61_from_mem   (ppe_stm_ppe_stm_mod_tbl_61_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_62_from_mem   (ppe_stm_ppe_stm_mod_tbl_62_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_63_from_mem   (ppe_stm_ppe_stm_mod_tbl_63_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_64_from_mem   (ppe_stm_ppe_stm_mod_tbl_64_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_65_from_mem   (ppe_stm_ppe_stm_mod_tbl_65_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_66_from_mem   (ppe_stm_ppe_stm_mod_tbl_66_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_67_from_mem   (ppe_stm_ppe_stm_mod_tbl_67_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_68_from_mem   (ppe_stm_ppe_stm_mod_tbl_68_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_69_from_mem   (ppe_stm_ppe_stm_mod_tbl_69_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_6_from_mem    (ppe_stm_ppe_stm_mod_tbl_6_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_70_from_mem   (ppe_stm_ppe_stm_mod_tbl_70_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_71_from_mem   (ppe_stm_ppe_stm_mod_tbl_71_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_72_from_mem   (ppe_stm_ppe_stm_mod_tbl_72_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_73_from_mem   (ppe_stm_ppe_stm_mod_tbl_73_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_74_from_mem   (ppe_stm_ppe_stm_mod_tbl_74_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_75_from_mem   (ppe_stm_ppe_stm_mod_tbl_75_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_76_from_mem   (ppe_stm_ppe_stm_mod_tbl_76_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_77_from_mem   (ppe_stm_ppe_stm_mod_tbl_77_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_78_from_mem   (ppe_stm_ppe_stm_mod_tbl_78_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_79_from_mem   (ppe_stm_ppe_stm_mod_tbl_79_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_7_from_mem    (ppe_stm_ppe_stm_mod_tbl_7_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_8_from_mem    (ppe_stm_ppe_stm_mod_tbl_8_from_mem),              
/* output logic   [72:0] */ .ppe_stm_ppe_stm_mod_tbl_9_from_mem    (ppe_stm_ppe_stm_mod_tbl_9_from_mem),              
/* output logic   [40:0] */ .ppe_stm_ppe_stm_shcp_tbl_from_mem     (ppe_stm_ppe_stm_shcp_tbl_from_mem),               
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_191_from_mem (ppe_stm_ppe_stm_fwd_tbl0_191_from_mem),           
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_19_from_mem  (ppe_stm_ppe_stm_fwd_tbl0_19_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl0_1_from_mem   (ppe_stm_ppe_stm_fwd_tbl0_1_from_mem),             
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_45_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_45_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_46_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_46_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_47_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_47_from_mem),            
/* output logic   [72:0] */ .ppe_stm_ppe_stm_fwd_tbl1_48_from_mem  (ppe_stm_ppe_stm_fwd_tbl1_48_from_mem));            
// End of module ppe_stm_sram_mems from ppe_stm_sram_mems

endmodule // ppe_stm_top
