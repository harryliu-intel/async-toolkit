magic
tech scmos
timestamp 970030343
<< ndiffusion >>
rect -25 148 -9 149
rect -25 140 -9 145
rect -25 132 -9 137
rect -25 124 -9 129
rect -50 117 -46 122
rect -58 116 -46 117
rect -25 120 -9 121
rect -58 108 -46 113
rect -25 111 -9 112
rect -58 103 -46 105
rect -50 95 -46 103
rect -25 103 -9 108
rect -25 95 -9 100
rect -58 94 -46 95
rect -58 90 -46 91
rect -50 82 -46 90
rect -25 87 -9 92
rect -58 81 -46 82
rect -25 83 -9 84
rect -58 73 -46 78
rect -25 74 -9 75
rect -58 69 -46 70
rect -58 61 -56 69
rect -58 59 -46 61
rect -58 55 -46 56
<< pdiffusion >>
rect 21 150 52 151
rect 66 151 74 156
rect 58 150 74 151
rect 21 146 52 147
rect 44 138 52 146
rect 21 137 52 138
rect 58 146 74 147
rect 58 138 66 146
rect 58 137 74 138
rect 21 133 52 134
rect 21 124 52 125
rect 58 133 74 134
rect 66 125 74 133
rect 58 124 74 125
rect 21 120 52 121
rect 58 120 74 121
rect 58 112 64 120
rect 72 112 74 120
rect 58 111 74 112
rect 58 107 74 108
rect 21 98 37 99
rect 72 99 74 107
rect 58 98 74 99
rect 21 94 37 95
rect 21 86 29 94
rect 58 92 74 95
rect 58 88 71 92
rect 21 85 37 86
rect 21 81 37 82
rect 21 72 37 73
rect 59 73 67 78
rect 51 72 67 73
rect 21 68 37 69
rect 51 68 67 69
rect 21 59 37 60
<< ntransistor >>
rect -25 145 -9 148
rect -25 137 -9 140
rect -25 129 -9 132
rect -25 121 -9 124
rect -58 113 -46 116
rect -25 108 -9 111
rect -58 105 -46 108
rect -25 100 -9 103
rect -58 91 -46 94
rect -25 92 -9 95
rect -58 78 -46 81
rect -25 84 -9 87
rect -58 70 -46 73
rect -58 56 -46 59
<< ptransistor >>
rect 21 147 52 150
rect 58 147 74 150
rect 21 134 52 137
rect 58 134 74 137
rect 21 121 52 124
rect 58 121 74 124
rect 58 108 74 111
rect 21 95 37 98
rect 58 95 74 98
rect 21 82 37 85
rect 21 69 37 72
rect 51 69 67 72
<< polysilicon >>
rect -29 145 -25 148
rect -9 145 -5 148
rect 8 147 21 150
rect 52 147 58 150
rect 74 147 78 150
rect 8 140 11 147
rect -55 137 -25 140
rect -9 137 11 140
rect 16 134 21 137
rect 52 134 58 137
rect 74 134 78 137
rect 16 132 19 134
rect -63 116 -60 132
rect -36 129 -25 132
rect -9 129 19 132
rect -29 121 -25 124
rect -9 121 -4 124
rect -63 113 -58 116
rect -46 113 -28 116
rect -31 111 -28 113
rect 4 121 21 124
rect 52 121 58 124
rect 74 121 78 124
rect -31 108 -25 111
rect -9 108 19 111
rect 54 108 58 111
rect 74 108 76 111
rect -62 105 -58 108
rect -46 105 -44 108
rect -36 100 -25 103
rect -9 100 11 103
rect -43 94 -25 95
rect -62 91 -58 94
rect -46 92 -25 94
rect -9 92 3 95
rect -46 91 -39 92
rect -33 86 -25 87
rect -62 78 -58 81
rect -46 78 -38 81
rect -30 84 -25 86
rect -9 84 -5 87
rect 0 77 3 92
rect 8 85 11 100
rect 16 98 19 108
rect 16 95 21 98
rect 37 95 41 98
rect 54 95 58 98
rect 74 95 78 98
rect 8 82 21 85
rect 37 82 41 85
rect 0 74 4 77
rect -60 70 -58 73
rect -46 70 -42 73
rect 12 69 21 72
rect 37 69 41 72
rect 47 69 51 72
rect 67 69 74 72
rect 71 67 74 69
rect -62 56 -58 59
rect -46 57 -39 59
rect -46 56 -42 57
<< ndcontact >>
rect -25 149 -9 157
rect -58 117 -50 125
rect -25 112 -9 120
rect -58 95 -50 103
rect -58 82 -50 90
rect -25 75 -9 83
rect -56 61 -46 69
rect -58 47 -46 55
<< pdcontact >>
rect 21 151 52 159
rect 58 151 66 159
rect 21 138 44 146
rect 66 138 74 146
rect 21 125 52 133
rect 58 125 66 133
rect 21 112 52 120
rect 64 112 72 120
rect 21 99 37 107
rect 58 99 72 107
rect 29 86 37 94
rect 71 84 79 92
rect 21 73 37 81
rect 51 73 59 81
rect 21 60 37 68
rect 51 60 67 68
<< psubstratepcontact >>
rect -25 66 -9 74
<< nsubstratencontact >>
rect 21 51 37 59
<< polycontact >>
rect -37 145 -29 153
rect -63 132 -55 140
rect -44 124 -36 132
rect -4 116 4 124
rect -44 100 -36 108
rect -38 78 -30 86
rect 76 103 84 111
rect 46 90 54 98
rect -68 65 -60 73
rect 4 69 12 77
rect 71 59 79 67
rect -42 49 -34 57
<< metal1 >>
rect -37 145 -29 155
rect -25 155 -21 157
rect -25 149 -9 155
rect 10 146 16 155
rect 21 151 52 159
rect -63 132 -55 143
rect 10 138 44 146
rect 48 133 52 151
rect -58 121 -50 125
rect -66 117 -50 121
rect -66 90 -62 117
rect -58 95 -50 107
rect -44 100 -36 131
rect 21 125 52 133
rect 56 151 66 159
rect 56 133 60 151
rect 66 138 74 146
rect 56 125 66 133
rect -25 113 -9 120
rect 56 120 60 125
rect 70 120 74 138
rect 4 119 8 120
rect -4 116 8 119
rect -13 103 -9 107
rect -13 99 0 103
rect -66 86 -50 90
rect -58 82 -50 86
rect -38 78 -30 83
rect -68 65 -60 71
rect -25 69 -9 83
rect -65 55 -60 65
rect -56 65 -9 69
rect -56 61 -21 65
rect -42 55 -34 57
rect -4 55 0 99
rect 4 77 8 116
rect 21 113 60 120
rect 64 116 74 120
rect 21 112 41 113
rect 64 112 72 116
rect 21 99 37 107
rect 21 81 25 99
rect 46 94 54 107
rect 58 99 72 107
rect 76 103 84 111
rect 29 86 55 94
rect 51 81 55 86
rect 4 69 12 77
rect 21 73 37 81
rect 51 73 59 81
rect 63 68 67 99
rect 76 92 81 103
rect 71 84 81 92
rect 76 77 81 84
rect 21 60 67 68
rect 71 65 79 67
rect -65 50 -46 55
rect -58 47 -46 50
rect -42 51 0 55
rect 21 51 37 60
rect -42 49 -34 51
<< m2contact >>
rect -37 155 -29 161
rect -63 143 -55 149
rect -21 155 -3 161
rect 3 155 16 161
rect -44 131 -36 137
rect -58 107 -50 113
rect -4 119 4 125
rect -25 107 -9 113
rect -38 83 -30 89
rect -68 71 -60 77
rect -21 59 -9 65
rect 41 107 54 113
rect 73 71 81 77
rect 8 59 21 65
rect 71 59 79 65
<< metal2 >>
rect -37 155 -26 161
rect -63 143 0 149
rect -44 131 0 137
rect -6 119 6 125
rect -58 107 54 113
rect -38 83 -27 89
rect -68 71 81 77
rect 27 59 79 65
<< m3contact >>
rect -21 155 -3 161
rect 3 155 21 161
rect -21 59 -3 65
rect 3 59 21 65
<< metal3 >>
rect -21 44 -3 164
rect 3 44 21 164
<< labels >>
rlabel polysilicon 75 122 75 122 1 a
rlabel polysilicon 38 70 38 70 1 a
rlabel metal1 33 90 33 90 1 x
rlabel metal1 29 64 29 64 1 Vdd!
rlabel metal1 -13 79 -13 79 1 GND!
rlabel metal1 -13 153 -13 153 5 GND!
rlabel metal1 58 64 58 64 1 Vdd!
rlabel polysilicon 68 70 68 70 1 _PReset!
rlabel metal1 67 103 67 103 1 Vdd!
rlabel polysilicon -26 138 -26 138 1 _b1
rlabel polysilicon -26 130 -26 130 1 _b0
rlabel polysilicon -26 146 -26 146 1 _SReset!
rlabel metal1 -13 116 -13 116 5 x
rlabel metal1 33 116 33 116 1 x
rlabel metal2 0 119 0 125 1 a
rlabel metal2 75 62 75 62 1 _PReset!
rlabel polysilicon -59 79 -59 79 1 _SReset!
rlabel metal1 -52 65 -52 65 1 GND!
rlabel polysilicon -59 114 -59 114 1 _b1
rlabel polysilicon -59 106 -59 106 1 _b0
rlabel metal1 -54 99 -54 99 1 x
rlabel metal2 0 131 0 137 7 _b0
rlabel metal2 0 143 0 149 7 _b1
rlabel metal2 -34 86 -34 86 1 _SReset!
rlabel metal2 -33 158 -33 158 1 _SReset!
rlabel metal1 40 142 40 142 1 Vdd!
rlabel metal1 62 155 62 155 5 x
rlabel metal1 62 129 62 129 1 x
rlabel space 36 50 85 160 3 ^p
rlabel space -69 47 -24 162 7 ^n
rlabel metal2 -27 83 -27 89 3 ^n
rlabel metal2 -26 155 -26 161 3 ^n
rlabel metal2 -54 110 -54 110 1 x
rlabel metal2 -59 146 -59 146 1 _b1
rlabel metal2 -40 134 -40 134 1 _b0
rlabel metal2 48 110 48 110 1 x
rlabel metal2 0 107 0 113 1 x
<< end >>
