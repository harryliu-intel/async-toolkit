    package svt_ahb_bfm_pkg;

        import sla_pkg::*;
        `include "uvm_macros.svh"
        `include "slu_macros.svh"
        import svt_uvm_pkg::*;
        import uvm_pkg::*;
        import svt_ahb_uvm_pkg::*;
        
        import svt_amba_common_uvm_pkg::*;

        
        `include "cust_svt_ahb_system_configuration.sv"
        `include "cust_svt_master_transaction.sv"
        `include "cust_svt_ahb_slave_transaction.sv"
        `include "ahb_virtual_sequencer.sv"
        `include "ahb_slave_random_response_sequence.sv"
        `include "ahb_master_directed_sequence.sv"
        `include "ahb_bfm_env.sv"

    endpackage


