//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2021 - 2021 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related
// to the source code ("Material") are owned by Intel Corporation or its
// suppliers or licensors. Title to the Material remains with Intel
// Corporation or its suppliers and licensors. The Material contains trade
// secrets and proprietary and confidential information of Intel or its
// suppliers and licensors. The Material is protected by worldwide copyright
// and trade secret laws and treaty provisions. No part of the Material may
// be used, copied, reproduced, modified, published, uploaded, posted,
// transmitted, distributed, or disclosed in any way without Intel's prior
// express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or
// delivery of the Materials, either expressly, by implication, inducement,
// estoppel or otherwise. Any license under such intellectual property rights
// must be express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//
// LATCH primitive
//
// Author : mika.nystroem@intel.com
// April, 2022
//


`resetall
`default_nettype wire  // needed for primitive?

`ifndef _LATCH_SV
`define _LATCH_SV

primitive LATCH( Q, CK, D );
   output     Q;
   reg        Q;
   input      CK;
   input      D;
table
//     CK  D  :  Q  :  Q
        0  ?  :  ?  :  -;
        1  1  :  ?  :  1;
        ?  1  :  1  :  1;
        1  0  :  ?  :  0;
        ?  0  :  0  :  0;

endtable
endprimitive

`endif // !_LATCH_SV

`default_nettype none
`default_nettype wire
