magic
tech scmos
timestamp 982687028
<< nselect >>
rect -50 58 0 96
rect -32 11 0 53
<< pselect >>
rect 0 58 62 95
rect 0 19 32 53
<< ndiffusion >>
rect -46 82 -42 85
rect -16 81 -8 82
rect -16 77 -8 78
rect -46 72 -42 77
rect -46 66 -42 69
rect -28 44 -8 45
rect -28 36 -8 41
rect -28 28 -8 33
rect -28 24 -8 25
<< pdiffusion >>
rect 54 82 58 87
rect 8 81 16 82
rect 8 77 16 78
rect 23 73 27 82
rect 46 81 58 82
rect 46 77 58 78
rect 54 72 58 77
rect 23 66 27 69
rect 8 44 28 45
rect 8 36 28 41
rect 8 32 28 33
<< ntransistor >>
rect -46 77 -42 82
rect -16 78 -8 81
rect -46 69 -42 72
rect -28 41 -8 44
rect -28 33 -8 36
rect -28 25 -8 28
<< ptransistor >>
rect 8 78 16 81
rect 46 78 58 81
rect 23 69 27 73
rect 8 41 28 44
rect 8 33 28 36
<< polysilicon >>
rect -50 77 -46 82
rect -42 77 -38 82
rect -20 78 -16 81
rect -8 78 -4 81
rect -50 69 -46 72
rect -42 69 -33 72
rect 4 78 8 81
rect 16 78 20 81
rect 42 78 46 81
rect 58 78 62 81
rect 18 69 23 73
rect 27 70 29 73
rect 27 69 31 70
rect 18 67 21 69
rect -28 64 21 67
rect -32 41 -28 44
rect -8 41 8 44
rect 28 41 32 44
rect -32 33 -28 36
rect -8 33 8 36
rect 28 33 32 36
rect -32 25 -28 28
rect -8 25 -4 28
<< ndcontact >>
rect -50 85 -42 93
rect -16 82 -8 90
rect -16 69 -8 77
rect -50 58 -42 66
rect -28 45 -8 53
rect -28 16 -8 24
<< pdcontact >>
rect 8 82 16 90
rect 22 82 30 90
rect 46 82 54 90
rect 8 69 16 77
rect 46 69 54 77
rect 23 58 31 66
rect 8 45 28 53
rect 8 24 28 32
<< polycontact >>
rect -33 67 -25 75
rect -4 73 4 81
rect 29 70 37 78
<< metal1 >>
rect -50 90 -42 93
rect -50 88 -8 90
rect -50 85 -27 88
rect -9 82 -8 88
rect 8 88 54 90
rect 8 82 9 88
rect 27 82 54 88
rect -16 75 -8 77
rect -33 71 -8 75
rect -33 67 -25 71
rect -16 69 -8 71
rect -50 62 -42 66
rect -4 62 4 81
rect 8 75 16 77
rect 29 75 37 78
rect 8 71 37 75
rect 8 69 16 71
rect 29 70 37 71
rect 46 69 54 77
rect 46 66 50 69
rect 23 62 50 66
rect -50 58 31 62
rect -4 53 4 58
rect -28 46 28 53
rect -28 45 -8 46
rect 8 45 28 46
rect 8 24 28 32
rect -28 19 -8 24
rect -28 16 -27 19
rect -9 16 -8 19
rect 9 19 27 24
<< m2contact >>
rect -27 82 -9 88
rect 9 82 27 88
rect -27 13 -9 19
rect 9 13 27 19
<< m3contact >>
rect -27 82 -9 88
rect 9 82 27 88
rect -27 13 -9 19
rect 9 13 27 19
<< metal3 >>
rect -27 11 -9 96
rect 9 11 27 96
<< labels >>
rlabel metal1 -46 63 -46 63 3 x
rlabel space -33 11 -28 53 7 ^n
rlabel space 28 19 33 53 3 ^p
rlabel metal3 -27 11 -9 96 1 GND!|pin|s|0
rlabel metal3 9 11 27 96 1 Vdd!|pin|s|1
rlabel metal1 -28 16 -8 24 1 GND!|pin|s|0
rlabel metal1 -50 85 -8 90 1 GND!|pin|s|0
rlabel metal1 8 82 54 90 1 Vdd!|pin|s|1
rlabel metal1 8 24 28 32 1 Vdd!|pin|s|1
rlabel metal1 9 13 27 32 1 Vdd!|pin|s|1
rlabel metal1 -4 46 4 81 1 x|pin|s|2
rlabel metal1 -28 46 28 53 1 x|pin|s|2
rlabel polysilicon 28 33 32 36 1 a|pin|w|3|poly
rlabel polysilicon 0 33 4 36 1 a|pin|w|3|poly
rlabel polysilicon -32 33 -28 36 1 a|pin|w|3|poly
rlabel polysilicon -32 41 -28 44 1 b|pin|w|4|poly
rlabel polysilicon 28 41 32 44 1 b|pin|w|4|poly
rlabel polysilicon -32 25 -28 28 1 _SReset!|pin|w|5|poly
rlabel polysilicon -8 25 -4 28 1 _SReset!|pin|w|5|poly
rlabel polysilicon -50 77 -46 82 1 _SReset!|pin|w|6|poly
rlabel polysilicon -42 77 -38 82 1 _SReset!|pin|w|6|poly
rlabel polysilicon 42 78 46 81 1 _PReset!|pin|w|7|poly
rlabel polysilicon 58 78 62 81 1 _PReset!|pin|w|7|poly
<< end >>
