magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect -225 -698 -217 -697
rect -225 -706 -217 -701
rect -225 -714 -217 -709
rect -225 -722 -217 -717
rect -225 -730 -217 -725
rect -225 -738 -217 -733
rect -225 -742 -217 -741
rect -225 -751 -217 -750
rect -225 -759 -217 -754
rect -225 -767 -217 -762
rect -225 -775 -217 -770
rect -225 -783 -217 -778
rect -225 -791 -217 -786
rect -225 -795 -217 -794
<< pdiffusion >>
rect -194 -673 -186 -672
rect -194 -677 -186 -676
rect -194 -686 -186 -685
rect -194 -690 -186 -689
rect -194 -699 -186 -698
rect -194 -703 -186 -702
rect -194 -712 -186 -711
rect -194 -716 -186 -715
rect -194 -725 -186 -724
rect -194 -729 -186 -728
rect -194 -738 -186 -737
rect -194 -742 -186 -741
rect -194 -751 -186 -750
rect -194 -755 -186 -754
rect -194 -764 -186 -763
rect -194 -768 -186 -767
rect -194 -777 -186 -776
rect -194 -781 -186 -780
rect -194 -790 -186 -789
rect -194 -794 -186 -793
rect -194 -803 -186 -802
rect -194 -807 -186 -806
rect -194 -816 -186 -815
rect -194 -820 -186 -819
<< ntransistor >>
rect -225 -701 -217 -698
rect -225 -709 -217 -706
rect -225 -717 -217 -714
rect -225 -725 -217 -722
rect -225 -733 -217 -730
rect -225 -741 -217 -738
rect -225 -754 -217 -751
rect -225 -762 -217 -759
rect -225 -770 -217 -767
rect -225 -778 -217 -775
rect -225 -786 -217 -783
rect -225 -794 -217 -791
<< ptransistor >>
rect -194 -676 -186 -673
rect -194 -689 -186 -686
rect -194 -702 -186 -699
rect -194 -715 -186 -712
rect -194 -728 -186 -725
rect -194 -741 -186 -738
rect -194 -754 -186 -751
rect -194 -767 -186 -764
rect -194 -780 -186 -777
rect -194 -793 -186 -790
rect -194 -806 -186 -803
rect -194 -819 -186 -816
<< polysilicon >>
rect -215 -676 -194 -673
rect -186 -676 -182 -673
rect -215 -698 -212 -676
rect -229 -701 -225 -698
rect -217 -701 -212 -698
rect -199 -689 -194 -686
rect -186 -689 -182 -686
rect -199 -699 -196 -689
rect -207 -702 -194 -699
rect -186 -702 -182 -699
rect -207 -706 -204 -702
rect -229 -709 -225 -706
rect -217 -709 -204 -706
rect -199 -714 -194 -712
rect -229 -717 -225 -714
rect -217 -715 -194 -714
rect -186 -715 -182 -712
rect -217 -717 -196 -715
rect -229 -725 -225 -722
rect -217 -725 -196 -722
rect -199 -728 -194 -725
rect -186 -728 -182 -725
rect -229 -733 -225 -730
rect -217 -733 -213 -730
rect -229 -741 -225 -738
rect -217 -741 -194 -738
rect -186 -741 -182 -738
rect -229 -754 -225 -751
rect -217 -754 -194 -751
rect -186 -754 -182 -751
rect -229 -762 -225 -759
rect -217 -762 -213 -759
rect -199 -767 -194 -764
rect -186 -767 -182 -764
rect -229 -770 -225 -767
rect -217 -770 -196 -767
rect -229 -778 -225 -775
rect -217 -777 -196 -775
rect -217 -778 -194 -777
rect -199 -780 -194 -778
rect -186 -780 -182 -777
rect -229 -786 -225 -783
rect -217 -786 -204 -783
rect -207 -790 -204 -786
rect -229 -794 -225 -791
rect -217 -794 -212 -791
rect -207 -793 -194 -790
rect -186 -793 -182 -790
rect -215 -816 -212 -794
rect -199 -803 -196 -793
rect -199 -806 -194 -803
rect -186 -806 -182 -803
rect -215 -819 -194 -816
rect -186 -819 -182 -816
<< ndcontact >>
rect -225 -697 -217 -689
rect -225 -750 -217 -742
rect -225 -803 -217 -795
<< pdcontact >>
rect -194 -672 -186 -664
rect -194 -685 -186 -677
rect -194 -698 -186 -690
rect -194 -711 -186 -703
rect -194 -724 -186 -716
rect -194 -737 -186 -729
rect -194 -750 -186 -742
rect -194 -763 -186 -755
rect -194 -776 -186 -768
rect -194 -789 -186 -781
rect -194 -802 -186 -794
rect -194 -815 -186 -807
rect -194 -828 -186 -820
<< metal1 >>
rect -194 -672 -186 -664
rect -206 -685 -186 -677
rect -225 -697 -217 -689
rect -206 -703 -198 -685
rect -194 -698 -186 -690
rect -206 -711 -186 -703
rect -206 -729 -198 -711
rect -194 -724 -186 -716
rect -206 -737 -186 -729
rect -206 -742 -198 -737
rect -225 -750 -198 -742
rect -194 -750 -186 -742
rect -206 -755 -198 -750
rect -206 -763 -186 -755
rect -206 -781 -198 -763
rect -194 -776 -186 -768
rect -206 -789 -186 -781
rect -225 -803 -217 -795
rect -206 -807 -198 -789
rect -194 -802 -186 -794
rect -206 -815 -186 -807
rect -194 -828 -186 -820
<< labels >>
rlabel metal1 -190 -745 -190 -745 5 Vdd!
rlabel metal1 -190 -771 -190 -771 5 Vdd!
rlabel metal1 -190 -824 -190 -824 1 Vdd!
rlabel metal1 -190 -733 -190 -733 5 x
rlabel metal1 -190 -695 -190 -695 1 Vdd!
rlabel metal1 -190 -707 -190 -707 5 x
rlabel metal1 -190 -720 -190 -720 1 Vdd!
rlabel metal1 -190 -759 -190 -759 1 x
rlabel metal1 -190 -785 -190 -785 5 x
rlabel metal1 -190 -811 -190 -811 1 x
rlabel metal1 -190 -798 -190 -798 1 Vdd!
rlabel metal1 -190 -669 -190 -669 1 Vdd!
rlabel metal1 -190 -681 -190 -681 5 x
rlabel polysilicon -226 -700 -226 -700 3 f
rlabel polysilicon -226 -753 -226 -753 3 f
rlabel polysilicon -226 -761 -226 -761 3 e
rlabel polysilicon -226 -769 -226 -769 1 d
rlabel polysilicon -226 -793 -226 -793 3 a
rlabel polysilicon -226 -785 -226 -785 3 b
rlabel polysilicon -226 -777 -226 -777 3 c
rlabel metal1 -221 -799 -221 -799 1 GND!
rlabel metal1 -221 -693 -221 -693 5 GND!
rlabel polysilicon -226 -708 -226 -708 3 e
rlabel polysilicon -226 -716 -226 -716 1 d
rlabel metal1 -221 -746 -221 -746 5 x
rlabel polysilicon -226 -724 -226 -724 3 c
rlabel polysilicon -226 -732 -226 -732 3 b
rlabel polysilicon -226 -740 -226 -740 3 a
rlabel polysilicon -185 -818 -185 -818 7 a
rlabel polysilicon -185 -805 -185 -805 7 b
rlabel polysilicon -185 -792 -185 -792 7 b
rlabel polysilicon -185 -779 -185 -779 7 c
rlabel polysilicon -185 -766 -185 -766 7 d
rlabel polysilicon -185 -753 -185 -753 7 f
rlabel polysilicon -185 -740 -185 -740 7 a
rlabel polysilicon -185 -727 -185 -727 7 c
rlabel polysilicon -185 -714 -185 -714 7 d
rlabel polysilicon -185 -701 -185 -701 7 e
rlabel polysilicon -185 -688 -185 -688 7 e
rlabel polysilicon -185 -675 -185 -675 7 f
rlabel space -230 -803 -225 -689 7 ^n
rlabel space -186 -828 -181 -664 3 ^p
<< end >>
