//                                                                             
// File:       mby_regs_ral_env.svh                                            
// Creator:    kmoses1                                                         
// Time:       Sunday Feb 2, 2014 [8:09:00 am]                                 
//                                                                             
// Path:       /tmp/kmoses1/nebulon_run/24391                                  
// Arguments:  /p/com/eda/denali/blueprint/3.7.4/Linux/blueprint -html -I      
//             /p/com/eda/intel/nebulon/2.07p2/include -I source/rdl/ -ovm     
//             mby_ip.rdl                                                      
//                                                                             
// Sources:    /nfs/iil/proj/mpg/kmoses1_wa1/ip_template-nhdk-x0_new/source/rdl/mby_cfg.rdl:02df54a73913bfd13bbaa467d89a076e
//             /nfs/iil/proj/mpg/kmoses1_wa1/ip_template-nhdk-x0_new/source/rdl/mby_mem.rdl:14594b1f2ecfcc36a63682f03cdcd2a5
//             /nfs/iil/proj/mpg/kmoses1_wa1/ip_template-nhdk-x0_new/source/rdl/mby_ip.rdl:7e800c616354c3f9ffd5f5ffffc8f907
//             /p/com/eda/intel/nebulon/2.07p2/generators/generator_common.pm:4973c402c43f97e18c4aba02585df570
//             /p/com/eda/intel/nebulon/2.07p2/generators/html.pm:a408055bdb3ba8a9656d793e9472104f
//             /p/com/eda/intel/nebulon/2.07p2/generators/ovm.pm:e21c7be001887ff41e17c43b43b1fcdc
//             /p/com/eda/intel/nebulon/2.07p2/include/lib_udp.rdl:34d6f45292e06a11e6a71125356fa028
//             /usr/intel/pkgs/perl/5.8.7/lib64/5.8.7/Digest/base.pm:54bebd0439900c1d44d212cba39747b5
//             /usr/intel/pkgs/perl/5.8.7/lib64/site_perl/Devel/StackTrace.pm:3b99e973435e2dea00aa3a8d6f1b9ddd
//                                                                             
// Blueprint:   3.7.4 (Tue Jun 23 00:17:01 PDT 2009)                           
// Machine:    icsl0104                                                        
// OS:         Linux 2.6.16.60-0.58.1.3835.0.PTF.638363-smp                    
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2014 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY DENALI BLUEPRINT, DO NOT EDIT       
//                                                                             


//RAL code compatible with Saola versions: v20131113 and newer 

`ifndef SLA_PATH_TO_STRING
`define SLA_PATH_TO_STRING(SIG_PATH) `"SIG_PATH`"
`endif

`include "mby_regs_regs.svh"


class mby_regs_ral_env extends sla_ral_env;

  `ovm_component_utils(mby_regs_ral_env);

  rand mby_regs_file mby_regs;

  // --------------------------
  function new( string n="mby_regs_ral_env", ovm_component p = null, string hdl_path = "");
    super.new( n, p, hdl_path);
  endfunction : new


  // --------------------------
  virtual function void build();
    super.build();

    mby_regs = mby_regs_file::type_id::create("mby_regs", this);
    add_file("mby_regs",mby_regs);

  endfunction : build

  // --------------------------
  function void connect();
    mby_regs.set_base(4'h0);


    set_bit_blasting(1);
  endfunction : connect


  virtual function string sprint_sv_ral_env();  
     return({"Generated SV RAL Env ---> ", `__FILE__}); 
  endfunction  
endclass : mby_regs_ral_env
