magic
tech scmos
timestamp 982685391
<< nselect >>
rect -33 25 0 88
<< pselect >>
rect 0 17 46 96
<< ndiffusion >>
rect -28 74 -8 75
rect -28 66 -8 71
rect -28 58 -8 63
rect -28 50 -8 55
rect -28 42 -8 47
rect -28 38 -8 39
<< pdiffusion >>
rect 8 84 40 85
rect 8 80 40 81
rect 8 71 40 72
rect 8 67 40 68
rect 28 59 40 67
rect 8 58 40 59
rect 8 54 40 55
rect 8 45 40 46
rect 8 41 40 42
rect 28 33 40 41
rect 8 32 40 33
rect 8 28 40 29
<< ntransistor >>
rect -28 71 -8 74
rect -28 63 -8 66
rect -28 55 -8 58
rect -28 47 -8 50
rect -28 39 -8 42
<< ptransistor >>
rect 8 81 40 84
rect 8 68 40 71
rect 8 55 40 58
rect 8 42 40 45
rect 8 29 40 32
<< polysilicon >>
rect -5 81 8 84
rect 40 81 44 84
rect -5 74 -2 81
rect -32 71 -28 74
rect -8 71 -2 74
rect 3 68 8 71
rect 40 68 44 71
rect 3 66 6 68
rect -32 63 -28 66
rect -8 63 6 66
rect -32 55 -28 58
rect -8 55 8 58
rect 40 55 44 58
rect -32 47 -28 50
rect -8 47 6 50
rect 3 45 6 47
rect 3 42 8 45
rect 40 42 44 45
rect -32 39 -28 42
rect -8 39 -2 42
rect -5 32 -2 39
rect -5 29 8 32
rect 40 29 44 32
<< ndcontact >>
rect -28 75 -8 83
rect -28 30 -8 38
<< pdcontact >>
rect 8 85 40 93
rect 8 72 40 80
rect 8 59 28 67
rect 8 46 40 54
rect 8 33 28 41
rect 8 20 40 28
<< metal1 >>
rect -4 85 40 93
rect -4 83 4 85
rect -28 75 4 83
rect -4 67 4 75
rect 8 79 40 80
rect 8 73 9 79
rect 27 73 40 79
rect 8 72 40 73
rect -4 59 28 67
rect -4 41 4 59
rect 32 54 40 72
rect 8 46 40 54
rect -28 30 -8 38
rect -4 33 28 41
rect -27 25 -9 30
rect 32 28 40 46
rect 8 25 40 28
rect 8 20 9 25
rect 27 20 40 25
<< m2contact >>
rect 9 73 27 79
rect -27 19 -9 25
rect 9 19 27 25
<< m3contact >>
rect 9 73 27 79
rect -27 19 -9 25
rect 9 19 27 25
<< metal3 >>
rect -27 17 -9 96
rect 9 17 27 96
<< labels >>
rlabel space -34 24 -28 89 7 ^n
rlabel space 28 17 47 96 3 ^p
rlabel metal3 -27 17 -9 96 1 GND!|pin|s|0
rlabel metal1 -28 30 -8 38 1 GND!|pin|s|0
rlabel metal1 -27 19 -9 38 1 GND!|pin|s|0
rlabel metal3 9 17 27 96 1 Vdd!|pin|s|1
rlabel metal1 8 72 40 80 1 Vdd!|pin|s|1
rlabel metal1 8 46 40 54 1 Vdd!|pin|s|1
rlabel metal1 8 20 40 28 1 Vdd!|pin|s|1
rlabel metal1 32 20 40 80 1 Vdd!|pin|s|1
rlabel metal1 -4 33 4 93 1 x|pin|s|2
rlabel metal1 -28 75 4 83 1 x|pin|s|2
rlabel metal1 -4 85 40 93 1 x|pin|s|2
rlabel metal1 -4 59 28 67 1 x|pin|s|2
rlabel metal1 -4 33 28 41 1 x|pin|s|2
rlabel polysilicon 40 29 44 32 1 a|pin|w|3|poly
rlabel polysilicon -2 29 2 32 1 a|pin|w|3|poly
rlabel polysilicon -32 39 -28 42 1 a|pin|w|3|poly
rlabel polysilicon 40 42 44 45 1 b|pin|w|4|poly
rlabel polysilicon -32 47 -28 50 1 b|pin|w|4|poly
rlabel polysilicon 40 55 44 58 1 c|pin|w|5|poly
rlabel polysilicon -32 55 -28 58 1 c|pin|w|5|poly
rlabel polysilicon -32 63 -28 66 1 d|pin|w|6|poly
rlabel polysilicon 40 68 44 71 1 d|pin|w|6|poly
rlabel polysilicon 40 81 44 84 1 e|pin|w|7|poly
rlabel polysilicon -2 81 2 84 1 e|pin|w|7|poly
rlabel polysilicon -32 71 -28 74 1 e|pin|w|7|poly
<< end >>
