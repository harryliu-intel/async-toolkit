magic
tech scmos
timestamp 962519129
<< ndiffusion >>
rect 24 108 36 109
rect 24 102 36 106
rect 1 90 9 91
rect 24 96 36 100
rect 24 90 36 94
rect 1 84 9 88
rect 24 84 36 88
rect 1 81 9 82
rect 1 77 5 81
rect 1 76 9 77
rect 24 81 36 82
rect 24 76 36 77
rect 1 70 9 74
rect 24 70 36 74
rect 1 67 9 68
rect 1 63 3 67
rect 1 62 9 63
rect 1 56 9 60
rect 24 64 36 68
rect 24 58 36 62
rect 1 53 9 54
rect 1 49 2 53
rect 24 52 36 56
rect 24 49 36 50
rect 28 43 36 45
rect 28 40 36 41
<< pdiffusion >>
rect 74 118 82 121
rect 74 117 86 118
rect 74 113 86 115
rect 83 109 86 113
rect 56 108 86 109
rect 90 109 92 113
rect 90 108 96 109
rect 56 105 86 106
rect 83 101 86 105
rect 56 100 86 101
rect 90 105 96 106
rect 94 101 96 105
rect 90 100 96 101
rect 56 97 86 98
rect 56 93 63 97
rect 56 92 86 93
rect 90 97 96 98
rect 90 93 92 97
rect 90 92 96 93
rect 56 89 86 90
rect 83 85 86 89
rect 56 84 86 85
rect 90 89 96 90
rect 94 85 96 89
rect 90 84 96 85
rect 56 81 86 82
rect 83 77 86 81
rect 56 76 86 77
rect 90 81 96 82
rect 90 77 92 81
rect 90 76 96 77
rect 56 73 86 74
rect 81 69 86 73
rect 56 68 86 69
rect 90 73 96 74
rect 94 69 96 73
rect 90 68 96 69
rect 56 65 86 66
rect 56 61 63 65
rect 56 60 86 61
rect 90 65 96 66
rect 90 61 92 65
rect 90 60 96 61
rect 56 57 86 58
rect 83 53 86 57
rect 56 52 86 53
rect 90 57 96 58
rect 94 53 96 57
rect 90 52 96 53
rect 56 49 86 50
rect 90 48 96 50
rect 56 43 68 45
rect 90 43 102 44
rect 56 40 68 41
rect 90 40 102 41
<< ntransistor >>
rect 24 106 36 108
rect 24 100 36 102
rect 24 94 36 96
rect 1 88 9 90
rect 24 88 36 90
rect 1 82 9 84
rect 24 82 36 84
rect 1 74 9 76
rect 24 74 36 76
rect 1 68 9 70
rect 24 68 36 70
rect 1 60 9 62
rect 24 62 36 64
rect 24 56 36 58
rect 1 54 9 56
rect 24 50 36 52
rect 28 41 36 43
<< ptransistor >>
rect 74 115 86 117
rect 56 106 86 108
rect 90 106 96 108
rect 56 98 86 100
rect 90 98 96 100
rect 56 90 86 92
rect 90 90 96 92
rect 56 82 86 84
rect 90 82 96 84
rect 56 74 86 76
rect 90 74 96 76
rect 56 66 86 68
rect 90 66 96 68
rect 56 58 86 60
rect 90 58 96 60
rect 56 50 86 52
rect 90 50 96 52
rect 56 41 68 43
rect 90 41 102 43
<< polysilicon >>
rect 71 115 74 117
rect 86 115 89 117
rect 21 106 24 108
rect 36 106 39 108
rect 42 106 56 108
rect 86 106 90 108
rect 96 106 99 108
rect 42 102 44 106
rect 16 100 24 102
rect 36 100 44 102
rect 16 90 18 100
rect 47 98 56 100
rect 86 98 90 100
rect 96 98 99 100
rect 47 96 49 98
rect 21 94 24 96
rect 36 94 49 96
rect 52 90 56 92
rect 86 90 90 92
rect 96 90 99 92
rect -2 88 1 90
rect 9 88 18 90
rect 21 88 24 90
rect 36 88 54 90
rect -2 82 1 84
rect 9 82 24 84
rect 36 82 56 84
rect 86 82 90 84
rect 96 82 99 84
rect -2 74 1 76
rect 9 74 24 76
rect 36 74 56 76
rect 86 74 90 76
rect 96 74 99 76
rect -2 68 1 70
rect 9 68 18 70
rect 21 68 24 70
rect 36 68 54 70
rect -1 60 1 62
rect 9 60 13 62
rect 16 58 18 68
rect 52 66 56 68
rect 86 66 90 68
rect 96 66 99 68
rect 21 62 24 64
rect 36 62 49 64
rect 47 60 49 62
rect 47 58 56 60
rect 86 58 90 60
rect 96 58 99 60
rect 16 56 24 58
rect 36 56 44 58
rect -2 54 1 56
rect 9 54 13 56
rect 11 52 13 54
rect 42 55 44 56
rect 42 53 54 55
rect 52 52 54 53
rect 11 50 24 52
rect 36 50 39 52
rect 52 50 56 52
rect 86 50 90 52
rect 96 50 99 52
rect 25 41 28 43
rect 36 41 56 43
rect 68 41 71 43
rect 77 41 90 43
rect 102 41 105 43
<< ndcontact >>
rect 24 109 36 113
rect 1 91 9 95
rect 5 77 9 81
rect 24 77 36 81
rect 3 63 9 67
rect 2 49 9 53
rect 24 45 36 49
rect 28 36 36 40
<< pdcontact >>
rect 82 118 86 122
rect 56 109 83 113
rect 92 109 96 113
rect 56 101 83 105
rect 90 101 94 105
rect 63 93 86 97
rect 92 93 96 97
rect 56 85 83 89
rect 90 85 94 89
rect 56 77 83 81
rect 92 77 96 81
rect 56 69 81 73
rect 90 69 94 73
rect 63 61 86 65
rect 92 61 96 65
rect 56 53 83 57
rect 90 53 94 57
rect 56 45 86 49
rect 90 44 102 48
rect 56 36 68 40
rect 90 36 102 40
<< polycontact >>
rect -5 60 -1 64
rect 43 43 47 47
rect 75 37 79 41
<< metal1 >>
rect 82 121 86 122
rect 82 118 89 121
rect 24 109 36 113
rect 56 109 83 113
rect 86 105 89 118
rect 92 109 100 113
rect 56 101 83 105
rect 86 101 94 105
rect -1 91 9 95
rect -1 70 2 91
rect 56 89 60 101
rect 86 97 89 101
rect 97 97 100 109
rect 63 93 89 97
rect 92 93 100 97
rect 86 89 89 93
rect 56 85 83 89
rect 86 85 94 89
rect 5 77 47 81
rect 56 77 83 81
rect 43 73 47 77
rect 86 73 89 85
rect 97 81 100 93
rect 92 77 100 81
rect -1 67 6 70
rect 56 69 81 73
rect -5 60 -1 64
rect 3 63 9 67
rect -5 40 -2 60
rect 2 49 19 53
rect 15 45 36 49
rect 43 43 47 68
rect 56 57 60 69
rect 89 69 94 73
rect 86 65 89 68
rect 97 65 100 77
rect 63 61 89 65
rect 92 61 100 65
rect 86 57 89 61
rect 56 53 83 57
rect 86 54 94 57
rect 90 53 94 54
rect 56 45 86 49
rect 97 48 100 61
rect 75 40 79 41
rect -5 37 79 40
rect 82 40 86 45
rect 90 44 102 48
rect 28 36 36 37
rect 56 36 68 37
rect 82 36 102 40
<< m2contact >>
rect 43 68 48 73
rect 84 68 89 73
<< metal2 >>
rect 43 69 89 73
rect 43 68 48 69
rect 84 68 89 69
<< labels >>
rlabel polysilicon 97 91 97 91 7 _a0
rlabel polysilicon 97 99 97 99 7 _a1
rlabel polysilicon 97 83 97 83 7 _b0
rlabel polysilicon 97 107 97 107 7 _b1
rlabel polysilicon 97 51 97 51 1 _a0
rlabel polysilicon 97 75 97 75 1 _a1
rlabel polysilicon 97 59 97 59 1 _b0
rlabel polysilicon 97 67 97 67 1 _b1
rlabel space 74 36 106 122 3 ^p
rlabel polysilicon 69 42 69 42 7 x
rlabel polysilicon 23 107 23 107 1 _SReset!
rlabel polysilicon 27 42 27 42 7 x
rlabel polysilicon 0 55 0 55 3 _SReset!
rlabel space -6 35 28 114 7 ^n
rlabel polysilicon 73 116 73 116 3 _PReset!
rlabel space 70 115 73 118 3 ^p
rlabel pdcontact 71 47 71 47 1 Vdd!
rlabel pdcontact 71 111 71 111 1 Vdd!
rlabel pdcontact 71 79 71 79 1 Vdd!
rlabel pdcontact 93 55 93 55 1 x
rlabel pdcontact 92 71 92 71 1 x
rlabel pdcontact 92 103 92 103 1 x
rlabel pdcontact 92 87 92 87 1 x
rlabel pdcontact 71 95 71 95 1 x
rlabel pdcontact 71 63 71 63 1 x
rlabel pdcontact 95 38 95 38 1 Vdd!
rlabel ndcontact 30 47 30 47 1 GND!
rlabel ndcontact 30 79 30 79 1 x
rlabel ndcontact 30 111 30 111 1 GND!
rlabel ndcontact 7 79 7 79 1 x
rlabel ndcontact 6 51 6 51 1 GND!
rlabel pdcontact 84 120 84 120 1 x
<< end >>
