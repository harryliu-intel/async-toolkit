// -----------------------------------------------------------------------------
// INTEL CONFIDENTIAL
// Copyright(c) 2018, Intel Corporation. All Rights Reserved
// -----------------------------------------------------------------------------
//
// Created By   :  Raghu P Gudla
// Created On   :  09/22/2018
// Description  :  Include all test island connections for each of the block
//------------------------------------------------------------------------------

`include "hvl_fc_conns.svh"
`include "hvl_igr_ti_conns.svh"

/*
 *  ----------------
 *    End of file
 *  ----------------
*/

// <<< VIM SETTINGS
// vim: ts=4 et
// >>>
