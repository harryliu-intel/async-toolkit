.SUBCKT nch_elvt_mac s g d b 
.ENDS

.SUBCKT pch_elvt_mac s g d b 
.ENDS

.SUBCKT ppode_elvt_mac s g b 
.ENDS

.SUBCKT npode_elvt_mac s g b 
.ENDS
