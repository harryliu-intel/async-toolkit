module write_ecc
  (
input  logic [1013-1:0] i_data,

output logic [1013-1:0] o_data
,output logic [11-1:0] o_chk
  );
logic  xor0000;
logic  xor0001;
logic  xor0002;
logic  xor0003;
logic  xor0004;
logic  xor0005;
logic  xor0006;
logic  xor0007;
logic  xor0008;
logic  xor0009;
logic  xor0010;
logic  xor0011;
logic  xor0012;
logic  xor0013;
logic  xor0014;
logic  xor0015;
logic  xor0016;
logic  xor0017;
logic  xor0018;
logic  xor0019;
logic  xor0020;
logic  xor0021;
logic  xor0022;
logic  xor0023;
logic  xor0024;
logic  xor0025;
logic  xor0026;
logic  xor0027;
logic  xor0028;
logic  xor0029;
logic  xor0030;
logic  xor0031;
logic  xor0032;
logic  xor0033;
logic  xor0034;
logic  xor0035;
logic  xor0036;
logic  xor0037;
logic  xor0038;
logic  xor0039;
logic  xor0040;
logic  xor0041;
logic  xor0042;
logic  xor0043;
logic  xor0044;
logic  xor0045;
logic  xor0046;
logic  xor0047;
logic  xor0048;
logic  xor0049;
logic  xor0050;
logic  xor0051;
logic  xor0052;
logic  xor0053;
logic  xor0054;
logic  xor0055;
logic  xor0056;
logic  xor0057;
logic  xor0058;
logic  xor0059;
logic  xor0060;
logic  xor0061;
logic  xor0062;
logic  xor0063;
logic  xor0064;
logic  xor0065;
logic  xor0066;
logic  xor0067;
logic  xor0068;
logic  xor0069;
logic  xor0070;
logic  xor0071;
logic  xor0072;
logic  xor0073;
logic  xor0074;
logic  xor0075;
logic  xor0076;
logic  xor0077;
logic  xor0078;
logic  xor0079;
logic  xor0080;
logic  xor0081;
logic  xor0082;
logic  xor0083;
logic  xor0084;
logic  xor0085;
logic  xor0086;
logic  xor0087;
logic  xor0088;
logic  xor0089;
logic  xor0090;
logic  xor0091;
logic  xor0092;
logic  xor0093;
logic  xor0094;
logic  xor0095;
logic  xor0096;
logic  xor0097;
logic  xor0098;
logic  xor0099;
logic  xor0100;
logic  xor0101;
logic  xor0102;
logic  xor0103;
logic  xor0104;
logic  xor0105;
logic  xor0106;
logic  xor0107;
logic  xor0108;
logic  xor0109;
logic  xor0110;
logic  xor0111;
logic  xor0112;
logic  xor0113;
logic  xor0114;
logic  xor0115;
logic  xor0116;
logic  xor0117;
logic  xor0118;
logic  xor0119;
logic  xor0120;
logic  xor0121;
logic  xor0122;
logic  xor0123;
logic  xor0124;
logic  xor0125;
logic  xor0126;
logic  xor0127;
logic  xor0128;
logic  xor0129;
logic  xor0130;
logic  xor0131;
logic  xor0132;
logic  xor0133;
logic  xor0134;
logic  xor0135;
logic  xor0136;
logic  xor0137;
logic  xor0138;
logic  xor0139;
logic  xor0140;
logic  xor0141;
logic  xor0142;
logic  xor0143;
logic  xor0144;
logic  xor0145;
logic  xor0146;
logic  xor0147;
logic  xor0148;
logic  xor0149;
logic  xor0150;
logic  xor0151;
logic  xor0152;
logic  xor0153;
logic  xor0154;
logic  xor0155;
logic  xor0156;
logic  xor0157;
logic  xor0158;
logic  xor0159;
logic  xor0160;
logic  xor0161;
logic  xor0162;
logic  xor0163;
logic  xor0164;
logic  xor0165;
logic  xor0166;
logic  xor0167;
logic  xor0168;
logic  xor0169;
logic  xor0170;
logic  xor0171;
logic  xor0172;
logic  xor0173;
logic  xor0174;
logic  xor0175;
logic  xor0176;
logic  xor0177;
logic  xor0178;
logic  xor0179;
logic  xor0180;
logic  xor0181;
logic  xor0182;
logic  xor0183;
logic  xor0184;
logic  xor0185;
logic  xor0186;
logic  xor0187;
logic  xor0188;
logic  xor0189;
logic  xor0190;
logic  xor0191;
logic  xor0192;
logic  xor0193;
logic  xor0194;
logic  xor0195;
logic  xor0196;
logic  xor0197;
logic  xor0198;
logic  xor0199;
logic  xor0200;
logic  xor0201;
logic  xor0202;
logic  xor0203;
logic  xor0204;
logic  xor0205;
logic  xor0206;
logic  xor0207;
logic  xor0208;
logic  xor0209;
logic  xor0210;
logic  xor0211;
logic  xor0212;
logic  xor0213;
logic  xor0214;
logic  xor0215;
logic  xor0216;
logic  xor0217;
logic  xor0218;
logic  xor0219;
logic  xor0220;
logic  xor0221;
logic  xor0222;
logic  xor0223;
logic  xor0224;
logic  xor0225;
logic  xor0226;
logic  xor0227;
logic  xor0228;
logic  xor0229;
logic  xor0230;
logic  xor0231;
logic  xor0232;
logic  xor0233;
logic  xor0234;
logic  xor0235;
logic  xor0236;
logic  xor0237;
logic  xor0238;
logic  xor0239;
logic  xor0240;
logic  xor0241;
logic  xor0242;
logic  xor0243;
logic  xor0244;
logic  xor0245;
logic  xor0246;
logic  xor0247;
logic  xor0248;
logic  xor0249;
logic  xor0250;
logic  xor0251;
logic  xor0252;
logic  xor0253;
logic  xor0254;
logic  xor0255;
logic  xor0256;
logic  xor0257;
logic  xor0258;
logic  xor0259;
logic  xor0260;
logic  xor0261;
logic  xor0262;
logic  xor0263;
logic  xor0264;
logic  xor0265;
logic  xor0266;
logic  xor0267;
logic  xor0268;
logic  xor0269;
logic  xor0270;
logic  xor0271;
logic  xor0272;
logic  xor0273;
logic  xor0274;
logic  xor0275;
logic  xor0276;
logic  xor0277;
logic  xor0278;
logic  xor0279;
logic  xor0280;
logic  xor0281;
logic  xor0282;
logic  xor0283;
logic  xor0284;
logic  xor0285;
logic  xor0286;
logic  xor0287;
logic  xor0288;
logic  xor0289;
logic  xor0290;
logic  xor0291;
logic  xor0292;
logic  xor0293;
logic  xor0294;
logic  xor0295;
logic  xor0296;
logic  xor0297;
logic  xor0298;
logic  xor0299;
logic  xor0300;
logic  xor0301;
logic  xor0302;
logic  xor0303;
logic  xor0304;
logic  xor0305;
logic  xor0306;
logic  xor0307;
logic  xor0308;
logic  xor0309;
logic  xor0310;
logic  xor0311;
logic  xor0312;
logic  xor0313;
logic  xor0314;
logic  xor0315;
logic  xor0316;
logic  xor0317;
logic  xor0318;
logic  xor0319;
logic  xor0320;
logic  xor0321;
logic  xor0322;
logic  xor0323;
logic  xor0324;
logic  xor0325;
logic  xor0326;
logic  xor0327;
logic  xor0328;
logic  xor0329;
logic  xor0330;
logic  xor0331;
logic  xor0332;
logic  xor0333;
logic  xor0334;
logic  xor0335;
logic  xor0336;
logic  xor0337;
logic  xor0338;
logic  xor0339;
logic  xor0340;
logic  xor0341;
logic  xor0342;
logic  xor0343;
logic  xor0344;
logic  xor0345;
logic  xor0346;
logic  xor0347;
logic  xor0348;
logic  xor0349;
logic  xor0350;
logic  xor0351;
logic  xor0352;
logic  xor0353;
logic  xor0354;
logic  xor0355;
logic  xor0356;
logic  xor0357;
logic  xor0358;
logic  xor0359;
logic  xor0360;
logic  xor0361;
logic  xor0362;
logic  xor0363;
logic  xor0364;
logic  xor0365;
logic  xor0366;
logic  xor0367;
logic  xor0368;
logic  xor0369;
logic  xor0370;
logic  xor0371;
logic  xor0372;
logic  xor0373;
logic  xor0374;
logic  xor0375;
logic  xor0376;
logic  xor0377;
logic  xor0378;
logic  xor0379;
logic  xor0380;
logic  xor0381;
logic  xor0382;
logic  xor0383;
logic  xor0384;
logic  xor0385;
logic  xor0386;
logic  xor0387;
logic  xor0388;
logic  xor0389;
logic  xor0390;
logic  xor0391;
logic  xor0392;
logic  xor0393;
logic  xor0394;
logic  xor0395;
logic  xor0396;
logic  xor0397;
logic  xor0398;
logic  xor0399;
logic  xor0400;
logic  xor0401;
logic  xor0402;
logic  xor0403;
logic  xor0404;
logic  xor0405;
logic  xor0406;
logic  xor0407;
logic  xor0408;
logic  xor0409;
logic  xor0410;
logic  xor0411;
logic  xor0412;
logic  xor0413;
logic  xor0414;
logic  xor0415;
logic  xor0416;
logic  xor0417;
logic  xor0418;
logic  xor0419;
logic  xor0420;
logic  xor0421;
logic  xor0422;
logic  xor0423;
logic  xor0424;
logic  xor0425;
logic  xor0426;
logic  xor0427;
logic  xor0428;
logic  xor0429;
logic  xor0430;
logic  xor0431;
logic  xor0432;
logic  xor0433;
logic  xor0434;
logic  xor0435;
logic  xor0436;
logic  xor0437;
logic  xor0438;
logic  xor0439;
logic  xor0440;
logic  xor0441;
logic  xor0442;
logic  xor0443;
logic  xor0444;
logic  xor0445;
logic  xor0446;
logic  xor0447;
logic  xor0448;
logic  xor0449;
logic  xor0450;
logic  xor0451;
logic  xor0452;
logic  xor0453;
logic  xor0454;
logic  xor0455;
logic  xor0456;
logic  xor0457;
logic  xor0458;
logic  xor0459;
logic  xor0460;
logic  xor0461;
logic  xor0462;
logic  xor0463;
logic  xor0464;
logic  xor0465;
logic  xor0466;
logic  xor0467;
logic  xor0468;
logic  xor0469;
logic  xor0470;
logic  xor0471;
logic  xor0472;
logic  xor0473;
logic  xor0474;
logic  xor0475;
logic  xor0476;
logic  xor0477;
logic  xor0478;
logic  xor0479;
logic  xor0480;
logic  xor0481;
logic  xor0482;
logic  xor0483;
logic  xor0484;
logic  xor0485;
logic  xor0486;
logic  xor0487;
logic  xor0488;
logic  xor0489;
logic  xor0490;
logic  xor0491;
logic  xor0492;
logic  xor0493;
logic  xor0494;
logic  xor0495;
logic  xor0496;
logic  xor0497;
logic  xor0498;
logic  xor0499;
logic  xor0500;
logic  xor0501;
logic  xor0502;
logic  xor0503;
logic  xor0504;
logic  xor0505;
logic  xor0506;
logic  xor0507;
logic  xor0508;
logic  xor0509;
logic  xor0510;
logic  xor0511;
logic  xor0512;
logic  xor0513;
logic  xor0514;
logic  xor0515;
logic  xor0516;
logic  xor0517;
logic  xor0518;
logic  xor0519;
logic  xor0520;
logic  xor0521;
logic  xor0522;
logic  xor0523;
logic  xor0524;
logic  xor0525;
logic  xor0526;
logic  xor0527;
logic  xor0528;
logic  xor0529;
logic  xor0530;
logic  xor0531;
logic  xor0532;
logic  xor0533;
logic  xor0534;
logic  xor0535;
logic  xor0536;
logic  xor0537;
logic  xor0538;
logic  xor0539;
logic  xor0540;
logic  xor0541;
logic  xor0542;
logic  xor0543;
logic  xor0544;
logic  xor0545;
logic  xor0546;
logic  xor0547;
logic  xor0548;
logic  xor0549;
logic  xor0550;
logic  xor0551;
logic  xor0552;
logic  xor0553;
logic  xor0554;
logic  xor0555;
logic  xor0556;
logic  xor0557;
logic  xor0558;
logic  xor0559;
logic  xor0560;
logic  xor0561;
logic  xor0562;
logic  xor0563;
logic  xor0564;
logic  xor0565;
logic  xor0566;
logic  xor0567;
logic  xor0568;
logic  xor0569;
logic  xor0570;
logic  xor0571;
logic  xor0572;
logic  xor0573;
logic  xor0574;
logic  xor0575;
logic  xor0576;
logic  xor0577;
logic  xor0578;
logic  xor0579;
logic  xor0580;
logic  xor0581;
logic  xor0582;
logic  xor0583;
logic  xor0584;
logic  xor0585;
logic  xor0586;
logic  xor0587;
logic  xor0588;
logic  xor0589;
logic  xor0590;
logic  xor0591;
logic  xor0592;
logic  xor0593;
logic  xor0594;
logic  xor0595;
logic  xor0596;
logic  xor0597;
logic  xor0598;
logic  xor0599;
logic  xor0600;
logic  xor0601;
logic  xor0602;
logic  xor0603;
logic  xor0604;
logic  xor0605;
logic  xor0606;
logic  xor0607;
logic  xor0608;
logic  xor0609;
logic  xor0610;
logic  xor0611;
logic  xor0612;
logic  xor0613;
logic  xor0614;
logic  xor0615;
logic  xor0616;
logic  xor0617;
logic  xor0618;
logic  xor0619;
logic  xor0620;
logic  xor0621;
logic  xor0622;
logic  xor0623;
logic  xor0624;
logic  xor0625;
logic  xor0626;
logic  xor0627;
logic  xor0628;
logic  xor0629;
logic  xor0630;
logic  xor0631;
logic  xor0632;
logic  xor0633;
logic  xor0634;
logic  xor0635;
logic  xor0636;
logic  xor0637;
logic  xor0638;
logic  xor0639;
logic  xor0640;
logic  xor0641;
logic  xor0642;
logic  xor0643;
logic  xor0644;
logic  xor0645;
logic  xor0646;
logic  xor0647;
logic  xor0648;
logic  xor0649;
logic  xor0650;
logic  xor0651;
logic  xor0652;
logic  xor0653;
logic  xor0654;
logic  xor0655;
logic  xor0656;
logic  xor0657;
logic  xor0658;
logic  xor0659;
logic  xor0660;
logic  xor0661;
logic  xor0662;
logic  xor0663;
logic  xor0664;
logic  xor0665;
logic  xor0666;
logic  xor0667;
logic  xor0668;
logic  xor0669;
logic  xor0670;
logic  xor0671;
logic  xor0672;
logic  xor0673;
logic  xor0674;
logic  xor0675;
logic  xor0676;
logic  xor0677;
logic  xor0678;
logic  xor0679;
logic  xor0680;
logic  xor0681;
logic  xor0682;
logic  xor0683;
logic  xor0684;
logic  xor0685;
logic  xor0686;
logic  xor0687;
logic  xor0688;
logic  xor0689;
logic  xor0690;
logic  xor0691;
logic  xor0692;
logic  xor0693;
logic  xor0694;
logic  xor0695;
logic  xor0696;
logic  xor0697;
logic  xor0698;
logic  xor0699;
logic  xor0700;
logic  xor0701;
logic  xor0702;
logic  xor0703;
logic  xor0704;
logic  xor0705;
logic  xor0706;
logic  xor0707;
logic  xor0708;
logic  xor0709;
logic  xor0710;
logic  xor0711;
logic  xor0712;
logic  xor0713;
logic  xor0714;
logic  xor0715;
logic  xor0716;
logic  xor0717;
logic  xor0718;
logic  xor0719;
logic  xor0720;
logic  xor0721;
logic  xor0722;
logic  xor0723;
logic  xor0724;
logic  xor0725;
logic  xor0726;
logic  xor0727;
logic  xor0728;
logic  xor0729;
logic  xor0730;
logic  xor0731;
logic  xor0732;
logic  xor0733;
logic  xor0734;
logic  xor0735;
logic  xor0736;
logic  xor0737;
logic  xor0738;
logic  xor0739;
logic  xor0740;
logic  xor0741;
logic  xor0742;
logic  xor0743;
logic  xor0744;
logic  xor0745;
logic  xor0746;
logic  xor0747;
logic  xor0748;
logic  xor0749;
logic  xor0750;
logic  xor0751;
logic  xor0752;
logic  xor0753;
logic  xor0754;
logic  xor0755;
logic  xor0756;
logic  xor0757;
logic  xor0758;
logic  xor0759;
logic  xor0760;
logic  xor0761;
logic  xor0762;
logic  xor0763;
logic  xor0764;
logic  xor0765;
logic  xor0766;
logic  xor0767;
logic  xor0768;
logic  xor0769;
logic  xor0770;
logic  xor0771;
logic  xor0772;
logic  xor0773;
logic  xor0774;
logic  xor0775;
logic  xor0776;
logic  xor0777;
logic  xor0778;
logic  xor0779;
logic  xor0780;
logic  xor0781;
logic  xor0782;
logic  xor0783;
logic  xor0784;
logic  xor0785;
logic  xor0786;
logic  xor0787;
logic  xor0788;
logic  xor0789;
logic  xor0790;
logic  xor0791;
logic  xor0792;
logic  xor0793;
logic  xor0794;
logic  xor0795;
logic  xor0796;
logic  xor0797;
logic  xor0798;
logic  xor0799;
logic  xor0800;
logic  xor0801;
logic  xor0802;
logic  xor0803;
logic  xor0804;
logic  xor0805;
logic  xor0806;
logic  xor0807;
logic  xor0808;
logic  xor0809;
logic  xor0810;
logic  xor0811;
logic  xor0812;
logic  xor0813;
logic  xor0814;
logic  xor0815;
logic  xor0816;
logic  xor0817;
logic  xor0818;
logic  xor0819;
logic  xor0820;
logic  xor0821;
logic  xor0822;
logic  xor0823;
logic  xor0824;
logic  xor0825;
logic  xor0826;
logic  xor0827;
logic  xor0828;
logic  xor0829;
logic  xor0830;
logic  xor0831;
logic  xor0832;
logic  xor0833;
logic  xor0834;
logic  xor0835;
logic  xor0836;
logic  xor0837;
logic  xor0838;
logic  xor0839;
logic  xor0840;
logic  xor0841;
logic  xor0842;
logic  xor0843;
logic  xor0844;
logic  xor0845;
logic  xor0846;
logic  xor0847;
logic  xor0848;
logic  xor0849;
logic  xor0850;
logic  xor0851;
logic  xor0852;
logic  xor0853;
logic  xor0854;
logic  xor0855;
logic  xor0856;
logic  xor0857;
logic  xor0858;
logic  xor0859;
logic  xor0860;
logic  xor0861;
logic  xor0862;
logic  xor0863;
logic  xor0864;
logic  xor0865;
logic  xor0866;
logic  xor0867;
logic  xor0868;
logic  xor0869;
logic  xor0870;
logic  xor0871;
logic  xor0872;
logic  xor0873;
logic  xor0874;
logic  xor0875;
logic  xor0876;
logic  xor0877;
logic  xor0878;
logic  xor0879;
logic  xor0880;
logic  xor0881;
logic  xor0882;
logic  xor0883;
logic  xor0884;
logic  xor0885;
logic  xor0886;
logic  xor0887;
logic  xor0888;
logic  xor0889;
logic  xor0890;
logic  xor0891;
logic  xor0892;
logic  xor0893;
logic  xor0894;
logic  xor0895;
logic  xor0896;
logic  xor0897;
logic  xor0898;
logic  xor0899;
logic  xor0900;
logic  xor0901;
logic  xor0902;
logic  xor0903;
logic  xor0904;
logic  xor0905;
logic  xor0906;
logic  xor0907;
logic  xor0908;
logic  xor0909;
logic  xor0910;
logic  xor0911;
logic  xor0912;
logic  xor0913;
logic  xor0914;
logic  xor0915;
logic  xor0916;
logic  xor0917;
logic  xor0918;
logic  xor0919;
logic  xor0920;
logic  xor0921;
logic  xor0922;
logic  xor0923;
logic  xor0924;
logic  xor0925;
logic  xor0926;
logic  xor0927;
logic  xor0928;
logic  xor0929;
logic  xor0930;
logic  xor0931;
logic  xor0932;
logic  xor0933;
logic  xor0934;
logic  xor0935;
logic  xor0936;
logic  xor0937;
logic  xor0938;
logic  xor0939;
logic  xor0940;
logic  xor0941;
logic  xor0942;
logic  xor0943;
logic  xor0944;
logic  xor0945;
logic  xor0946;
logic  xor0947;
logic  xor0948;
logic  xor0949;
logic  xor0950;
logic  xor0951;
logic  xor0952;
logic  xor0953;
logic  xor0954;
logic  xor0955;
logic  xor0956;
logic  xor0957;
logic  xor0958;
logic  xor0959;
logic  xor0960;
logic  xor0961;
logic  xor0962;
logic  xor0963;
logic  xor0964;
logic  xor0965;
logic  xor0966;
logic  xor0967;
logic  xor0968;
logic  xor0969;
logic  xor0970;
logic  xor0971;
logic  xor0972;
logic  xor0973;
logic  xor0974;
logic  xor0975;
logic  xor0976;
logic  xor0977;
logic  xor0978;
logic  xor0979;
logic  xor0980;
logic  xor0981;
logic  xor0982;
logic  xor0983;
logic  xor0984;
logic  xor0985;
logic  xor0986;
logic  xor0987;
logic  xor0988;
logic  xor0989;
logic  xor0990;
logic  xor0991;
logic  xor0992;
logic  xor0993;
logic  xor0994;
logic  xor0995;
logic  xor0996;
logic  xor0997;
logic  xor0998;
logic  xor0999;
logic  xor1000;
logic  xor1001;
logic  xor1002;
logic  xor1003;
logic  xor1004;
logic  xor1005;
logic  xor1006;
logic  xor1007;
logic  xor1008;
logic  xor1009;
logic  xor1010;
logic  xor1011;
logic  xor1012;
logic  xor1013;
logic  xor1014;
logic  xor1015;
logic  xor1016;
logic  xor1017;
logic  xor1018;
logic  xor1019;
logic  xor1020;
logic  xor1021;
logic  xor1022;
logic  xor1023;
logic  xor1024;
logic  xor1025;
logic  xor1026;
logic  xor1027;
logic  xor1028;
logic  xor1029;
logic  xor1030;
logic  xor1031;
logic  xor1032;
logic  xor1033;
logic  xor1034;
logic  xor1035;
logic  xor1036;
logic  xor1037;
logic  xor1038;
logic  xor1039;
logic  xor1040;
logic  xor1041;
logic  xor1042;
logic  xor1043;
logic  xor1044;
logic  xor1045;
logic  xor1046;
logic  xor1047;
logic  xor1048;
logic  xor1049;
logic  xor1050;
logic  xor1051;
logic  xor1052;
logic  xor1053;
logic  xor1054;
logic  xor1055;
logic  xor1056;
logic  xor1057;
logic  xor1058;
logic  xor1059;
logic  xor1060;
logic  xor1061;
logic  xor1062;
logic  xor1063;
logic  xor1064;
logic  xor1065;
logic  xor1066;
logic  xor1067;
logic  xor1068;
logic  xor1069;
logic  xor1070;
logic  xor1071;
logic  xor1072;
logic  xor1073;
logic  xor1074;
logic  xor1075;
logic  xor1076;
logic  xor1077;
logic  xor1078;
logic  xor1079;
logic  xor1080;
logic  xor1081;
logic  xor1082;
logic  xor1083;
logic  xor1084;
logic  xor1085;
logic  xor1086;
logic  xor1087;
logic  xor1088;
logic  xor1089;
logic  xor1090;
logic  xor1091;
logic  xor1092;
logic  xor1093;
logic  xor1094;
logic  xor1095;
logic  xor1096;
logic  xor1097;
logic  xor1098;
logic  xor1099;
logic  xor1100;
logic  xor1101;
logic  xor1102;
logic  xor1103;
logic  xor1104;
logic  xor1105;
logic  xor1106;
logic  xor1107;
logic  xor1108;
logic  xor1109;
logic  xor1110;
logic  xor1111;
logic  xor1112;
logic  xor1113;
logic  xor1114;
logic  xor1115;
logic  xor1116;
logic  xor1117;
logic  xor1118;
logic  xor1119;
logic  xor1120;
logic  xor1121;
logic  xor1122;
logic  xor1123;
logic  xor1124;
logic  xor1125;
logic  xor1126;
logic  xor1127;
logic  xor1128;
logic  xor1129;
logic  xor1130;
logic  xor1131;
logic[9:-1] ecc_parity;
logic[1023:0] input_data;
// BuildXorTrees
// BuildXorTrees, FirstLevel, f = -1
assign xor0000 = (input_data[0001]^input_data[0000]^input_data[0003]^input_data[0002]); // EmitInputXorGate
assign xor0001 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); // EmitInputXorGate
assign xor0002 = (input_data[0009]^input_data[0008]^input_data[0011]^input_data[0010]); // EmitInputXorGate
assign xor0003 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); // EmitInputXorGate
assign xor0004 = (input_data[0019]^input_data[0018]^input_data[0017]^input_data[0016]); // EmitInputXorGate
assign xor0005 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); // EmitInputXorGate
assign xor0006 = (input_data[0025]^input_data[0024]^input_data[0027]^input_data[0026]); // EmitInputXorGate
assign xor0007 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); // EmitInputXorGate
assign xor0008 = (input_data[0035]^input_data[0034]^input_data[0033]^input_data[0032]); // EmitInputXorGate
assign xor0009 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); // EmitInputXorGate
assign xor0010 = (input_data[0041]^input_data[0040]^input_data[0043]^input_data[0042]); // EmitInputXorGate
assign xor0011 = (input_data[0046]^input_data[0045]^input_data[0044]^input_data[0047]); // EmitInputXorGate
assign xor0012 = (input_data[0051]^input_data[0050]^input_data[0049]^input_data[0048]); // EmitInputXorGate
assign xor0013 = (input_data[0053]^input_data[0052]^input_data[0055]^input_data[0054]); // EmitInputXorGate
assign xor0014 = (input_data[0059]^input_data[0058]^input_data[0057]^input_data[0056]); // EmitInputXorGate
assign xor0015 = (input_data[0063]^input_data[0062]^input_data[0061]^input_data[0060]); // EmitInputXorGate
assign xor0016 = (input_data[0065]^input_data[0064]^input_data[0067]^input_data[0066]); // EmitInputXorGate
assign xor0017 = (input_data[0069]^input_data[0068]^input_data[0071]^input_data[0070]); // EmitInputXorGate
assign xor0018 = (input_data[0072]^input_data[0075]^input_data[0074]^input_data[0073]); // EmitInputXorGate
assign xor0019 = (input_data[0079]^input_data[0078]^input_data[0077]^input_data[0076]); // EmitInputXorGate
assign xor0020 = (input_data[0081]^input_data[0080]^input_data[0083]^input_data[0082]); // EmitInputXorGate
assign xor0021 = (input_data[0085]^input_data[0084]^input_data[0087]^input_data[0086]); // EmitInputXorGate
assign xor0022 = (input_data[0088]^input_data[0091]^input_data[0090]^input_data[0089]); // EmitInputXorGate
assign xor0023 = (input_data[0095]^input_data[0094]^input_data[0093]^input_data[0092]); // EmitInputXorGate
assign xor0024 = (input_data[0097]^input_data[0096]^input_data[0099]^input_data[0098]); // EmitInputXorGate
assign xor0025 = (input_data[0101]^input_data[0100]^input_data[0103]^input_data[0102]); // EmitInputXorGate
assign xor0026 = (input_data[0105]^input_data[0104]^input_data[0107]^input_data[0106]); // EmitInputXorGate
assign xor0027 = (input_data[0111]^input_data[0110]^input_data[0109]^input_data[0108]); // EmitInputXorGate
assign xor0028 = (input_data[0114]^input_data[0113]^input_data[0112]^input_data[0115]); // EmitInputXorGate
assign xor0029 = (input_data[0117]^input_data[0116]^input_data[0119]^input_data[0118]); // EmitInputXorGate
assign xor0030 = (input_data[0121]^input_data[0120]^input_data[0123]^input_data[0122]); // EmitInputXorGate
assign xor0031 = (input_data[0127]^input_data[0126]^input_data[0125]^input_data[0124]); // EmitInputXorGate
assign xor0032 = (input_data[0131]^input_data[0130]^input_data[0129]^input_data[0128]); // EmitInputXorGate
assign xor0033 = (input_data[0133]^input_data[0132]^input_data[0135]^input_data[0134]); // EmitInputXorGate
assign xor0034 = (input_data[0139]^input_data[0138]^input_data[0137]^input_data[0136]); // EmitInputXorGate
assign xor0035 = (input_data[0141]^input_data[0140]^input_data[0143]^input_data[0142]); // EmitInputXorGate
assign xor0036 = (input_data[0145]^input_data[0144]^input_data[0147]^input_data[0146]); // EmitInputXorGate
assign xor0037 = (input_data[0149]^input_data[0148]^input_data[0151]^input_data[0150]); // EmitInputXorGate
assign xor0038 = (input_data[0155]^input_data[0154]^input_data[0153]^input_data[0152]); // EmitInputXorGate
assign xor0039 = (input_data[0159]^input_data[0158]^input_data[0157]^input_data[0156]); // EmitInputXorGate
assign xor0040 = (input_data[0161]^input_data[0160]^input_data[0163]^input_data[0162]); // EmitInputXorGate
assign xor0041 = (input_data[0165]^input_data[0164]^input_data[0167]^input_data[0166]); // EmitInputXorGate
assign xor0042 = (input_data[0169]^input_data[0168]^input_data[0171]^input_data[0170]); // EmitInputXorGate
assign xor0043 = (input_data[0175]^input_data[0174]^input_data[0173]^input_data[0172]); // EmitInputXorGate
assign xor0044 = (input_data[0177]^input_data[0176]^input_data[0179]^input_data[0178]); // EmitInputXorGate
assign xor0045 = (input_data[0181]^input_data[0180]^input_data[0183]^input_data[0182]); // EmitInputXorGate
assign xor0046 = (input_data[0187]^input_data[0186]^input_data[0185]^input_data[0184]); // EmitInputXorGate
assign xor0047 = (input_data[0191]^input_data[0190]^input_data[0189]^input_data[0188]); // EmitInputXorGate
assign xor0048 = (input_data[0193]^input_data[0192]^input_data[0195]^input_data[0194]); // EmitInputXorGate
assign xor0049 = (input_data[0196]^input_data[0199]^input_data[0198]^input_data[0197]); // EmitInputXorGate
assign xor0050 = (input_data[0201]^input_data[0200]^input_data[0203]^input_data[0202]); // EmitInputXorGate
assign xor0051 = (input_data[0205]^input_data[0204]^input_data[0207]^input_data[0206]); // EmitInputXorGate
assign xor0052 = (input_data[0211]^input_data[0210]^input_data[0209]^input_data[0208]); // EmitInputXorGate
assign xor0053 = (input_data[0215]^input_data[0214]^input_data[0213]^input_data[0212]); // EmitInputXorGate
assign xor0054 = (input_data[0217]^input_data[0216]^input_data[0219]^input_data[0218]); // EmitInputXorGate
assign xor0055 = (input_data[0221]^input_data[0220]^input_data[0223]^input_data[0222]); // EmitInputXorGate
assign xor0056 = (input_data[0224]^input_data[0227]^input_data[0226]^input_data[0225]); // EmitInputXorGate
assign xor0057 = (input_data[0231]^input_data[0230]^input_data[0229]^input_data[0228]); // EmitInputXorGate
assign xor0058 = (input_data[0233]^input_data[0232]^input_data[0235]^input_data[0234]); // EmitInputXorGate
assign xor0059 = (input_data[0236]^input_data[0239]^input_data[0238]^input_data[0237]); // EmitInputXorGate
assign xor0060 = (input_data[0242]^input_data[0241]^input_data[0240]^input_data[0243]); // EmitInputXorGate
assign xor0061 = (input_data[0245]^input_data[0244]^input_data[0247]^input_data[0246]); // EmitInputXorGate
assign xor0062 = (input_data[0249]^input_data[0248]^input_data[0251]^input_data[0250]); // EmitInputXorGate
assign xor0063 = (input_data[0255]^input_data[0254]^input_data[0253]^input_data[0252]); // EmitInputXorGate
assign xor0064 = (input_data[0259]^input_data[0258]^input_data[0257]^input_data[0256]); // EmitInputXorGate
assign xor0065 = (input_data[0261]^input_data[0260]^input_data[0263]^input_data[0262]); // EmitInputXorGate
assign xor0066 = (input_data[0265]^input_data[0264]^input_data[0267]^input_data[0266]); // EmitInputXorGate
assign xor0067 = (input_data[0269]^input_data[0268]^input_data[0271]^input_data[0270]); // EmitInputXorGate
assign xor0068 = (input_data[0275]^input_data[0274]^input_data[0273]^input_data[0272]); // EmitInputXorGate
assign xor0069 = (input_data[0278]^input_data[0277]^input_data[0276]^input_data[0279]); // EmitInputXorGate
assign xor0070 = (input_data[0281]^input_data[0280]^input_data[0283]^input_data[0282]); // EmitInputXorGate
assign xor0071 = (input_data[0284]^input_data[0287]^input_data[0286]^input_data[0285]); // EmitInputXorGate
assign xor0072 = (input_data[0291]^input_data[0290]^input_data[0289]^input_data[0288]); // EmitInputXorGate
assign xor0073 = (input_data[0293]^input_data[0292]^input_data[0295]^input_data[0294]); // EmitInputXorGate
assign xor0074 = (input_data[0296]^input_data[0299]^input_data[0298]^input_data[0297]); // EmitInputXorGate
assign xor0075 = (input_data[0301]^input_data[0300]^input_data[0303]^input_data[0302]); // EmitInputXorGate
assign xor0076 = (input_data[0305]^input_data[0304]^input_data[0307]^input_data[0306]); // EmitInputXorGate
assign xor0077 = (input_data[0310]^input_data[0309]^input_data[0308]^input_data[0311]); // EmitInputXorGate
assign xor0078 = (input_data[0313]^input_data[0312]^input_data[0315]^input_data[0314]); // EmitInputXorGate
assign xor0079 = (input_data[0319]^input_data[0318]^input_data[0317]^input_data[0316]); // EmitInputXorGate
assign xor0080 = (input_data[0322]^input_data[0321]^input_data[0320]^input_data[0323]); // EmitInputXorGate
assign xor0081 = (input_data[0325]^input_data[0324]^input_data[0327]^input_data[0326]); // EmitInputXorGate
assign xor0082 = (input_data[0329]^input_data[0328]^input_data[0331]^input_data[0330]); // EmitInputXorGate
assign xor0083 = (input_data[0335]^input_data[0334]^input_data[0333]^input_data[0332]); // EmitInputXorGate
assign xor0084 = (input_data[0339]^input_data[0338]^input_data[0337]^input_data[0336]); // EmitInputXorGate
assign xor0085 = (input_data[0341]^input_data[0340]^input_data[0343]^input_data[0342]); // EmitInputXorGate
assign xor0086 = (input_data[0345]^input_data[0344]^input_data[0347]^input_data[0346]); // EmitInputXorGate
assign xor0087 = (input_data[0348]^input_data[0351]^input_data[0350]^input_data[0349]); // EmitInputXorGate
assign xor0088 = (input_data[0355]^input_data[0354]^input_data[0353]^input_data[0352]); // EmitInputXorGate
assign xor0089 = (input_data[0357]^input_data[0356]^input_data[0359]^input_data[0358]); // EmitInputXorGate
assign xor0090 = (input_data[0361]^input_data[0360]^input_data[0363]^input_data[0362]); // EmitInputXorGate
assign xor0091 = (input_data[0365]^input_data[0364]^input_data[0367]^input_data[0366]); // EmitInputXorGate
assign xor0092 = (input_data[0371]^input_data[0370]^input_data[0369]^input_data[0368]); // EmitInputXorGate
assign xor0093 = (input_data[0373]^input_data[0372]^input_data[0375]^input_data[0374]); // EmitInputXorGate
assign xor0094 = (input_data[0377]^input_data[0376]^input_data[0379]^input_data[0378]); // EmitInputXorGate
assign xor0095 = (input_data[0383]^input_data[0382]^input_data[0381]^input_data[0380]); // EmitInputXorGate
assign xor0096 = (input_data[0385]^input_data[0384]^input_data[0387]^input_data[0386]); // EmitInputXorGate
assign xor0097 = (input_data[0389]^input_data[0388]^input_data[0391]^input_data[0390]); // EmitInputXorGate
assign xor0098 = (input_data[0395]^input_data[0394]^input_data[0393]^input_data[0392]); // EmitInputXorGate
assign xor0099 = (input_data[0399]^input_data[0398]^input_data[0397]^input_data[0396]); // EmitInputXorGate
assign xor0100 = (input_data[0401]^input_data[0400]^input_data[0403]^input_data[0402]); // EmitInputXorGate
assign xor0101 = (input_data[0405]^input_data[0404]^input_data[0407]^input_data[0406]); // EmitInputXorGate
assign xor0102 = (input_data[0411]^input_data[0410]^input_data[0409]^input_data[0408]); // EmitInputXorGate
assign xor0103 = (input_data[0413]^input_data[0412]^input_data[0415]^input_data[0414]); // EmitInputXorGate
assign xor0104 = (input_data[0417]^input_data[0416]^input_data[0419]^input_data[0418]); // EmitInputXorGate
assign xor0105 = (input_data[0421]^input_data[0420]^input_data[0423]^input_data[0422]); // EmitInputXorGate
assign xor0106 = (input_data[0426]^input_data[0425]^input_data[0424]^input_data[0427]); // EmitInputXorGate
assign xor0107 = (input_data[0430]^input_data[0429]^input_data[0428]^input_data[0431]); // EmitInputXorGate
assign xor0108 = (input_data[0433]^input_data[0432]^input_data[0435]^input_data[0434]); // EmitInputXorGate
assign xor0109 = (input_data[0439]^input_data[0438]^input_data[0437]^input_data[0436]); // EmitInputXorGate
assign xor0110 = (input_data[0441]^input_data[0440]^input_data[0443]^input_data[0442]); // EmitInputXorGate
assign xor0111 = (input_data[0445]^input_data[0444]^input_data[0447]^input_data[0446]); // EmitInputXorGate
assign xor0112 = (input_data[0449]^input_data[0448]^input_data[0451]^input_data[0450]); // EmitInputXorGate
assign xor0113 = (input_data[0455]^input_data[0454]^input_data[0453]^input_data[0452]); // EmitInputXorGate
assign xor0114 = (input_data[0459]^input_data[0458]^input_data[0457]^input_data[0456]); // EmitInputXorGate
assign xor0115 = (input_data[0461]^input_data[0460]^input_data[0463]^input_data[0462]); // EmitInputXorGate
assign xor0116 = (input_data[0465]^input_data[0464]^input_data[0467]^input_data[0466]); // EmitInputXorGate
assign xor0117 = (input_data[0468]^input_data[0471]^input_data[0470]^input_data[0469]); // EmitInputXorGate
assign xor0118 = (input_data[0475]^input_data[0474]^input_data[0473]^input_data[0472]); // EmitInputXorGate
assign xor0119 = (input_data[0477]^input_data[0476]^input_data[0479]^input_data[0478]); // EmitInputXorGate
assign xor0120 = (input_data[0481]^input_data[0480]^input_data[0483]^input_data[0482]); // EmitInputXorGate
assign xor0121 = (input_data[0486]^input_data[0485]^input_data[0484]^input_data[0487]); // EmitInputXorGate
assign xor0122 = (input_data[0491]^input_data[0490]^input_data[0489]^input_data[0488]); // EmitInputXorGate
assign xor0123 = (input_data[0493]^input_data[0492]^input_data[0495]^input_data[0494]); // EmitInputXorGate
assign xor0124 = (input_data[0499]^input_data[0498]^input_data[0497]^input_data[0496]); // EmitInputXorGate
assign xor0125 = (input_data[0500]^input_data[0503]^input_data[0502]^input_data[0501]); // EmitInputXorGate
assign xor0126 = (input_data[0505]^input_data[0504]^input_data[0507]^input_data[0506]); // EmitInputXorGate
assign xor0127 = (input_data[0509]^input_data[0508]^input_data[0511]^input_data[0510]); // EmitInputXorGate
assign xor0128 = (input_data[0512]^input_data[0515]^input_data[0514]^input_data[0513]); // EmitInputXorGate
assign xor0129 = (input_data[0519]^input_data[0518]^input_data[0517]^input_data[0516]); // EmitInputXorGate
assign xor0130 = (input_data[0521]^input_data[0520]^input_data[0523]^input_data[0522]); // EmitInputXorGate
assign xor0131 = (input_data[0525]^input_data[0524]^input_data[0527]^input_data[0526]); // EmitInputXorGate
assign xor0132 = (input_data[0529]^input_data[0528]^input_data[0531]^input_data[0530]); // EmitInputXorGate
assign xor0133 = (input_data[0535]^input_data[0534]^input_data[0533]^input_data[0532]); // EmitInputXorGate
assign xor0134 = (input_data[0539]^input_data[0538]^input_data[0537]^input_data[0536]); // EmitInputXorGate
assign xor0135 = (input_data[0541]^input_data[0540]^input_data[0543]^input_data[0542]); // EmitInputXorGate
assign xor0136 = (input_data[0545]^input_data[0544]^input_data[0547]^input_data[0546]); // EmitInputXorGate
assign xor0137 = (input_data[0551]^input_data[0550]^input_data[0549]^input_data[0548]); // EmitInputXorGate
assign xor0138 = (input_data[0554]^input_data[0553]^input_data[0552]^input_data[0555]); // EmitInputXorGate
assign xor0139 = (input_data[0557]^input_data[0556]^input_data[0559]^input_data[0558]); // EmitInputXorGate
assign xor0140 = (input_data[0561]^input_data[0560]^input_data[0563]^input_data[0562]); // EmitInputXorGate
assign xor0141 = (input_data[0567]^input_data[0566]^input_data[0565]^input_data[0564]); // EmitInputXorGate
assign xor0142 = (input_data[0571]^input_data[0570]^input_data[0569]^input_data[0568]); // EmitInputXorGate
assign xor0143 = (input_data[0573]^input_data[0572]^input_data[0575]^input_data[0574]); // EmitInputXorGate
assign xor0144 = (input_data[0579]^input_data[0578]^input_data[0577]^input_data[0576]); // EmitInputXorGate
assign xor0145 = (input_data[0581]^input_data[0580]^input_data[0583]^input_data[0582]); // EmitInputXorGate
assign xor0146 = (input_data[0585]^input_data[0584]^input_data[0587]^input_data[0586]); // EmitInputXorGate
assign xor0147 = (input_data[0589]^input_data[0588]^input_data[0591]^input_data[0590]); // EmitInputXorGate
assign xor0148 = (input_data[0595]^input_data[0594]^input_data[0593]^input_data[0592]); // EmitInputXorGate
assign xor0149 = (input_data[0599]^input_data[0598]^input_data[0597]^input_data[0596]); // EmitInputXorGate
assign xor0150 = (input_data[0601]^input_data[0600]^input_data[0603]^input_data[0602]); // EmitInputXorGate
assign xor0151 = (input_data[0605]^input_data[0604]^input_data[0607]^input_data[0606]); // EmitInputXorGate
assign xor0152 = (input_data[0609]^input_data[0608]^input_data[0611]^input_data[0610]); // EmitInputXorGate
assign xor0153 = (input_data[0613]^input_data[0612]^input_data[0615]^input_data[0614]); // EmitInputXorGate
assign xor0154 = (input_data[0619]^input_data[0618]^input_data[0617]^input_data[0616]); // EmitInputXorGate
assign xor0155 = (input_data[0621]^input_data[0620]^input_data[0623]^input_data[0622]); // EmitInputXorGate
assign xor0156 = (input_data[0625]^input_data[0624]^input_data[0627]^input_data[0626]); // EmitInputXorGate
assign xor0157 = (input_data[0629]^input_data[0628]^input_data[0631]^input_data[0630]); // EmitInputXorGate
assign xor0158 = (input_data[0635]^input_data[0634]^input_data[0633]^input_data[0632]); // EmitInputXorGate
assign xor0159 = (input_data[0639]^input_data[0638]^input_data[0637]^input_data[0636]); // EmitInputXorGate
assign xor0160 = (input_data[0641]^input_data[0640]^input_data[0643]^input_data[0642]); // EmitInputXorGate
assign xor0161 = (input_data[0645]^input_data[0644]^input_data[0647]^input_data[0646]); // EmitInputXorGate
assign xor0162 = (input_data[0651]^input_data[0650]^input_data[0649]^input_data[0648]); // EmitInputXorGate
assign xor0163 = (input_data[0655]^input_data[0654]^input_data[0653]^input_data[0652]); // EmitInputXorGate
assign xor0164 = (input_data[0657]^input_data[0656]^input_data[0659]^input_data[0658]); // EmitInputXorGate
assign xor0165 = (input_data[0661]^input_data[0660]^input_data[0663]^input_data[0662]); // EmitInputXorGate
assign xor0166 = (input_data[0664]^input_data[0667]^input_data[0666]^input_data[0665]); // EmitInputXorGate
assign xor0167 = (input_data[0671]^input_data[0670]^input_data[0669]^input_data[0668]); // EmitInputXorGate
assign xor0168 = (input_data[0673]^input_data[0672]^input_data[0675]^input_data[0674]); // EmitInputXorGate
assign xor0169 = (input_data[0676]^input_data[0679]^input_data[0678]^input_data[0677]); // EmitInputXorGate
assign xor0170 = (input_data[0682]^input_data[0681]^input_data[0680]^input_data[0683]); // EmitInputXorGate
assign xor0171 = (input_data[0685]^input_data[0684]^input_data[0687]^input_data[0686]); // EmitInputXorGate
assign xor0172 = (input_data[0689]^input_data[0688]^input_data[0691]^input_data[0690]); // EmitInputXorGate
assign xor0173 = (input_data[0695]^input_data[0694]^input_data[0693]^input_data[0692]); // EmitInputXorGate
assign xor0174 = (input_data[0699]^input_data[0698]^input_data[0697]^input_data[0696]); // EmitInputXorGate
assign xor0175 = (input_data[0701]^input_data[0700]^input_data[0703]^input_data[0702]); // EmitInputXorGate
assign xor0176 = (input_data[0705]^input_data[0704]^input_data[0707]^input_data[0706]); // EmitInputXorGate
assign xor0177 = (input_data[0709]^input_data[0708]^input_data[0711]^input_data[0710]); // EmitInputXorGate
assign xor0178 = (input_data[0715]^input_data[0714]^input_data[0713]^input_data[0712]); // EmitInputXorGate
assign xor0179 = (input_data[0719]^input_data[0718]^input_data[0717]^input_data[0716]); // EmitInputXorGate
assign xor0180 = (input_data[0721]^input_data[0720]^input_data[0723]^input_data[0722]); // EmitInputXorGate
assign xor0181 = (input_data[0725]^input_data[0724]^input_data[0727]^input_data[0726]); // EmitInputXorGate
assign xor0182 = (input_data[0731]^input_data[0730]^input_data[0729]^input_data[0728]); // EmitInputXorGate
assign xor0183 = (input_data[0735]^input_data[0734]^input_data[0733]^input_data[0732]); // EmitInputXorGate
assign xor0184 = (input_data[0737]^input_data[0736]^input_data[0739]^input_data[0738]); // EmitInputXorGate
assign xor0185 = (input_data[0741]^input_data[0740]^input_data[0743]^input_data[0742]); // EmitInputXorGate
assign xor0186 = (input_data[0745]^input_data[0744]^input_data[0747]^input_data[0746]); // EmitInputXorGate
assign xor0187 = (input_data[0750]^input_data[0749]^input_data[0748]^input_data[0751]); // EmitInputXorGate
assign xor0188 = (input_data[0753]^input_data[0752]^input_data[0755]^input_data[0754]); // EmitInputXorGate
assign xor0189 = (input_data[0759]^input_data[0758]^input_data[0757]^input_data[0756]); // EmitInputXorGate
assign xor0190 = (input_data[0762]^input_data[0761]^input_data[0760]^input_data[0763]); // EmitInputXorGate
assign xor0191 = (input_data[0765]^input_data[0764]^input_data[0767]^input_data[0766]); // EmitInputXorGate
assign xor0192 = (input_data[0769]^input_data[0768]^input_data[0771]^input_data[0770]); // EmitInputXorGate
assign xor0193 = (input_data[0775]^input_data[0774]^input_data[0773]^input_data[0772]); // EmitInputXorGate
assign xor0194 = (input_data[0779]^input_data[0778]^input_data[0777]^input_data[0776]); // EmitInputXorGate
assign xor0195 = (input_data[0781]^input_data[0780]^input_data[0783]^input_data[0782]); // EmitInputXorGate
assign xor0196 = (input_data[0785]^input_data[0784]^input_data[0787]^input_data[0786]); // EmitInputXorGate
assign xor0197 = (input_data[0788]^input_data[0791]^input_data[0790]^input_data[0789]); // EmitInputXorGate
assign xor0198 = (input_data[0795]^input_data[0794]^input_data[0793]^input_data[0792]); // EmitInputXorGate
assign xor0199 = (input_data[0797]^input_data[0796]^input_data[0799]^input_data[0798]); // EmitInputXorGate
assign xor0200 = (input_data[0803]^input_data[0802]^input_data[0801]^input_data[0800]); // EmitInputXorGate
assign xor0201 = (input_data[0805]^input_data[0804]^input_data[0807]^input_data[0806]); // EmitInputXorGate
assign xor0202 = (input_data[0809]^input_data[0808]^input_data[0811]^input_data[0810]); // EmitInputXorGate
assign xor0203 = (input_data[0815]^input_data[0814]^input_data[0813]^input_data[0812]); // EmitInputXorGate
assign xor0204 = (input_data[0819]^input_data[0818]^input_data[0817]^input_data[0816]); // EmitInputXorGate
assign xor0205 = (input_data[0821]^input_data[0820]^input_data[0823]^input_data[0822]); // EmitInputXorGate
assign xor0206 = (input_data[0825]^input_data[0824]^input_data[0827]^input_data[0826]); // EmitInputXorGate
assign xor0207 = (input_data[0829]^input_data[0828]^input_data[0831]^input_data[0830]); // EmitInputXorGate
assign xor0208 = (input_data[0835]^input_data[0834]^input_data[0833]^input_data[0832]); // EmitInputXorGate
assign xor0209 = (input_data[0839]^input_data[0838]^input_data[0837]^input_data[0836]); // EmitInputXorGate
assign xor0210 = (input_data[0841]^input_data[0840]^input_data[0843]^input_data[0842]); // EmitInputXorGate
assign xor0211 = (input_data[0845]^input_data[0844]^input_data[0847]^input_data[0846]); // EmitInputXorGate
assign xor0212 = (input_data[0851]^input_data[0850]^input_data[0849]^input_data[0848]); // EmitInputXorGate
assign xor0213 = (input_data[0853]^input_data[0852]^input_data[0855]^input_data[0854]); // EmitInputXorGate
assign xor0214 = (input_data[0857]^input_data[0856]^input_data[0859]^input_data[0858]); // EmitInputXorGate
assign xor0215 = (input_data[0861]^input_data[0860]^input_data[0863]^input_data[0862]); // EmitInputXorGate
assign xor0216 = (input_data[0866]^input_data[0865]^input_data[0864]^input_data[0867]); // EmitInputXorGate
assign xor0217 = (input_data[0870]^input_data[0869]^input_data[0868]^input_data[0871]); // EmitInputXorGate
assign xor0218 = (input_data[0873]^input_data[0872]^input_data[0875]^input_data[0874]); // EmitInputXorGate
assign xor0219 = (input_data[0879]^input_data[0878]^input_data[0877]^input_data[0876]); // EmitInputXorGate
assign xor0220 = (input_data[0881]^input_data[0880]^input_data[0883]^input_data[0882]); // EmitInputXorGate
assign xor0221 = (input_data[0885]^input_data[0884]^input_data[0887]^input_data[0886]); // EmitInputXorGate
assign xor0222 = (input_data[0889]^input_data[0888]^input_data[0891]^input_data[0890]); // EmitInputXorGate
assign xor0223 = (input_data[0895]^input_data[0894]^input_data[0893]^input_data[0892]); // EmitInputXorGate
assign xor0224 = (input_data[0899]^input_data[0898]^input_data[0897]^input_data[0896]); // EmitInputXorGate
assign xor0225 = (input_data[0901]^input_data[0900]^input_data[0903]^input_data[0902]); // EmitInputXorGate
assign xor0226 = (input_data[0905]^input_data[0904]^input_data[0907]^input_data[0906]); // EmitInputXorGate
assign xor0227 = (input_data[0908]^input_data[0911]^input_data[0910]^input_data[0909]); // EmitInputXorGate
assign xor0228 = (input_data[0915]^input_data[0914]^input_data[0913]^input_data[0912]); // EmitInputXorGate
assign xor0229 = (input_data[0917]^input_data[0916]^input_data[0919]^input_data[0918]); // EmitInputXorGate
assign xor0230 = (input_data[0921]^input_data[0920]^input_data[0923]^input_data[0922]); // EmitInputXorGate
assign xor0231 = (input_data[0925]^input_data[0924]^input_data[0927]^input_data[0926]); // EmitInputXorGate
assign xor0232 = (input_data[0931]^input_data[0930]^input_data[0929]^input_data[0928]); // EmitInputXorGate
assign xor0233 = (input_data[0934]^input_data[0933]^input_data[0932]^input_data[0935]); // EmitInputXorGate
assign xor0234 = (input_data[0937]^input_data[0936]^input_data[0939]^input_data[0938]); // EmitInputXorGate
assign xor0235 = (input_data[0943]^input_data[0942]^input_data[0941]^input_data[0940]); // EmitInputXorGate
assign xor0236 = (input_data[0945]^input_data[0944]^input_data[0947]^input_data[0946]); // EmitInputXorGate
assign xor0237 = (input_data[0949]^input_data[0948]^input_data[0951]^input_data[0950]); // EmitInputXorGate
assign xor0238 = (input_data[0952]^input_data[0955]^input_data[0954]^input_data[0953]); // EmitInputXorGate
assign xor0239 = (input_data[0959]^input_data[0958]^input_data[0957]^input_data[0956]); // EmitInputXorGate
assign xor0240 = (input_data[0961]^input_data[0960]^input_data[0963]^input_data[0962]); // EmitInputXorGate
assign xor0241 = (input_data[0965]^input_data[0964]^input_data[0967]^input_data[0966]); // EmitInputXorGate
assign xor0242 = (input_data[0969]^input_data[0968]^input_data[0971]^input_data[0970]); // EmitInputXorGate
assign xor0243 = (input_data[0975]^input_data[0974]^input_data[0973]^input_data[0972]); // EmitInputXorGate
assign xor0244 = (input_data[0979]^input_data[0978]^input_data[0977]^input_data[0976]); // EmitInputXorGate
assign xor0245 = (input_data[0981]^input_data[0980]^input_data[0983]^input_data[0982]); // EmitInputXorGate
assign xor0246 = (input_data[0985]^input_data[0984]^input_data[0987]^input_data[0986]); // EmitInputXorGate
assign xor0247 = (input_data[0991]^input_data[0990]^input_data[0989]^input_data[0988]); // EmitInputXorGate
assign xor0248 = (input_data[0994]^input_data[0993]^input_data[0992]^input_data[0995]); // EmitInputXorGate
assign xor0249 = (input_data[0997]^input_data[0996]^input_data[0999]^input_data[0998]); // EmitInputXorGate
assign xor0250 = (input_data[1001]^input_data[1000]^input_data[1003]^input_data[1002]); // EmitInputXorGate
assign xor0251 = (input_data[1005]^input_data[1004]^input_data[1007]^input_data[1006]); // EmitInputXorGate
assign xor0252 = (input_data[1008]^input_data[1011]^input_data[1010]^input_data[1009]); // EmitInputXorGate
assign xor0253 = (input_data[1015]^input_data[1014]^input_data[1013]^input_data[1012]); // EmitInputXorGate
assign xor0254 = (input_data[1017]^input_data[1016]^input_data[1019]^input_data[1018]); // EmitInputXorGate
assign xor0255 = (input_data[1021]^input_data[1020]^input_data[1023]^input_data[1022]); // EmitInputXorGate
// BuildXorTrees, FirstLevel, f = 0
assign xor0256 = (input_data[0005]^input_data[0007]^input_data[0001]^input_data[0003]); // EmitInputXorGate
assign xor0257 = (input_data[0009]^input_data[0015]^input_data[0011]^input_data[0013]); // EmitInputXorGate
assign xor0258 = (input_data[0019]^input_data[0017]^input_data[0021]^input_data[0023]); // EmitInputXorGate
assign xor0259 = (input_data[0025]^input_data[0027]^input_data[0031]^input_data[0029]); // EmitInputXorGate
assign xor0260 = (input_data[0035]^input_data[0037]^input_data[0033]^input_data[0039]); // EmitInputXorGate
assign xor0261 = (input_data[0041]^input_data[0043]^input_data[0045]^input_data[0047]); // EmitInputXorGate
assign xor0262 = (input_data[0051]^input_data[0053]^input_data[0049]^input_data[0055]); // EmitInputXorGate
assign xor0263 = (input_data[0063]^input_data[0059]^input_data[0061]^input_data[0057]); // EmitInputXorGate
assign xor0264 = (input_data[0069]^input_data[0065]^input_data[0071]^input_data[0067]); // EmitInputXorGate
assign xor0265 = (input_data[0079]^input_data[0075]^input_data[0077]^input_data[0073]); // EmitInputXorGate
assign xor0266 = (input_data[0085]^input_data[0087]^input_data[0081]^input_data[0083]); // EmitInputXorGate
assign xor0267 = (input_data[0095]^input_data[0091]^input_data[0093]^input_data[0089]); // EmitInputXorGate
assign xor0268 = (input_data[0097]^input_data[0101]^input_data[0103]^input_data[0099]); // EmitInputXorGate
assign xor0269 = (input_data[0105]^input_data[0107]^input_data[0111]^input_data[0109]); // EmitInputXorGate
assign xor0270 = (input_data[0117]^input_data[0113]^input_data[0119]^input_data[0115]); // EmitInputXorGate
assign xor0271 = (input_data[0127]^input_data[0121]^input_data[0123]^input_data[0125]); // EmitInputXorGate
assign xor0272 = (input_data[0131]^input_data[0133]^input_data[0129]^input_data[0135]); // EmitInputXorGate
assign xor0273 = (input_data[0139]^input_data[0141]^input_data[0137]^input_data[0143]); // EmitInputXorGate
assign xor0274 = (input_data[0149]^input_data[0145]^input_data[0147]^input_data[0151]); // EmitInputXorGate
assign xor0275 = (input_data[0159]^input_data[0155]^input_data[0157]^input_data[0153]); // EmitInputXorGate
assign xor0276 = (input_data[0165]^input_data[0167]^input_data[0161]^input_data[0163]); // EmitInputXorGate
assign xor0277 = (input_data[0169]^input_data[0175]^input_data[0171]^input_data[0173]); // EmitInputXorGate
assign xor0278 = (input_data[0181]^input_data[0183]^input_data[0177]^input_data[0179]); // EmitInputXorGate
assign xor0279 = (input_data[0187]^input_data[0191]^input_data[0189]^input_data[0185]); // EmitInputXorGate
assign xor0280 = (input_data[0193]^input_data[0199]^input_data[0195]^input_data[0197]); // EmitInputXorGate
assign xor0281 = (input_data[0205]^input_data[0207]^input_data[0201]^input_data[0203]); // EmitInputXorGate
assign xor0282 = (input_data[0215]^input_data[0211]^input_data[0213]^input_data[0209]); // EmitInputXorGate
assign xor0283 = (input_data[0217]^input_data[0221]^input_data[0223]^input_data[0219]); // EmitInputXorGate
assign xor0284 = (input_data[0231]^input_data[0227]^input_data[0229]^input_data[0225]); // EmitInputXorGate
assign xor0285 = (input_data[0233]^input_data[0239]^input_data[0235]^input_data[0237]); // EmitInputXorGate
assign xor0286 = (input_data[0245]^input_data[0247]^input_data[0241]^input_data[0243]); // EmitInputXorGate
assign xor0287 = (input_data[0249]^input_data[0255]^input_data[0251]^input_data[0253]); // EmitInputXorGate
assign xor0288 = (input_data[0259]^input_data[0257]^input_data[0261]^input_data[0263]); // EmitInputXorGate
assign xor0289 = (input_data[0269]^input_data[0265]^input_data[0267]^input_data[0271]); // EmitInputXorGate
assign xor0290 = (input_data[0275]^input_data[0277]^input_data[0273]^input_data[0279]); // EmitInputXorGate
assign xor0291 = (input_data[0287]^input_data[0281]^input_data[0283]^input_data[0285]); // EmitInputXorGate
assign xor0292 = (input_data[0291]^input_data[0293]^input_data[0289]^input_data[0295]); // EmitInputXorGate
assign xor0293 = (input_data[0301]^input_data[0303]^input_data[0299]^input_data[0297]); // EmitInputXorGate
assign xor0294 = (input_data[0309]^input_data[0305]^input_data[0307]^input_data[0311]); // EmitInputXorGate
assign xor0295 = (input_data[0313]^input_data[0319]^input_data[0315]^input_data[0317]); // EmitInputXorGate
assign xor0296 = (input_data[0325]^input_data[0327]^input_data[0321]^input_data[0323]); // EmitInputXorGate
assign xor0297 = (input_data[0329]^input_data[0335]^input_data[0331]^input_data[0333]); // EmitInputXorGate
assign xor0298 = (input_data[0339]^input_data[0341]^input_data[0343]^input_data[0337]); // EmitInputXorGate
assign xor0299 = (input_data[0345]^input_data[0351]^input_data[0347]^input_data[0349]); // EmitInputXorGate
assign xor0300 = (input_data[0355]^input_data[0357]^input_data[0353]^input_data[0359]); // EmitInputXorGate
assign xor0301 = (input_data[0365]^input_data[0367]^input_data[0361]^input_data[0363]); // EmitInputXorGate
assign xor0302 = (input_data[0371]^input_data[0373]^input_data[0369]^input_data[0375]); // EmitInputXorGate
assign xor0303 = (input_data[0377]^input_data[0383]^input_data[0379]^input_data[0381]); // EmitInputXorGate
assign xor0304 = (input_data[0389]^input_data[0385]^input_data[0387]^input_data[0391]); // EmitInputXorGate
assign xor0305 = (input_data[0399]^input_data[0395]^input_data[0397]^input_data[0393]); // EmitInputXorGate
assign xor0306 = (input_data[0405]^input_data[0407]^input_data[0401]^input_data[0403]); // EmitInputXorGate
assign xor0307 = (input_data[0411]^input_data[0413]^input_data[0409]^input_data[0415]); // EmitInputXorGate
assign xor0308 = (input_data[0417]^input_data[0421]^input_data[0423]^input_data[0419]); // EmitInputXorGate
assign xor0309 = (input_data[0429]^input_data[0425]^input_data[0427]^input_data[0431]); // EmitInputXorGate
assign xor0310 = (input_data[0433]^input_data[0439]^input_data[0435]^input_data[0437]); // EmitInputXorGate
assign xor0311 = (input_data[0445]^input_data[0447]^input_data[0441]^input_data[0443]); // EmitInputXorGate
assign xor0312 = (input_data[0449]^input_data[0455]^input_data[0451]^input_data[0453]); // EmitInputXorGate
assign xor0313 = (input_data[0459]^input_data[0461]^input_data[0457]^input_data[0463]); // EmitInputXorGate
assign xor0314 = (input_data[0465]^input_data[0467]^input_data[0471]^input_data[0469]); // EmitInputXorGate
assign xor0315 = (input_data[0475]^input_data[0477]^input_data[0473]^input_data[0479]); // EmitInputXorGate
assign xor0316 = (input_data[0481]^input_data[0483]^input_data[0485]^input_data[0487]); // EmitInputXorGate
assign xor0317 = (input_data[0491]^input_data[0493]^input_data[0489]^input_data[0495]); // EmitInputXorGate
assign xor0318 = (input_data[0503]^input_data[0499]^input_data[0497]^input_data[0501]); // EmitInputXorGate
assign xor0319 = (input_data[0509]^input_data[0505]^input_data[0507]^input_data[0511]); // EmitInputXorGate
assign xor0320 = (input_data[0519]^input_data[0515]^input_data[0517]^input_data[0513]); // EmitInputXorGate
assign xor0321 = (input_data[0525]^input_data[0527]^input_data[0521]^input_data[0523]); // EmitInputXorGate
assign xor0322 = (input_data[0529]^input_data[0535]^input_data[0531]^input_data[0533]); // EmitInputXorGate
assign xor0323 = (input_data[0539]^input_data[0541]^input_data[0543]^input_data[0537]); // EmitInputXorGate
assign xor0324 = (input_data[0545]^input_data[0551]^input_data[0547]^input_data[0549]); // EmitInputXorGate
assign xor0325 = (input_data[0557]^input_data[0553]^input_data[0559]^input_data[0555]); // EmitInputXorGate
assign xor0326 = (input_data[0567]^input_data[0561]^input_data[0563]^input_data[0565]); // EmitInputXorGate
assign xor0327 = (input_data[0571]^input_data[0573]^input_data[0569]^input_data[0575]); // EmitInputXorGate
assign xor0328 = (input_data[0579]^input_data[0581]^input_data[0577]^input_data[0583]); // EmitInputXorGate
assign xor0329 = (input_data[0589]^input_data[0585]^input_data[0587]^input_data[0591]); // EmitInputXorGate
assign xor0330 = (input_data[0599]^input_data[0595]^input_data[0597]^input_data[0593]); // EmitInputXorGate
assign xor0331 = (input_data[0601]^input_data[0603]^input_data[0605]^input_data[0607]); // EmitInputXorGate
assign xor0332 = (input_data[0613]^input_data[0609]^input_data[0615]^input_data[0611]); // EmitInputXorGate
assign xor0333 = (input_data[0619]^input_data[0621]^input_data[0617]^input_data[0623]); // EmitInputXorGate
assign xor0334 = (input_data[0629]^input_data[0625]^input_data[0627]^input_data[0631]); // EmitInputXorGate
assign xor0335 = (input_data[0639]^input_data[0635]^input_data[0637]^input_data[0633]); // EmitInputXorGate
assign xor0336 = (input_data[0645]^input_data[0647]^input_data[0641]^input_data[0643]); // EmitInputXorGate
assign xor0337 = (input_data[0655]^input_data[0651]^input_data[0653]^input_data[0649]); // EmitInputXorGate
assign xor0338 = (input_data[0657]^input_data[0661]^input_data[0663]^input_data[0659]); // EmitInputXorGate
assign xor0339 = (input_data[0671]^input_data[0667]^input_data[0669]^input_data[0665]); // EmitInputXorGate
assign xor0340 = (input_data[0673]^input_data[0679]^input_data[0675]^input_data[0677]); // EmitInputXorGate
assign xor0341 = (input_data[0685]^input_data[0687]^input_data[0681]^input_data[0683]); // EmitInputXorGate
assign xor0342 = (input_data[0689]^input_data[0695]^input_data[0691]^input_data[0693]); // EmitInputXorGate
assign xor0343 = (input_data[0699]^input_data[0697]^input_data[0701]^input_data[0703]); // EmitInputXorGate
assign xor0344 = (input_data[0709]^input_data[0705]^input_data[0707]^input_data[0711]); // EmitInputXorGate
assign xor0345 = (input_data[0719]^input_data[0715]^input_data[0717]^input_data[0713]); // EmitInputXorGate
assign xor0346 = (input_data[0725]^input_data[0727]^input_data[0721]^input_data[0723]); // EmitInputXorGate
assign xor0347 = (input_data[0735]^input_data[0731]^input_data[0733]^input_data[0729]); // EmitInputXorGate
assign xor0348 = (input_data[0741]^input_data[0743]^input_data[0737]^input_data[0739]); // EmitInputXorGate
assign xor0349 = (input_data[0749]^input_data[0745]^input_data[0747]^input_data[0751]); // EmitInputXorGate
assign xor0350 = (input_data[0753]^input_data[0759]^input_data[0755]^input_data[0757]); // EmitInputXorGate
assign xor0351 = (input_data[0765]^input_data[0767]^input_data[0761]^input_data[0763]); // EmitInputXorGate
assign xor0352 = (input_data[0769]^input_data[0775]^input_data[0771]^input_data[0773]); // EmitInputXorGate
assign xor0353 = (input_data[0779]^input_data[0781]^input_data[0783]^input_data[0777]); // EmitInputXorGate
assign xor0354 = (input_data[0785]^input_data[0791]^input_data[0787]^input_data[0789]); // EmitInputXorGate
assign xor0355 = (input_data[0795]^input_data[0797]^input_data[0793]^input_data[0799]); // EmitInputXorGate
assign xor0356 = (input_data[0803]^input_data[0805]^input_data[0807]^input_data[0801]); // EmitInputXorGate
assign xor0357 = (input_data[0809]^input_data[0815]^input_data[0811]^input_data[0813]); // EmitInputXorGate
assign xor0358 = (input_data[0819]^input_data[0817]^input_data[0821]^input_data[0823]); // EmitInputXorGate
assign xor0359 = (input_data[0829]^input_data[0825]^input_data[0827]^input_data[0831]); // EmitInputXorGate
assign xor0360 = (input_data[0839]^input_data[0835]^input_data[0837]^input_data[0833]); // EmitInputXorGate
assign xor0361 = (input_data[0845]^input_data[0847]^input_data[0841]^input_data[0843]); // EmitInputXorGate
assign xor0362 = (input_data[0851]^input_data[0853]^input_data[0849]^input_data[0855]); // EmitInputXorGate
assign xor0363 = (input_data[0857]^input_data[0861]^input_data[0863]^input_data[0859]); // EmitInputXorGate
assign xor0364 = (input_data[0869]^input_data[0865]^input_data[0867]^input_data[0871]); // EmitInputXorGate
assign xor0365 = (input_data[0873]^input_data[0879]^input_data[0875]^input_data[0877]); // EmitInputXorGate
assign xor0366 = (input_data[0885]^input_data[0887]^input_data[0881]^input_data[0883]); // EmitInputXorGate
assign xor0367 = (input_data[0889]^input_data[0895]^input_data[0891]^input_data[0893]); // EmitInputXorGate
assign xor0368 = (input_data[0899]^input_data[0897]^input_data[0901]^input_data[0903]); // EmitInputXorGate
assign xor0369 = (input_data[0905]^input_data[0907]^input_data[0911]^input_data[0909]); // EmitInputXorGate
assign xor0370 = (input_data[0915]^input_data[0917]^input_data[0913]^input_data[0919]); // EmitInputXorGate
assign xor0371 = (input_data[0925]^input_data[0927]^input_data[0921]^input_data[0923]); // EmitInputXorGate
assign xor0372 = (input_data[0931]^input_data[0933]^input_data[0929]^input_data[0935]); // EmitInputXorGate
assign xor0373 = (input_data[0943]^input_data[0937]^input_data[0939]^input_data[0941]); // EmitInputXorGate
assign xor0374 = (input_data[0949]^input_data[0945]^input_data[0947]^input_data[0951]); // EmitInputXorGate
assign xor0375 = (input_data[0959]^input_data[0955]^input_data[0957]^input_data[0953]); // EmitInputXorGate
assign xor0376 = (input_data[0965]^input_data[0967]^input_data[0961]^input_data[0963]); // EmitInputXorGate
assign xor0377 = (input_data[0969]^input_data[0975]^input_data[0971]^input_data[0973]); // EmitInputXorGate
assign xor0378 = (input_data[0979]^input_data[0981]^input_data[0977]^input_data[0983]); // EmitInputXorGate
assign xor0379 = (input_data[0985]^input_data[0987]^input_data[0991]^input_data[0989]); // EmitInputXorGate
assign xor0380 = (input_data[0997]^input_data[0993]^input_data[0999]^input_data[0995]); // EmitInputXorGate
assign xor0381 = (input_data[1005]^input_data[1007]^input_data[1001]^input_data[1003]); // EmitInputXorGate
assign xor0382 = (input_data[1015]^input_data[1011]^input_data[1013]^input_data[1009]); // EmitInputXorGate
assign xor0383 = (input_data[1017]^input_data[1021]^input_data[1023]^input_data[1019]); // EmitInputXorGate
// BuildXorTrees, FirstLevel, f = 1
assign xor0384 = (input_data[0007]^input_data[0006]^input_data[0003]^input_data[0002]); // EmitInputXorGate
assign xor0385 = (input_data[0015]^input_data[0014]^input_data[0011]^input_data[0010]); // EmitInputXorGate
assign xor0386 = (input_data[0019]^input_data[0018]^input_data[0023]^input_data[0022]); // EmitInputXorGate
assign xor0387 = (input_data[0027]^input_data[0031]^input_data[0030]^input_data[0026]); // EmitInputXorGate
assign xor0388 = (input_data[0035]^input_data[0034]^input_data[0039]^input_data[0038]); // EmitInputXorGate
assign xor0389 = (input_data[0046]^input_data[0043]^input_data[0042]^input_data[0047]); // EmitInputXorGate
assign xor0390 = (input_data[0051]^input_data[0050]^input_data[0055]^input_data[0054]); // EmitInputXorGate
assign xor0391 = (input_data[0063]^input_data[0062]^input_data[0059]^input_data[0058]); // EmitInputXorGate
assign xor0392 = (input_data[0071]^input_data[0067]^input_data[0066]^input_data[0070]); // EmitInputXorGate
assign xor0393 = (input_data[0079]^input_data[0078]^input_data[0075]^input_data[0074]); // EmitInputXorGate
assign xor0394 = (input_data[0087]^input_data[0086]^input_data[0083]^input_data[0082]); // EmitInputXorGate
assign xor0395 = (input_data[0095]^input_data[0094]^input_data[0091]^input_data[0090]); // EmitInputXorGate
assign xor0396 = (input_data[0103]^input_data[0102]^input_data[0099]^input_data[0098]); // EmitInputXorGate
assign xor0397 = (input_data[0107]^input_data[0111]^input_data[0106]^input_data[0110]); // EmitInputXorGate
assign xor0398 = (input_data[0114]^input_data[0119]^input_data[0118]^input_data[0115]); // EmitInputXorGate
assign xor0399 = (input_data[0127]^input_data[0126]^input_data[0123]^input_data[0122]); // EmitInputXorGate
assign xor0400 = (input_data[0131]^input_data[0130]^input_data[0135]^input_data[0134]); // EmitInputXorGate
assign xor0401 = (input_data[0139]^input_data[0138]^input_data[0143]^input_data[0142]); // EmitInputXorGate
assign xor0402 = (input_data[0147]^input_data[0151]^input_data[0150]^input_data[0146]); // EmitInputXorGate
assign xor0403 = (input_data[0159]^input_data[0158]^input_data[0155]^input_data[0154]); // EmitInputXorGate
assign xor0404 = (input_data[0167]^input_data[0166]^input_data[0163]^input_data[0162]); // EmitInputXorGate
assign xor0405 = (input_data[0175]^input_data[0174]^input_data[0171]^input_data[0170]); // EmitInputXorGate
assign xor0406 = (input_data[0183]^input_data[0182]^input_data[0179]^input_data[0178]); // EmitInputXorGate
assign xor0407 = (input_data[0187]^input_data[0186]^input_data[0191]^input_data[0190]); // EmitInputXorGate
assign xor0408 = (input_data[0199]^input_data[0198]^input_data[0195]^input_data[0194]); // EmitInputXorGate
assign xor0409 = (input_data[0207]^input_data[0206]^input_data[0203]^input_data[0202]); // EmitInputXorGate
assign xor0410 = (input_data[0215]^input_data[0214]^input_data[0211]^input_data[0210]); // EmitInputXorGate
assign xor0411 = (input_data[0223]^input_data[0222]^input_data[0219]^input_data[0218]); // EmitInputXorGate
assign xor0412 = (input_data[0231]^input_data[0227]^input_data[0226]^input_data[0230]); // EmitInputXorGate
assign xor0413 = (input_data[0239]^input_data[0238]^input_data[0235]^input_data[0234]); // EmitInputXorGate
assign xor0414 = (input_data[0242]^input_data[0247]^input_data[0246]^input_data[0243]); // EmitInputXorGate
assign xor0415 = (input_data[0255]^input_data[0254]^input_data[0251]^input_data[0250]); // EmitInputXorGate
assign xor0416 = (input_data[0259]^input_data[0258]^input_data[0263]^input_data[0262]); // EmitInputXorGate
assign xor0417 = (input_data[0267]^input_data[0271]^input_data[0266]^input_data[0270]); // EmitInputXorGate
assign xor0418 = (input_data[0278]^input_data[0275]^input_data[0274]^input_data[0279]); // EmitInputXorGate
assign xor0419 = (input_data[0287]^input_data[0286]^input_data[0283]^input_data[0282]); // EmitInputXorGate
assign xor0420 = (input_data[0291]^input_data[0290]^input_data[0295]^input_data[0294]); // EmitInputXorGate
assign xor0421 = (input_data[0303]^input_data[0302]^input_data[0299]^input_data[0298]); // EmitInputXorGate
assign xor0422 = (input_data[0310]^input_data[0307]^input_data[0311]^input_data[0306]); // EmitInputXorGate
assign xor0423 = (input_data[0319]^input_data[0318]^input_data[0315]^input_data[0314]); // EmitInputXorGate
assign xor0424 = (input_data[0322]^input_data[0327]^input_data[0326]^input_data[0323]); // EmitInputXorGate
assign xor0425 = (input_data[0335]^input_data[0334]^input_data[0331]^input_data[0330]); // EmitInputXorGate
assign xor0426 = (input_data[0339]^input_data[0338]^input_data[0343]^input_data[0342]); // EmitInputXorGate
assign xor0427 = (input_data[0351]^input_data[0347]^input_data[0346]^input_data[0350]); // EmitInputXorGate
assign xor0428 = (input_data[0355]^input_data[0354]^input_data[0359]^input_data[0358]); // EmitInputXorGate
assign xor0429 = (input_data[0367]^input_data[0366]^input_data[0363]^input_data[0362]); // EmitInputXorGate
assign xor0430 = (input_data[0371]^input_data[0370]^input_data[0375]^input_data[0374]); // EmitInputXorGate
assign xor0431 = (input_data[0383]^input_data[0382]^input_data[0379]^input_data[0378]); // EmitInputXorGate
assign xor0432 = (input_data[0387]^input_data[0391]^input_data[0386]^input_data[0390]); // EmitInputXorGate
assign xor0433 = (input_data[0399]^input_data[0398]^input_data[0395]^input_data[0394]); // EmitInputXorGate
assign xor0434 = (input_data[0407]^input_data[0406]^input_data[0403]^input_data[0402]); // EmitInputXorGate
assign xor0435 = (input_data[0411]^input_data[0410]^input_data[0415]^input_data[0414]); // EmitInputXorGate
assign xor0436 = (input_data[0423]^input_data[0422]^input_data[0419]^input_data[0418]); // EmitInputXorGate
assign xor0437 = (input_data[0430]^input_data[0426]^input_data[0427]^input_data[0431]); // EmitInputXorGate
assign xor0438 = (input_data[0439]^input_data[0438]^input_data[0435]^input_data[0434]); // EmitInputXorGate
assign xor0439 = (input_data[0447]^input_data[0446]^input_data[0443]^input_data[0442]); // EmitInputXorGate
assign xor0440 = (input_data[0455]^input_data[0454]^input_data[0451]^input_data[0450]); // EmitInputXorGate
assign xor0441 = (input_data[0459]^input_data[0458]^input_data[0463]^input_data[0462]); // EmitInputXorGate
assign xor0442 = (input_data[0467]^input_data[0471]^input_data[0466]^input_data[0470]); // EmitInputXorGate
assign xor0443 = (input_data[0475]^input_data[0474]^input_data[0479]^input_data[0478]); // EmitInputXorGate
assign xor0444 = (input_data[0486]^input_data[0483]^input_data[0482]^input_data[0487]); // EmitInputXorGate
assign xor0445 = (input_data[0491]^input_data[0490]^input_data[0495]^input_data[0494]); // EmitInputXorGate
assign xor0446 = (input_data[0503]^input_data[0502]^input_data[0499]^input_data[0498]); // EmitInputXorGate
assign xor0447 = (input_data[0507]^input_data[0511]^input_data[0506]^input_data[0510]); // EmitInputXorGate
assign xor0448 = (input_data[0519]^input_data[0518]^input_data[0515]^input_data[0514]); // EmitInputXorGate
assign xor0449 = (input_data[0527]^input_data[0526]^input_data[0523]^input_data[0522]); // EmitInputXorGate
assign xor0450 = (input_data[0535]^input_data[0534]^input_data[0531]^input_data[0530]); // EmitInputXorGate
assign xor0451 = (input_data[0539]^input_data[0538]^input_data[0543]^input_data[0542]); // EmitInputXorGate
assign xor0452 = (input_data[0551]^input_data[0547]^input_data[0550]^input_data[0546]); // EmitInputXorGate
assign xor0453 = (input_data[0554]^input_data[0559]^input_data[0558]^input_data[0555]); // EmitInputXorGate
assign xor0454 = (input_data[0567]^input_data[0566]^input_data[0563]^input_data[0562]); // EmitInputXorGate
assign xor0455 = (input_data[0571]^input_data[0570]^input_data[0575]^input_data[0574]); // EmitInputXorGate
assign xor0456 = (input_data[0579]^input_data[0578]^input_data[0583]^input_data[0582]); // EmitInputXorGate
assign xor0457 = (input_data[0587]^input_data[0591]^input_data[0586]^input_data[0590]); // EmitInputXorGate
assign xor0458 = (input_data[0599]^input_data[0598]^input_data[0595]^input_data[0594]); // EmitInputXorGate
assign xor0459 = (input_data[0603]^input_data[0602]^input_data[0607]^input_data[0606]); // EmitInputXorGate
assign xor0460 = (input_data[0615]^input_data[0614]^input_data[0611]^input_data[0610]); // EmitInputXorGate
assign xor0461 = (input_data[0619]^input_data[0618]^input_data[0623]^input_data[0622]); // EmitInputXorGate
assign xor0462 = (input_data[0627]^input_data[0631]^input_data[0626]^input_data[0630]); // EmitInputXorGate
assign xor0463 = (input_data[0639]^input_data[0638]^input_data[0635]^input_data[0634]); // EmitInputXorGate
assign xor0464 = (input_data[0647]^input_data[0646]^input_data[0643]^input_data[0642]); // EmitInputXorGate
assign xor0465 = (input_data[0655]^input_data[0654]^input_data[0651]^input_data[0650]); // EmitInputXorGate
assign xor0466 = (input_data[0663]^input_data[0662]^input_data[0659]^input_data[0658]); // EmitInputXorGate
assign xor0467 = (input_data[0671]^input_data[0667]^input_data[0666]^input_data[0670]); // EmitInputXorGate
assign xor0468 = (input_data[0679]^input_data[0678]^input_data[0675]^input_data[0674]); // EmitInputXorGate
assign xor0469 = (input_data[0682]^input_data[0687]^input_data[0686]^input_data[0683]); // EmitInputXorGate
assign xor0470 = (input_data[0695]^input_data[0694]^input_data[0691]^input_data[0690]); // EmitInputXorGate
assign xor0471 = (input_data[0699]^input_data[0698]^input_data[0703]^input_data[0702]); // EmitInputXorGate
assign xor0472 = (input_data[0707]^input_data[0711]^input_data[0710]^input_data[0706]); // EmitInputXorGate
assign xor0473 = (input_data[0719]^input_data[0718]^input_data[0715]^input_data[0714]); // EmitInputXorGate
assign xor0474 = (input_data[0727]^input_data[0726]^input_data[0723]^input_data[0722]); // EmitInputXorGate
assign xor0475 = (input_data[0735]^input_data[0734]^input_data[0731]^input_data[0730]); // EmitInputXorGate
assign xor0476 = (input_data[0743]^input_data[0742]^input_data[0739]^input_data[0738]); // EmitInputXorGate
assign xor0477 = (input_data[0750]^input_data[0747]^input_data[0751]^input_data[0746]); // EmitInputXorGate
assign xor0478 = (input_data[0759]^input_data[0758]^input_data[0755]^input_data[0754]); // EmitInputXorGate
assign xor0479 = (input_data[0762]^input_data[0767]^input_data[0766]^input_data[0763]); // EmitInputXorGate
assign xor0480 = (input_data[0775]^input_data[0774]^input_data[0771]^input_data[0770]); // EmitInputXorGate
assign xor0481 = (input_data[0779]^input_data[0778]^input_data[0783]^input_data[0782]); // EmitInputXorGate
assign xor0482 = (input_data[0791]^input_data[0787]^input_data[0786]^input_data[0790]); // EmitInputXorGate
assign xor0483 = (input_data[0795]^input_data[0794]^input_data[0799]^input_data[0798]); // EmitInputXorGate
assign xor0484 = (input_data[0803]^input_data[0802]^input_data[0807]^input_data[0806]); // EmitInputXorGate
assign xor0485 = (input_data[0815]^input_data[0814]^input_data[0811]^input_data[0810]); // EmitInputXorGate
assign xor0486 = (input_data[0819]^input_data[0818]^input_data[0823]^input_data[0822]); // EmitInputXorGate
assign xor0487 = (input_data[0827]^input_data[0831]^input_data[0826]^input_data[0830]); // EmitInputXorGate
assign xor0488 = (input_data[0839]^input_data[0838]^input_data[0835]^input_data[0834]); // EmitInputXorGate
assign xor0489 = (input_data[0847]^input_data[0846]^input_data[0843]^input_data[0842]); // EmitInputXorGate
assign xor0490 = (input_data[0851]^input_data[0850]^input_data[0855]^input_data[0854]); // EmitInputXorGate
assign xor0491 = (input_data[0863]^input_data[0862]^input_data[0859]^input_data[0858]); // EmitInputXorGate
assign xor0492 = (input_data[0870]^input_data[0866]^input_data[0867]^input_data[0871]); // EmitInputXorGate
assign xor0493 = (input_data[0879]^input_data[0878]^input_data[0875]^input_data[0874]); // EmitInputXorGate
assign xor0494 = (input_data[0887]^input_data[0886]^input_data[0883]^input_data[0882]); // EmitInputXorGate
assign xor0495 = (input_data[0895]^input_data[0894]^input_data[0891]^input_data[0890]); // EmitInputXorGate
assign xor0496 = (input_data[0899]^input_data[0898]^input_data[0903]^input_data[0902]); // EmitInputXorGate
assign xor0497 = (input_data[0907]^input_data[0911]^input_data[0906]^input_data[0910]); // EmitInputXorGate
assign xor0498 = (input_data[0915]^input_data[0914]^input_data[0919]^input_data[0918]); // EmitInputXorGate
assign xor0499 = (input_data[0927]^input_data[0926]^input_data[0923]^input_data[0922]); // EmitInputXorGate
assign xor0500 = (input_data[0934]^input_data[0931]^input_data[0930]^input_data[0935]); // EmitInputXorGate
assign xor0501 = (input_data[0943]^input_data[0942]^input_data[0939]^input_data[0938]); // EmitInputXorGate
assign xor0502 = (input_data[0947]^input_data[0951]^input_data[0946]^input_data[0950]); // EmitInputXorGate
assign xor0503 = (input_data[0959]^input_data[0958]^input_data[0955]^input_data[0954]); // EmitInputXorGate
assign xor0504 = (input_data[0967]^input_data[0966]^input_data[0963]^input_data[0962]); // EmitInputXorGate
assign xor0505 = (input_data[0975]^input_data[0974]^input_data[0971]^input_data[0970]); // EmitInputXorGate
assign xor0506 = (input_data[0979]^input_data[0978]^input_data[0983]^input_data[0982]); // EmitInputXorGate
assign xor0507 = (input_data[0987]^input_data[0991]^input_data[0990]^input_data[0986]); // EmitInputXorGate
assign xor0508 = (input_data[0994]^input_data[0999]^input_data[0998]^input_data[0995]); // EmitInputXorGate
assign xor0509 = (input_data[1007]^input_data[1006]^input_data[1003]^input_data[1002]); // EmitInputXorGate
assign xor0510 = (input_data[1015]^input_data[1014]^input_data[1011]^input_data[1010]); // EmitInputXorGate
assign xor0511 = (input_data[1023]^input_data[1022]^input_data[1019]^input_data[1018]); // EmitInputXorGate
// BuildXorTrees, FirstLevel, f = 2
assign xor0512 = (input_data[0005]^input_data[0004]^input_data[0007]^input_data[0006]); // EmitInputXorGate
assign xor0513 = (input_data[0015]^input_data[0014]^input_data[0013]^input_data[0012]); // EmitInputXorGate
assign xor0514 = (input_data[0021]^input_data[0020]^input_data[0023]^input_data[0022]); // EmitInputXorGate
assign xor0515 = (input_data[0028]^input_data[0031]^input_data[0030]^input_data[0029]); // EmitInputXorGate
assign xor0516 = (input_data[0037]^input_data[0036]^input_data[0039]^input_data[0038]); // EmitInputXorGate
assign xor0517 = (input_data[0046]^input_data[0045]^input_data[0044]^input_data[0047]); // EmitInputXorGate
assign xor0518 = (input_data[0053]^input_data[0052]^input_data[0055]^input_data[0054]); // EmitInputXorGate
assign xor0519 = (input_data[0063]^input_data[0062]^input_data[0061]^input_data[0060]); // EmitInputXorGate
assign xor0520 = (input_data[0069]^input_data[0068]^input_data[0071]^input_data[0070]); // EmitInputXorGate
assign xor0521 = (input_data[0079]^input_data[0078]^input_data[0077]^input_data[0076]); // EmitInputXorGate
assign xor0522 = (input_data[0085]^input_data[0084]^input_data[0087]^input_data[0086]); // EmitInputXorGate
assign xor0523 = (input_data[0095]^input_data[0094]^input_data[0093]^input_data[0092]); // EmitInputXorGate
assign xor0524 = (input_data[0101]^input_data[0100]^input_data[0103]^input_data[0102]); // EmitInputXorGate
assign xor0525 = (input_data[0111]^input_data[0110]^input_data[0109]^input_data[0108]); // EmitInputXorGate
assign xor0526 = (input_data[0117]^input_data[0116]^input_data[0119]^input_data[0118]); // EmitInputXorGate
assign xor0527 = (input_data[0127]^input_data[0126]^input_data[0125]^input_data[0124]); // EmitInputXorGate
assign xor0528 = (input_data[0133]^input_data[0132]^input_data[0135]^input_data[0134]); // EmitInputXorGate
assign xor0529 = (input_data[0141]^input_data[0140]^input_data[0143]^input_data[0142]); // EmitInputXorGate
assign xor0530 = (input_data[0149]^input_data[0148]^input_data[0151]^input_data[0150]); // EmitInputXorGate
assign xor0531 = (input_data[0159]^input_data[0158]^input_data[0157]^input_data[0156]); // EmitInputXorGate
assign xor0532 = (input_data[0165]^input_data[0164]^input_data[0167]^input_data[0166]); // EmitInputXorGate
assign xor0533 = (input_data[0175]^input_data[0174]^input_data[0173]^input_data[0172]); // EmitInputXorGate
assign xor0534 = (input_data[0181]^input_data[0180]^input_data[0183]^input_data[0182]); // EmitInputXorGate
assign xor0535 = (input_data[0191]^input_data[0190]^input_data[0189]^input_data[0188]); // EmitInputXorGate
assign xor0536 = (input_data[0196]^input_data[0199]^input_data[0198]^input_data[0197]); // EmitInputXorGate
assign xor0537 = (input_data[0205]^input_data[0204]^input_data[0207]^input_data[0206]); // EmitInputXorGate
assign xor0538 = (input_data[0215]^input_data[0214]^input_data[0213]^input_data[0212]); // EmitInputXorGate
assign xor0539 = (input_data[0221]^input_data[0220]^input_data[0223]^input_data[0222]); // EmitInputXorGate
assign xor0540 = (input_data[0231]^input_data[0230]^input_data[0229]^input_data[0228]); // EmitInputXorGate
assign xor0541 = (input_data[0236]^input_data[0239]^input_data[0238]^input_data[0237]); // EmitInputXorGate
assign xor0542 = (input_data[0245]^input_data[0244]^input_data[0247]^input_data[0246]); // EmitInputXorGate
assign xor0543 = (input_data[0255]^input_data[0254]^input_data[0253]^input_data[0252]); // EmitInputXorGate
assign xor0544 = (input_data[0261]^input_data[0260]^input_data[0263]^input_data[0262]); // EmitInputXorGate
assign xor0545 = (input_data[0269]^input_data[0268]^input_data[0271]^input_data[0270]); // EmitInputXorGate
assign xor0546 = (input_data[0278]^input_data[0277]^input_data[0276]^input_data[0279]); // EmitInputXorGate
assign xor0547 = (input_data[0284]^input_data[0287]^input_data[0286]^input_data[0285]); // EmitInputXorGate
assign xor0548 = (input_data[0293]^input_data[0292]^input_data[0295]^input_data[0294]); // EmitInputXorGate
assign xor0549 = (input_data[0301]^input_data[0300]^input_data[0303]^input_data[0302]); // EmitInputXorGate
assign xor0550 = (input_data[0310]^input_data[0309]^input_data[0308]^input_data[0311]); // EmitInputXorGate
assign xor0551 = (input_data[0319]^input_data[0318]^input_data[0317]^input_data[0316]); // EmitInputXorGate
assign xor0552 = (input_data[0325]^input_data[0324]^input_data[0327]^input_data[0326]); // EmitInputXorGate
assign xor0553 = (input_data[0335]^input_data[0334]^input_data[0333]^input_data[0332]); // EmitInputXorGate
assign xor0554 = (input_data[0341]^input_data[0340]^input_data[0343]^input_data[0342]); // EmitInputXorGate
assign xor0555 = (input_data[0348]^input_data[0351]^input_data[0350]^input_data[0349]); // EmitInputXorGate
assign xor0556 = (input_data[0357]^input_data[0356]^input_data[0359]^input_data[0358]); // EmitInputXorGate
assign xor0557 = (input_data[0365]^input_data[0364]^input_data[0367]^input_data[0366]); // EmitInputXorGate
assign xor0558 = (input_data[0373]^input_data[0372]^input_data[0375]^input_data[0374]); // EmitInputXorGate
assign xor0559 = (input_data[0383]^input_data[0382]^input_data[0381]^input_data[0380]); // EmitInputXorGate
assign xor0560 = (input_data[0389]^input_data[0388]^input_data[0391]^input_data[0390]); // EmitInputXorGate
assign xor0561 = (input_data[0399]^input_data[0398]^input_data[0397]^input_data[0396]); // EmitInputXorGate
assign xor0562 = (input_data[0405]^input_data[0404]^input_data[0407]^input_data[0406]); // EmitInputXorGate
assign xor0563 = (input_data[0413]^input_data[0412]^input_data[0415]^input_data[0414]); // EmitInputXorGate
assign xor0564 = (input_data[0421]^input_data[0420]^input_data[0423]^input_data[0422]); // EmitInputXorGate
assign xor0565 = (input_data[0430]^input_data[0429]^input_data[0428]^input_data[0431]); // EmitInputXorGate
assign xor0566 = (input_data[0439]^input_data[0438]^input_data[0437]^input_data[0436]); // EmitInputXorGate
assign xor0567 = (input_data[0445]^input_data[0444]^input_data[0447]^input_data[0446]); // EmitInputXorGate
assign xor0568 = (input_data[0455]^input_data[0454]^input_data[0453]^input_data[0452]); // EmitInputXorGate
assign xor0569 = (input_data[0461]^input_data[0460]^input_data[0463]^input_data[0462]); // EmitInputXorGate
assign xor0570 = (input_data[0468]^input_data[0471]^input_data[0470]^input_data[0469]); // EmitInputXorGate
assign xor0571 = (input_data[0477]^input_data[0476]^input_data[0479]^input_data[0478]); // EmitInputXorGate
assign xor0572 = (input_data[0486]^input_data[0485]^input_data[0484]^input_data[0487]); // EmitInputXorGate
assign xor0573 = (input_data[0493]^input_data[0492]^input_data[0495]^input_data[0494]); // EmitInputXorGate
assign xor0574 = (input_data[0500]^input_data[0503]^input_data[0502]^input_data[0501]); // EmitInputXorGate
assign xor0575 = (input_data[0509]^input_data[0508]^input_data[0511]^input_data[0510]); // EmitInputXorGate
assign xor0576 = (input_data[0519]^input_data[0518]^input_data[0517]^input_data[0516]); // EmitInputXorGate
assign xor0577 = (input_data[0525]^input_data[0524]^input_data[0527]^input_data[0526]); // EmitInputXorGate
assign xor0578 = (input_data[0535]^input_data[0534]^input_data[0533]^input_data[0532]); // EmitInputXorGate
assign xor0579 = (input_data[0541]^input_data[0540]^input_data[0543]^input_data[0542]); // EmitInputXorGate
assign xor0580 = (input_data[0551]^input_data[0550]^input_data[0549]^input_data[0548]); // EmitInputXorGate
assign xor0581 = (input_data[0557]^input_data[0556]^input_data[0559]^input_data[0558]); // EmitInputXorGate
assign xor0582 = (input_data[0567]^input_data[0566]^input_data[0565]^input_data[0564]); // EmitInputXorGate
assign xor0583 = (input_data[0573]^input_data[0572]^input_data[0575]^input_data[0574]); // EmitInputXorGate
assign xor0584 = (input_data[0581]^input_data[0580]^input_data[0583]^input_data[0582]); // EmitInputXorGate
assign xor0585 = (input_data[0589]^input_data[0588]^input_data[0591]^input_data[0590]); // EmitInputXorGate
assign xor0586 = (input_data[0599]^input_data[0598]^input_data[0597]^input_data[0596]); // EmitInputXorGate
assign xor0587 = (input_data[0605]^input_data[0604]^input_data[0607]^input_data[0606]); // EmitInputXorGate
assign xor0588 = (input_data[0613]^input_data[0612]^input_data[0615]^input_data[0614]); // EmitInputXorGate
assign xor0589 = (input_data[0621]^input_data[0620]^input_data[0623]^input_data[0622]); // EmitInputXorGate
assign xor0590 = (input_data[0629]^input_data[0628]^input_data[0631]^input_data[0630]); // EmitInputXorGate
assign xor0591 = (input_data[0639]^input_data[0638]^input_data[0637]^input_data[0636]); // EmitInputXorGate
assign xor0592 = (input_data[0645]^input_data[0644]^input_data[0647]^input_data[0646]); // EmitInputXorGate
assign xor0593 = (input_data[0655]^input_data[0654]^input_data[0653]^input_data[0652]); // EmitInputXorGate
assign xor0594 = (input_data[0661]^input_data[0660]^input_data[0663]^input_data[0662]); // EmitInputXorGate
assign xor0595 = (input_data[0671]^input_data[0670]^input_data[0669]^input_data[0668]); // EmitInputXorGate
assign xor0596 = (input_data[0676]^input_data[0679]^input_data[0678]^input_data[0677]); // EmitInputXorGate
assign xor0597 = (input_data[0685]^input_data[0684]^input_data[0687]^input_data[0686]); // EmitInputXorGate
assign xor0598 = (input_data[0695]^input_data[0694]^input_data[0693]^input_data[0692]); // EmitInputXorGate
assign xor0599 = (input_data[0701]^input_data[0700]^input_data[0703]^input_data[0702]); // EmitInputXorGate
assign xor0600 = (input_data[0709]^input_data[0708]^input_data[0711]^input_data[0710]); // EmitInputXorGate
assign xor0601 = (input_data[0719]^input_data[0718]^input_data[0717]^input_data[0716]); // EmitInputXorGate
assign xor0602 = (input_data[0725]^input_data[0724]^input_data[0727]^input_data[0726]); // EmitInputXorGate
assign xor0603 = (input_data[0735]^input_data[0734]^input_data[0733]^input_data[0732]); // EmitInputXorGate
assign xor0604 = (input_data[0741]^input_data[0740]^input_data[0743]^input_data[0742]); // EmitInputXorGate
assign xor0605 = (input_data[0750]^input_data[0749]^input_data[0748]^input_data[0751]); // EmitInputXorGate
assign xor0606 = (input_data[0759]^input_data[0758]^input_data[0757]^input_data[0756]); // EmitInputXorGate
assign xor0607 = (input_data[0765]^input_data[0764]^input_data[0767]^input_data[0766]); // EmitInputXorGate
assign xor0608 = (input_data[0775]^input_data[0774]^input_data[0773]^input_data[0772]); // EmitInputXorGate
assign xor0609 = (input_data[0781]^input_data[0780]^input_data[0783]^input_data[0782]); // EmitInputXorGate
assign xor0610 = (input_data[0788]^input_data[0791]^input_data[0790]^input_data[0789]); // EmitInputXorGate
assign xor0611 = (input_data[0797]^input_data[0796]^input_data[0799]^input_data[0798]); // EmitInputXorGate
assign xor0612 = (input_data[0805]^input_data[0804]^input_data[0807]^input_data[0806]); // EmitInputXorGate
assign xor0613 = (input_data[0815]^input_data[0814]^input_data[0813]^input_data[0812]); // EmitInputXorGate
assign xor0614 = (input_data[0821]^input_data[0820]^input_data[0823]^input_data[0822]); // EmitInputXorGate
assign xor0615 = (input_data[0829]^input_data[0828]^input_data[0831]^input_data[0830]); // EmitInputXorGate
assign xor0616 = (input_data[0839]^input_data[0838]^input_data[0837]^input_data[0836]); // EmitInputXorGate
assign xor0617 = (input_data[0845]^input_data[0844]^input_data[0847]^input_data[0846]); // EmitInputXorGate
assign xor0618 = (input_data[0853]^input_data[0852]^input_data[0855]^input_data[0854]); // EmitInputXorGate
assign xor0619 = (input_data[0861]^input_data[0860]^input_data[0863]^input_data[0862]); // EmitInputXorGate
assign xor0620 = (input_data[0870]^input_data[0869]^input_data[0868]^input_data[0871]); // EmitInputXorGate
assign xor0621 = (input_data[0879]^input_data[0878]^input_data[0877]^input_data[0876]); // EmitInputXorGate
assign xor0622 = (input_data[0885]^input_data[0884]^input_data[0887]^input_data[0886]); // EmitInputXorGate
assign xor0623 = (input_data[0895]^input_data[0894]^input_data[0893]^input_data[0892]); // EmitInputXorGate
assign xor0624 = (input_data[0901]^input_data[0900]^input_data[0903]^input_data[0902]); // EmitInputXorGate
assign xor0625 = (input_data[0908]^input_data[0911]^input_data[0910]^input_data[0909]); // EmitInputXorGate
assign xor0626 = (input_data[0917]^input_data[0916]^input_data[0919]^input_data[0918]); // EmitInputXorGate
assign xor0627 = (input_data[0925]^input_data[0924]^input_data[0927]^input_data[0926]); // EmitInputXorGate
assign xor0628 = (input_data[0934]^input_data[0933]^input_data[0932]^input_data[0935]); // EmitInputXorGate
assign xor0629 = (input_data[0943]^input_data[0942]^input_data[0941]^input_data[0940]); // EmitInputXorGate
assign xor0630 = (input_data[0949]^input_data[0948]^input_data[0951]^input_data[0950]); // EmitInputXorGate
assign xor0631 = (input_data[0959]^input_data[0958]^input_data[0957]^input_data[0956]); // EmitInputXorGate
assign xor0632 = (input_data[0965]^input_data[0964]^input_data[0967]^input_data[0966]); // EmitInputXorGate
assign xor0633 = (input_data[0975]^input_data[0974]^input_data[0973]^input_data[0972]); // EmitInputXorGate
assign xor0634 = (input_data[0981]^input_data[0980]^input_data[0983]^input_data[0982]); // EmitInputXorGate
assign xor0635 = (input_data[0991]^input_data[0990]^input_data[0989]^input_data[0988]); // EmitInputXorGate
assign xor0636 = (input_data[0997]^input_data[0996]^input_data[0999]^input_data[0998]); // EmitInputXorGate
assign xor0637 = (input_data[1005]^input_data[1004]^input_data[1007]^input_data[1006]); // EmitInputXorGate
assign xor0638 = (input_data[1015]^input_data[1014]^input_data[1013]^input_data[1012]); // EmitInputXorGate
assign xor0639 = (input_data[1021]^input_data[1020]^input_data[1023]^input_data[1022]); // EmitInputXorGate
// BuildXorTrees, ParityBits, i = 0
assign xor0640 = (xor0257^xor0258^xor0256^xor0259); // MakeXorFrom
assign xor0641 = (xor0260^xor0263^xor0261^xor0262); // MakeXorFrom
assign xor0642 = (xor0265^xor0266^xor0264^xor0267); // MakeXorFrom
assign xor0643 = (xor0270^xor0268^xor0271^xor0269); // MakeXorFrom
assign xor0644 = (xor0275^xor0273^xor0274^xor0272); // MakeXorFrom
assign xor0645 = (xor0278^xor0276^xor0279^xor0277); // MakeXorFrom
assign xor0646 = (xor0283^xor0281^xor0282^xor0280); // MakeXorFrom
assign xor0647 = (xor0285^xor0286^xor0284^xor0287); // MakeXorFrom
assign xor0648 = (xor0288^xor0291^xor0289^xor0290); // MakeXorFrom
assign xor0649 = (xor0295^xor0293^xor0294^xor0292); // MakeXorFrom
assign xor0650 = (xor0296^xor0299^xor0297^xor0298); // MakeXorFrom
assign xor0651 = (xor0302^xor0300^xor0303^xor0301); // MakeXorFrom
assign xor0652 = (xor0307^xor0305^xor0306^xor0304); // MakeXorFrom
assign xor0653 = (xor0309^xor0310^xor0308^xor0311); // MakeXorFrom
assign xor0654 = (xor0312^xor0315^xor0313^xor0314); // MakeXorFrom
assign xor0655 = (xor0317^xor0318^xor0316^xor0319); // MakeXorFrom
assign xor0656 = (xor0322^xor0320^xor0323^xor0321); // MakeXorFrom
assign xor0657 = (xor0327^xor0325^xor0326^xor0324); // MakeXorFrom
assign xor0658 = (xor0330^xor0328^xor0331^xor0329); // MakeXorFrom
assign xor0659 = (xor0335^xor0333^xor0334^xor0332); // MakeXorFrom
assign xor0660 = (xor0337^xor0338^xor0336^xor0339); // MakeXorFrom
assign xor0661 = (xor0340^xor0343^xor0341^xor0342); // MakeXorFrom
assign xor0662 = (xor0347^xor0345^xor0346^xor0344); // MakeXorFrom
assign xor0663 = (xor0350^xor0348^xor0351^xor0349); // MakeXorFrom
assign xor0664 = (xor0355^xor0353^xor0354^xor0352); // MakeXorFrom
assign xor0665 = (xor0358^xor0356^xor0359^xor0357); // MakeXorFrom
assign xor0666 = (xor0363^xor0361^xor0362^xor0360); // MakeXorFrom
assign xor0667 = (xor0365^xor0366^xor0364^xor0367); // MakeXorFrom
assign xor0668 = (xor0368^xor0371^xor0369^xor0370); // MakeXorFrom
assign xor0669 = (xor0375^xor0373^xor0374^xor0372); // MakeXorFrom
assign xor0670 = (xor0376^xor0379^xor0377^xor0378); // MakeXorFrom
assign xor0671 = (xor0383^xor0381^xor0382^xor0380); // MakeXorFrom
assign xor0672 = (xor0643^xor0641^xor0642^xor0640); // MakeXorFrom
assign xor0673 = (xor0644^xor0647^xor0645^xor0646); // MakeXorFrom
assign xor0674 = (xor0651^xor0649^xor0650^xor0648); // MakeXorFrom
assign xor0675 = (xor0654^xor0652^xor0655^xor0653); // MakeXorFrom
assign xor0676 = (xor0659^xor0657^xor0658^xor0656); // MakeXorFrom
assign xor0677 = (xor0661^xor0662^xor0660^xor0663); // MakeXorFrom
assign xor0678 = (xor0664^xor0667^xor0665^xor0666); // MakeXorFrom
assign xor0679 = (xor0671^xor0669^xor0670^xor0668); // MakeXorFrom
assign xor0680 = (xor0672^xor0675^xor0673^xor0674); // MakeXorFrom
assign xor0681 = (xor0679^xor0677^xor0678^xor0676); // MakeXorFrom
assign xor0682 = (xor0680^xor0681); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 1
assign xor0683 = (xor0386^xor0384^xor0387^xor0385); // MakeXorFrom
assign xor0684 = (xor0391^xor0389^xor0390^xor0388); // MakeXorFrom
assign xor0685 = (xor0393^xor0394^xor0392^xor0395); // MakeXorFrom
assign xor0686 = (xor0396^xor0399^xor0397^xor0398); // MakeXorFrom
assign xor0687 = (xor0403^xor0401^xor0402^xor0400); // MakeXorFrom
assign xor0688 = (xor0404^xor0407^xor0405^xor0406); // MakeXorFrom
assign xor0689 = (xor0411^xor0409^xor0410^xor0408); // MakeXorFrom
assign xor0690 = (xor0414^xor0412^xor0415^xor0413); // MakeXorFrom
assign xor0691 = (xor0419^xor0417^xor0418^xor0416); // MakeXorFrom
assign xor0692 = (xor0421^xor0422^xor0420^xor0423); // MakeXorFrom
assign xor0693 = (xor0424^xor0427^xor0425^xor0426); // MakeXorFrom
assign xor0694 = (xor0431^xor0429^xor0430^xor0428); // MakeXorFrom
assign xor0695 = (xor0434^xor0432^xor0435^xor0433); // MakeXorFrom
assign xor0696 = (xor0439^xor0437^xor0438^xor0436); // MakeXorFrom
assign xor0697 = (xor0441^xor0442^xor0440^xor0443); // MakeXorFrom
assign xor0698 = (xor0447^xor0445^xor0446^xor0444); // MakeXorFrom
assign xor0699 = (xor0449^xor0450^xor0448^xor0451); // MakeXorFrom
assign xor0700 = (xor0452^xor0455^xor0453^xor0454); // MakeXorFrom
assign xor0701 = (xor0459^xor0457^xor0458^xor0456); // MakeXorFrom
assign xor0702 = (xor0462^xor0460^xor0463^xor0461); // MakeXorFrom
assign xor0703 = (xor0467^xor0465^xor0466^xor0464); // MakeXorFrom
assign xor0704 = (xor0470^xor0468^xor0471^xor0469); // MakeXorFrom
assign xor0705 = (xor0475^xor0473^xor0474^xor0472); // MakeXorFrom
assign xor0706 = (xor0477^xor0478^xor0476^xor0479); // MakeXorFrom
assign xor0707 = (xor0480^xor0483^xor0481^xor0482); // MakeXorFrom
assign xor0708 = (xor0487^xor0485^xor0486^xor0484); // MakeXorFrom
assign xor0709 = (xor0490^xor0488^xor0491^xor0489); // MakeXorFrom
assign xor0710 = (xor0495^xor0493^xor0494^xor0492); // MakeXorFrom
assign xor0711 = (xor0498^xor0496^xor0499^xor0497); // MakeXorFrom
assign xor0712 = (xor0501^xor0502^xor0500^xor0503); // MakeXorFrom
assign xor0713 = (xor0504^xor0507^xor0505^xor0506); // MakeXorFrom
assign xor0714 = (xor0511^xor0509^xor0510^xor0508); // MakeXorFrom
assign xor0715 = (xor0685^xor0686^xor0683^xor0684); // MakeXorFrom
assign xor0716 = (xor0689^xor0690^xor0687^xor0688); // MakeXorFrom
assign xor0717 = (xor0692^xor0693^xor0694^xor0691); // MakeXorFrom
assign xor0718 = (xor0697^xor0698^xor0695^xor0696); // MakeXorFrom
assign xor0719 = (xor0701^xor0702^xor0700^xor0699); // MakeXorFrom
assign xor0720 = (xor0706^xor0703^xor0704^xor0705); // MakeXorFrom
assign xor0721 = (xor0709^xor0710^xor0707^xor0708); // MakeXorFrom
assign xor0722 = (xor0713^xor0714^xor0711^xor0712); // MakeXorFrom
assign xor0723 = (xor0716^xor0717^xor0718^xor0715); // MakeXorFrom
assign xor0724 = (xor0721^xor0722^xor0719^xor0720); // MakeXorFrom
assign xor0725 = (xor0723^xor0724); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 2
assign xor0726 = (xor0514^xor0512^xor0515^xor0513); // MakeXorFrom
assign xor0727 = (xor0519^xor0517^xor0518^xor0516); // MakeXorFrom
assign xor0728 = (xor0521^xor0522^xor0520^xor0523); // MakeXorFrom
assign xor0729 = (xor0527^xor0525^xor0526^xor0524); // MakeXorFrom
assign xor0730 = (xor0529^xor0530^xor0528^xor0531); // MakeXorFrom
assign xor0731 = (xor0532^xor0535^xor0533^xor0534); // MakeXorFrom
assign xor0732 = (xor0539^xor0537^xor0538^xor0536); // MakeXorFrom
assign xor0733 = (xor0542^xor0540^xor0543^xor0541); // MakeXorFrom
assign xor0734 = (xor0547^xor0545^xor0546^xor0544); // MakeXorFrom
assign xor0735 = (xor0550^xor0548^xor0551^xor0549); // MakeXorFrom
assign xor0736 = (xor0552^xor0555^xor0553^xor0554); // MakeXorFrom
assign xor0737 = (xor0557^xor0558^xor0556^xor0559); // MakeXorFrom
assign xor0738 = (xor0560^xor0563^xor0561^xor0562); // MakeXorFrom
assign xor0739 = (xor0567^xor0565^xor0566^xor0564); // MakeXorFrom
assign xor0740 = (xor0570^xor0568^xor0571^xor0569); // MakeXorFrom
assign xor0741 = (xor0575^xor0573^xor0574^xor0572); // MakeXorFrom
assign xor0742 = (xor0577^xor0578^xor0576^xor0579); // MakeXorFrom
assign xor0743 = (xor0580^xor0583^xor0581^xor0582); // MakeXorFrom
assign xor0744 = (xor0585^xor0586^xor0584^xor0587); // MakeXorFrom
assign xor0745 = (xor0588^xor0591^xor0589^xor0590); // MakeXorFrom
assign xor0746 = (xor0595^xor0593^xor0594^xor0592); // MakeXorFrom
assign xor0747 = (xor0598^xor0596^xor0599^xor0597); // MakeXorFrom
assign xor0748 = (xor0603^xor0601^xor0602^xor0600); // MakeXorFrom
assign xor0749 = (xor0605^xor0606^xor0604^xor0607); // MakeXorFrom
assign xor0750 = (xor0611^xor0609^xor0610^xor0608); // MakeXorFrom
assign xor0751 = (xor0613^xor0614^xor0612^xor0615); // MakeXorFrom
assign xor0752 = (xor0616^xor0619^xor0617^xor0618); // MakeXorFrom
assign xor0753 = (xor0623^xor0621^xor0622^xor0620); // MakeXorFrom
assign xor0754 = (xor0626^xor0624^xor0627^xor0625); // MakeXorFrom
assign xor0755 = (xor0631^xor0629^xor0630^xor0628); // MakeXorFrom
assign xor0756 = (xor0633^xor0634^xor0632^xor0635); // MakeXorFrom
assign xor0757 = (xor0639^xor0637^xor0638^xor0636); // MakeXorFrom
assign xor0758 = (xor0729^xor0727^xor0728^xor0726); // MakeXorFrom
assign xor0759 = (xor0731^xor0732^xor0730^xor0733); // MakeXorFrom
assign xor0760 = (xor0734^xor0737^xor0735^xor0736); // MakeXorFrom
assign xor0761 = (xor0741^xor0739^xor0740^xor0738); // MakeXorFrom
assign xor0762 = (xor0744^xor0742^xor0745^xor0743); // MakeXorFrom
assign xor0763 = (xor0749^xor0747^xor0748^xor0746); // MakeXorFrom
assign xor0764 = (xor0751^xor0752^xor0750^xor0753); // MakeXorFrom
assign xor0765 = (xor0757^xor0755^xor0756^xor0754); // MakeXorFrom
assign xor0766 = (xor0761^xor0759^xor0760^xor0758); // MakeXorFrom
assign xor0767 = (xor0762^xor0765^xor0763^xor0764); // MakeXorFrom
assign xor0768 = (xor0767^xor0766); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 3
assign xor0769 = (xor0002^xor0010^xor0006^xor0014); // MakeXorFrom
assign xor0770 = (xor0030^xor0018^xor0026^xor0022); // MakeXorFrom
assign xor0771 = (xor0038^xor0046^xor0034^xor0042); // MakeXorFrom
assign xor0772 = (xor0054^xor0062^xor0058^xor0050); // MakeXorFrom
assign xor0773 = (xor0066^xor0074^xor0078^xor0070); // MakeXorFrom
assign xor0774 = (xor0086^xor0094^xor0082^xor0090); // MakeXorFrom
assign xor0775 = (xor0110^xor0106^xor0098^xor0102); // MakeXorFrom
assign xor0776 = (xor0118^xor0126^xor0114^xor0122); // MakeXorFrom
assign xor0777 = (xor0138^xor0134^xor0142^xor0130); // MakeXorFrom
assign xor0778 = (xor0146^xor0154^xor0150^xor0158); // MakeXorFrom
assign xor0779 = (xor0166^xor0174^xor0162^xor0170); // MakeXorFrom
assign xor0780 = (xor0182^xor0190^xor0178^xor0186); // MakeXorFrom
assign xor0781 = (xor0194^xor0202^xor0198^xor0206); // MakeXorFrom
assign xor0782 = (xor0222^xor0210^xor0218^xor0214); // MakeXorFrom
assign xor0783 = (xor0230^xor0238^xor0226^xor0234); // MakeXorFrom
assign xor0784 = (xor0250^xor0246^xor0254^xor0242); // MakeXorFrom
assign xor0785 = (xor0519^xor0517^xor0515^xor0513); // MakeXorFrom
assign xor0786 = (xor0521^xor0527^xor0525^xor0523); // MakeXorFrom
assign xor0787 = (xor0529^xor0535^xor0533^xor0531); // MakeXorFrom
assign xor0788 = (xor0539^xor0537^xor0543^xor0541); // MakeXorFrom
assign xor0789 = (xor0547^xor0545^xor0551^xor0549); // MakeXorFrom
assign xor0790 = (xor0557^xor0555^xor0553^xor0559); // MakeXorFrom
assign xor0791 = (xor0567^xor0565^xor0563^xor0561); // MakeXorFrom
assign xor0792 = (xor0575^xor0573^xor0571^xor0569); // MakeXorFrom
assign xor0793 = (xor0577^xor0583^xor0581^xor0579); // MakeXorFrom
assign xor0794 = (xor0585^xor0591^xor0589^xor0587); // MakeXorFrom
assign xor0795 = (xor0595^xor0593^xor0599^xor0597); // MakeXorFrom
assign xor0796 = (xor0605^xor0603^xor0601^xor0607); // MakeXorFrom
assign xor0797 = (xor0613^xor0611^xor0609^xor0615); // MakeXorFrom
assign xor0798 = (xor0623^xor0621^xor0619^xor0617); // MakeXorFrom
assign xor0799 = (xor0631^xor0629^xor0627^xor0625); // MakeXorFrom
assign xor0800 = (xor0633^xor0639^xor0637^xor0635); // MakeXorFrom
assign xor0801 = (xor0769^xor0772^xor0770^xor0771); // MakeXorFrom
assign xor0802 = (xor0775^xor0776^xor0773^xor0774); // MakeXorFrom
assign xor0803 = (xor0777^xor0780^xor0778^xor0779); // MakeXorFrom
assign xor0804 = (xor0782^xor0783^xor0784^xor0781); // MakeXorFrom
assign xor0805 = (xor0787^xor0788^xor0785^xor0786); // MakeXorFrom
assign xor0806 = (xor0790^xor0791^xor0789^xor0792); // MakeXorFrom
assign xor0807 = (xor0795^xor0796^xor0793^xor0794); // MakeXorFrom
assign xor0808 = (xor0800^xor0797^xor0798^xor0799); // MakeXorFrom
assign xor0809 = (xor0803^xor0804^xor0801^xor0802); // MakeXorFrom
assign xor0810 = (xor0808^xor0805^xor0806^xor0807); // MakeXorFrom
assign xor0811 = (xor0810^xor0809); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 4
assign xor0812 = (xor0006^xor0014^xor0004^xor0012); // MakeXorFrom
assign xor0813 = (xor0030^xor0020^xor0028^xor0022); // MakeXorFrom
assign xor0814 = (xor0038^xor0046^xor0036^xor0044); // MakeXorFrom
assign xor0815 = (xor0054^xor0062^xor0052^xor0060); // MakeXorFrom
assign xor0816 = (xor0076^xor0078^xor0070^xor0068); // MakeXorFrom
assign xor0817 = (xor0086^xor0094^xor0084^xor0092); // MakeXorFrom
assign xor0818 = (xor0110^xor0100^xor0108^xor0102); // MakeXorFrom
assign xor0819 = (xor0118^xor0126^xor0116^xor0124); // MakeXorFrom
assign xor0820 = (xor0134^xor0142^xor0132^xor0140); // MakeXorFrom
assign xor0821 = (xor0156^xor0150^xor0158^xor0148); // MakeXorFrom
assign xor0822 = (xor0166^xor0174^xor0164^xor0172); // MakeXorFrom
assign xor0823 = (xor0182^xor0190^xor0180^xor0188); // MakeXorFrom
assign xor0824 = (xor0204^xor0198^xor0206^xor0196); // MakeXorFrom
assign xor0825 = (xor0222^xor0212^xor0220^xor0214); // MakeXorFrom
assign xor0826 = (xor0230^xor0238^xor0228^xor0236); // MakeXorFrom
assign xor0827 = (xor0246^xor0254^xor0244^xor0252); // MakeXorFrom
assign xor0828 = (xor0514^xor0519^xor0518^xor0515); // MakeXorFrom
assign xor0829 = (xor0522^xor0527^xor0526^xor0523); // MakeXorFrom
assign xor0830 = (xor0530^xor0535^xor0534^xor0531); // MakeXorFrom
assign xor0831 = (xor0539^xor0542^xor0538^xor0543); // MakeXorFrom
assign xor0832 = (xor0550^xor0547^xor0546^xor0551); // MakeXorFrom
assign xor0833 = (xor0558^xor0555^xor0554^xor0559); // MakeXorFrom
assign xor0834 = (xor0567^xor0566^xor0563^xor0562); // MakeXorFrom
assign xor0835 = (xor0570^xor0575^xor0574^xor0571); // MakeXorFrom
assign xor0836 = (xor0578^xor0583^xor0579^xor0582); // MakeXorFrom
assign xor0837 = (xor0586^xor0591^xor0590^xor0587); // MakeXorFrom
assign xor0838 = (xor0598^xor0595^xor0594^xor0599); // MakeXorFrom
assign xor0839 = (xor0606^xor0603^xor0602^xor0607); // MakeXorFrom
assign xor0840 = (xor0614^xor0611^xor0610^xor0615); // MakeXorFrom
assign xor0841 = (xor0623^xor0619^xor0622^xor0618); // MakeXorFrom
assign xor0842 = (xor0626^xor0631^xor0630^xor0627); // MakeXorFrom
assign xor0843 = (xor0634^xor0639^xor0638^xor0635); // MakeXorFrom
assign xor0844 = (xor0815^xor0813^xor0814^xor0812); // MakeXorFrom
assign xor0845 = (xor0818^xor0816^xor0819^xor0817); // MakeXorFrom
assign xor0846 = (xor0823^xor0821^xor0822^xor0820); // MakeXorFrom
assign xor0847 = (xor0825^xor0826^xor0824^xor0827); // MakeXorFrom
assign xor0848 = (xor0828^xor0831^xor0829^xor0830); // MakeXorFrom
assign xor0849 = (xor0835^xor0833^xor0834^xor0832); // MakeXorFrom
assign xor0850 = (xor0836^xor0839^xor0837^xor0838); // MakeXorFrom
assign xor0851 = (xor0843^xor0841^xor0842^xor0840); // MakeXorFrom
assign xor0852 = (xor0846^xor0844^xor0847^xor0845); // MakeXorFrom
assign xor0853 = (xor0851^xor0849^xor0850^xor0848); // MakeXorFrom
assign xor0854 = (xor0853^xor0852); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 5
assign xor0855 = (xor0010^xor0008^xor0014^xor0012); // MakeXorFrom
assign xor0856 = (xor0030^xor0028^xor0026^xor0024); // MakeXorFrom
assign xor0857 = (xor0040^xor0046^xor0044^xor0042); // MakeXorFrom
assign xor0858 = (xor0056^xor0062^xor0060^xor0058); // MakeXorFrom
assign xor0859 = (xor0076^xor0074^xor0072^xor0078); // MakeXorFrom
assign xor0860 = (xor0094^xor0092^xor0090^xor0088); // MakeXorFrom
assign xor0861 = (xor0110^xor0108^xor0106^xor0104); // MakeXorFrom
assign xor0862 = (xor0120^xor0126^xor0124^xor0122); // MakeXorFrom
assign xor0863 = (xor0138^xor0136^xor0142^xor0140); // MakeXorFrom
assign xor0864 = (xor0156^xor0154^xor0152^xor0158); // MakeXorFrom
assign xor0865 = (xor0174^xor0172^xor0170^xor0168); // MakeXorFrom
assign xor0866 = (xor0184^xor0190^xor0188^xor0186); // MakeXorFrom
assign xor0867 = (xor0204^xor0202^xor0200^xor0206); // MakeXorFrom
assign xor0868 = (xor0222^xor0220^xor0218^xor0216); // MakeXorFrom
assign xor0869 = (xor0232^xor0238^xor0236^xor0234); // MakeXorFrom
assign xor0870 = (xor0250^xor0248^xor0254^xor0252); // MakeXorFrom
assign xor0871 = (xor0731^xor0729^xor0727^xor0733); // MakeXorFrom
assign xor0872 = (xor0741^xor0739^xor0737^xor0735); // MakeXorFrom
assign xor0873 = (xor0749^xor0747^xor0745^xor0743); // MakeXorFrom
assign xor0874 = (xor0751^xor0757^xor0755^xor0753); // MakeXorFrom
assign xor0875 = (xor0856^xor0857^xor0858^xor0855); // MakeXorFrom
assign xor0876 = (xor0861^xor0859^xor0862^xor0860); // MakeXorFrom
assign xor0877 = (xor0863^xor0864^xor0865^xor0866); // MakeXorFrom
assign xor0878 = (xor0869^xor0867^xor0870^xor0868); // MakeXorFrom
assign xor0879 = (xor0873^xor0874^xor0871^xor0872); // MakeXorFrom
assign xor0880 = (xor0877^xor0878^xor0875^xor0876); // MakeXorFrom
assign xor0881 = xor0879;
assign xor0882 = (xor0881^xor0880); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 6
assign xor0883 = (xor0020^xor0018^xor0016^xor0022); // MakeXorFrom
assign xor0884 = (xor0048^xor0054^xor0052^xor0050); // MakeXorFrom
assign xor0885 = (xor0086^xor0084^xor0082^xor0080); // MakeXorFrom
assign xor0886 = (xor0118^xor0116^xor0114^xor0112); // MakeXorFrom
assign xor0887 = (xor0146^xor0144^xor0150^xor0148); // MakeXorFrom
assign xor0888 = (xor0176^xor0182^xor0180^xor0178); // MakeXorFrom
assign xor0889 = (xor0212^xor0210^xor0208^xor0214); // MakeXorFrom
assign xor0890 = (xor0240^xor0246^xor0244^xor0242); // MakeXorFrom
assign xor0891 = (xor0521^xor0520^xor0525^xor0524); // MakeXorFrom
assign xor0892 = (xor0537^xor0540^xor0536^xor0541); // MakeXorFrom
assign xor0893 = (xor0552^xor0557^xor0556^xor0553); // MakeXorFrom
assign xor0894 = (xor0568^xor0573^xor0569^xor0572); // MakeXorFrom
assign xor0895 = (xor0588^xor0585^xor0584^xor0589); // MakeXorFrom
assign xor0896 = (xor0605^xor0604^xor0601^xor0600); // MakeXorFrom
assign xor0897 = (xor0616^xor0621^xor0617^xor0620); // MakeXorFrom
assign xor0898 = (xor0633^xor0632^xor0637^xor0636); // MakeXorFrom
assign xor0899 = (xor0835^xor0833^xor0831^xor0829); // MakeXorFrom
assign xor0900 = (xor0843^xor0841^xor0839^xor0837); // MakeXorFrom
assign xor0901 = (xor0856^xor0862^xor0860^xor0858); // MakeXorFrom
assign xor0902 = (xor0864^xor0870^xor0868^xor0866); // MakeXorFrom
assign xor0903 = (xor0884^xor0885^xor0886^xor0883); // MakeXorFrom
assign xor0904 = (xor0889^xor0890^xor0887^xor0888); // MakeXorFrom
assign xor0905 = (xor0894^xor0891^xor0892^xor0893); // MakeXorFrom
assign xor0906 = (xor0897^xor0898^xor0895^xor0896); // MakeXorFrom
assign xor0907 = (xor0899^xor0901^xor0902^xor0900); // MakeXorFrom
assign xor0908 = (xor0905^xor0906^xor0903^xor0904); // MakeXorFrom
assign xor0909 = xor0907;
assign xor0910 = (xor0908^xor0909); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 7
assign xor0911 = (xor0038^xor0036^xor0034^xor0032); // MakeXorFrom
assign xor0912 = (xor0100^xor0098^xor0102^xor0096); // MakeXorFrom
assign xor0913 = (xor0166^xor0164^xor0162^xor0160); // MakeXorFrom
assign xor0914 = (xor0230^xor0228^xor0226^xor0224); // MakeXorFrom
assign xor0915 = (xor0529^xor0532^xor0528^xor0533); // MakeXorFrom
assign xor0916 = (xor0560^xor0565^xor0564^xor0561); // MakeXorFrom
assign xor0917 = (xor0596^xor0593^xor0592^xor0597); // MakeXorFrom
assign xor0918 = (xor0624^xor0629^xor0628^xor0625); // MakeXorFrom
assign xor0919 = (xor0835^xor0834^xor0831^xor0830); // MakeXorFrom
assign xor0920 = (xor0843^xor0839^xor0842^xor0838); // MakeXorFrom
assign xor0921 = (xor0861^xor0862^xor0857^xor0858); // MakeXorFrom
assign xor0922 = (xor0869^xor0870^xor0865^xor0866); // MakeXorFrom
assign xor0923 = (xor0884^xor0890^xor0888^xor0886); // MakeXorFrom
assign xor0924 = (xor0894^xor0892^xor0898^xor0896); // MakeXorFrom
assign xor0925 = (xor0913^xor0914^xor0911^xor0912); // MakeXorFrom
assign xor0926 = (xor0915^xor0916^xor0917^xor0918); // MakeXorFrom
assign xor0927 = (xor0921^xor0922^xor0919^xor0920); // MakeXorFrom
assign xor0928 = (xor0923^xor0924); // MakeXorFrom
assign xor0929 = (xor0926^xor0927^xor0928^xor0925); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 8
assign xor0930 = (xor0066^xor0064^xor0070^xor0068); // MakeXorFrom
assign xor0931 = (xor0194^xor0192^xor0198^xor0196); // MakeXorFrom
assign xor0932 = (xor0548^xor0545^xor0544^xor0549); // MakeXorFrom
assign xor0933 = (xor0613^xor0609^xor0612^xor0608); // MakeXorFrom
assign xor0934 = (xor0851^xor0849^xor0878^xor0876); // MakeXorFrom
assign xor0935 = (xor0889^xor0890^xor0885^xor0886); // MakeXorFrom
assign xor0936 = (xor0894^xor0897^xor0898^xor0893); // MakeXorFrom
assign xor0937 = (xor0916^xor0914^xor0912^xor0918); // MakeXorFrom
assign xor0938 = (xor0933^xor0931^xor0932^xor0930); // MakeXorFrom
assign xor0939 = (xor0936^xor0934^xor0937^xor0935); // MakeXorFrom
assign xor0940 = (xor0939^xor0938); // MakeXorFrom
// BuildXorTrees, ParityBits, i = 9
assign xor0941 = (xor0128^xor0134^xor0132^xor0130); // MakeXorFrom
assign xor0942 = (xor0580^xor0577^xor0576^xor0581); // MakeXorFrom
assign xor0943 = (xor0836^xor0841^xor0837^xor0840); // MakeXorFrom
assign xor0944 = (xor0863^xor0864^xor0867^xor0868); // MakeXorFrom
assign xor0945 = (xor0913^xor0906^xor0914^xor0904); // MakeXorFrom
assign xor0946 = (xor0922^xor0920^xor0917^xor0918); // MakeXorFrom
assign xor0947 = (xor0933^xor0931); // MakeXorFrom
assign xor0948 = (xor0943^xor0944^xor0941^xor0942); // MakeXorFrom
assign xor0949 = (xor0946^xor0947^xor0945); // MakeXorFrom
assign xor0950 = (xor0949^xor0948); // MakeXorFrom
// BuildXorTrees, BuildCheckBit
// BuildCheckBit: building inverse max-parity tree
assign xor0951 = (xor0002^xor0000^xor0006^xor0004); // MakeXorFrom
assign xor0952 = (xor0512^xor0517^xor0516^xor0513); // MakeXorFrom
assign xor0953 = (xor0828^xor0833^xor0832^xor0829); // MakeXorFrom
assign xor0954 = (xor0856^xor0859^xor0860^xor0855); // MakeXorFrom
assign xor0955 = (xor0905^xor0903^xor0911^xor0912); // MakeXorFrom
assign xor0956 = (xor0915^xor0916^xor0921^xor0919); // MakeXorFrom
assign xor0957 = (xor0932^xor0930); // MakeXorFrom
assign xor0958 = (xor0953^xor0954^xor0951^xor0952); // MakeXorFrom
assign xor0959 = (xor0957^xor0955^xor0956); // MakeXorFrom
assign xor0960 = (xor0959^xor0958); // MakeXorFrom
// BuildCheckBit: building check-bit tree
assign xor0961 = (input_data[0009]^input_data[0005]^input_data[0006]^input_data[0003]); // EmitInputXorGate
assign xor0962 = (input_data[0015]^input_data[0017]^input_data[0010]^input_data[0012]); // EmitInputXorGate
assign xor0963 = (input_data[0018]^input_data[0024]^input_data[0020]^input_data[0023]); // EmitInputXorGate
assign xor0964 = (input_data[0027]^input_data[0030]^input_data[0033]^input_data[0029]); // EmitInputXorGate
assign xor0965 = (input_data[0040]^input_data[0034]^input_data[0036]^input_data[0039]); // EmitInputXorGate
assign xor0966 = (input_data[0046]^input_data[0043]^input_data[0048]^input_data[0045]); // EmitInputXorGate
assign xor0967 = (input_data[0051]^input_data[0053]^input_data[0054]^input_data[0057]); // EmitInputXorGate
assign xor0968 = (input_data[0063]^input_data[0058]^input_data[0065]^input_data[0060]); // EmitInputXorGate
assign xor0969 = (input_data[0072]^input_data[0068]^input_data[0071]^input_data[0066]); // EmitInputXorGate
assign xor0970 = (input_data[0078]^input_data[0075]^input_data[0080]^input_data[0077]); // EmitInputXorGate
assign xor0971 = (input_data[0085]^input_data[0086]^input_data[0083]^input_data[0089]); // EmitInputXorGate
assign xor0972 = (input_data[0095]^input_data[0096]^input_data[0090]^input_data[0092]); // EmitInputXorGate
assign xor0973 = (input_data[0105]^input_data[0101]^input_data[0102]^input_data[0099]); // EmitInputXorGate
assign xor0974 = (input_data[0111]^input_data[0106]^input_data[0113]^input_data[0108]); // EmitInputXorGate
assign xor0975 = (input_data[0114]^input_data[0116]^input_data[0120]^input_data[0119]); // EmitInputXorGate
assign xor0976 = (input_data[0126]^input_data[0123]^input_data[0129]^input_data[0125]); // EmitInputXorGate
assign xor0977 = (input_data[0130]^input_data[0132]^input_data[0135]^input_data[0136]); // EmitInputXorGate
assign xor0978 = (input_data[0139]^input_data[0144]^input_data[0141]^input_data[0142]); // EmitInputXorGate
assign xor0979 = (input_data[0149]^input_data[0147]^input_data[0150]^input_data[0153]); // EmitInputXorGate
assign xor0980 = (input_data[0159]^input_data[0154]^input_data[0160]^input_data[0156]); // EmitInputXorGate
assign xor0981 = (input_data[0169]^input_data[0165]^input_data[0166]^input_data[0163]); // EmitInputXorGate
assign xor0982 = (input_data[0175]^input_data[0177]^input_data[0170]^input_data[0172]); // EmitInputXorGate
assign xor0983 = (input_data[0180]^input_data[0183]^input_data[0184]^input_data[0178]); // EmitInputXorGate
assign xor0984 = (input_data[0187]^input_data[0190]^input_data[0192]^input_data[0189]); // EmitInputXorGate
assign xor0985 = (input_data[0201]^input_data[0198]^input_data[0195]^input_data[0197]); // EmitInputXorGate
assign xor0986 = (input_data[0204]^input_data[0207]^input_data[0202]^input_data[0209]); // EmitInputXorGate
assign xor0987 = (input_data[0215]^input_data[0216]^input_data[0210]^input_data[0212]); // EmitInputXorGate
assign xor0988 = (input_data[0221]^input_data[0222]^input_data[0219]^input_data[0225]); // EmitInputXorGate
assign xor0989 = (input_data[0231]^input_data[0226]^input_data[0232]^input_data[0228]); // EmitInputXorGate
assign xor0990 = (input_data[0238]^input_data[0235]^input_data[0240]^input_data[0237]); // EmitInputXorGate
assign xor0991 = (input_data[0249]^input_data[0245]^input_data[0246]^input_data[0243]); // EmitInputXorGate
assign xor0992 = (input_data[0255]^input_data[0257]^input_data[0250]^input_data[0252]); // EmitInputXorGate
assign xor0993 = (input_data[0258]^input_data[0264]^input_data[0260]^input_data[0263]); // EmitInputXorGate
assign xor0994 = (input_data[0269]^input_data[0267]^input_data[0270]^input_data[0272]); // EmitInputXorGate
assign xor0995 = (input_data[0278]^input_data[0281]^input_data[0275]^input_data[0277]); // EmitInputXorGate
assign xor0996 = (input_data[0284]^input_data[0287]^input_data[0282]^input_data[0288]); // EmitInputXorGate
assign xor0997 = (input_data[0291]^input_data[0293]^input_data[0294]^input_data[0297]); // EmitInputXorGate
assign xor0998 = (input_data[0300]^input_data[0303]^input_data[0298]^input_data[0305]); // EmitInputXorGate
assign xor0999 = (input_data[0312]^input_data[0308]^input_data[0311]^input_data[0306]); // EmitInputXorGate
assign xor1000 = (input_data[0318]^input_data[0315]^input_data[0317]^input_data[0320]); // EmitInputXorGate
assign xor1001 = (input_data[0329]^input_data[0325]^input_data[0326]^input_data[0323]); // EmitInputXorGate
assign xor1002 = (input_data[0335]^input_data[0337]^input_data[0330]^input_data[0332]); // EmitInputXorGate
assign xor1003 = (input_data[0338]^input_data[0344]^input_data[0340]^input_data[0343]); // EmitInputXorGate
assign xor1004 = (input_data[0347]^input_data[0350]^input_data[0353]^input_data[0349]); // EmitInputXorGate
assign xor1005 = (input_data[0354]^input_data[0356]^input_data[0360]^input_data[0359]); // EmitInputXorGate
assign xor1006 = (input_data[0365]^input_data[0366]^input_data[0363]^input_data[0368]); // EmitInputXorGate
assign xor1007 = (input_data[0377]^input_data[0371]^input_data[0373]^input_data[0374]); // EmitInputXorGate
assign xor1008 = (input_data[0383]^input_data[0384]^input_data[0378]^input_data[0380]); // EmitInputXorGate
assign xor1009 = (input_data[0389]^input_data[0387]^input_data[0390]^input_data[0393]); // EmitInputXorGate
assign xor1010 = (input_data[0401]^input_data[0399]^input_data[0394]^input_data[0396]); // EmitInputXorGate
assign xor1011 = (input_data[0404]^input_data[0407]^input_data[0402]^input_data[0408]); // EmitInputXorGate
assign xor1012 = (input_data[0417]^input_data[0411]^input_data[0413]^input_data[0414]); // EmitInputXorGate
assign xor1013 = (input_data[0420]^input_data[0423]^input_data[0418]^input_data[0424]); // EmitInputXorGate
assign xor1014 = (input_data[0430]^input_data[0432]^input_data[0429]^input_data[0427]); // EmitInputXorGate
assign xor1015 = (input_data[0438]^input_data[0435]^input_data[0441]^input_data[0437]); // EmitInputXorGate
assign xor1016 = (input_data[0449]^input_data[0444]^input_data[0447]^input_data[0442]); // EmitInputXorGate
assign xor1017 = (input_data[0455]^input_data[0456]^input_data[0450]^input_data[0452]); // EmitInputXorGate
assign xor1018 = (input_data[0459]^input_data[0464]^input_data[0461]^input_data[0462]); // EmitInputXorGate
assign xor1019 = (input_data[0467]^input_data[0470]^input_data[0473]^input_data[0469]); // EmitInputXorGate
assign xor1020 = (input_data[0480]^input_data[0474]^input_data[0476]^input_data[0479]); // EmitInputXorGate
assign xor1021 = (input_data[0486]^input_data[0483]^input_data[0489]^input_data[0485]); // EmitInputXorGate
assign xor1022 = (input_data[0490]^input_data[0492]^input_data[0495]^input_data[0497]); // EmitInputXorGate
assign xor1023 = (input_data[0500]^input_data[0503]^input_data[0498]^input_data[0504]); // EmitInputXorGate
assign xor1024 = (input_data[0509]^input_data[0507]^input_data[0510]^input_data[0513]); // EmitInputXorGate
assign xor1025 = (input_data[0519]^input_data[0514]^input_data[0516]^input_data[0520]); // EmitInputXorGate
assign xor1026 = (input_data[0528]^input_data[0525]^input_data[0526]^input_data[0523]); // EmitInputXorGate
assign xor1027 = (input_data[0534]^input_data[0537]^input_data[0531]^input_data[0533]); // EmitInputXorGate
assign xor1028 = (input_data[0538]^input_data[0544]^input_data[0540]^input_data[0543]); // EmitInputXorGate
assign xor1029 = (input_data[0547]^input_data[0550]^input_data[0553]^input_data[0549]); // EmitInputXorGate
assign xor1030 = (input_data[0554]^input_data[0561]^input_data[0556]^input_data[0559]); // EmitInputXorGate
assign xor1031 = (input_data[0567]^input_data[0562]^input_data[0568]^input_data[0564]); // EmitInputXorGate
assign xor1032 = (input_data[0571]^input_data[0573]^input_data[0574]^input_data[0576]); // EmitInputXorGate
assign xor1033 = (input_data[0585]^input_data[0579]^input_data[0581]^input_data[0582]); // EmitInputXorGate
assign xor1034 = (input_data[0588]^input_data[0591]^input_data[0586]^input_data[0593]); // EmitInputXorGate
assign xor1035 = (input_data[0600]^input_data[0599]^input_data[0594]^input_data[0596]); // EmitInputXorGate
assign xor1036 = (input_data[0603]^input_data[0609]^input_data[0605]^input_data[0606]); // EmitInputXorGate
assign xor1037 = (input_data[0612]^input_data[0615]^input_data[0616]^input_data[0610]); // EmitInputXorGate
assign xor1038 = (input_data[0619]^input_data[0624]^input_data[0621]^input_data[0622]); // EmitInputXorGate
assign xor1039 = (input_data[0629]^input_data[0627]^input_data[0630]^input_data[0633]); // EmitInputXorGate
assign xor1040 = (input_data[0639]^input_data[0634]^input_data[0640]^input_data[0636]); // EmitInputXorGate
assign xor1041 = (input_data[0645]^input_data[0646]^input_data[0643]^input_data[0649]); // EmitInputXorGate
assign xor1042 = (input_data[0655]^input_data[0657]^input_data[0650]^input_data[0652]); // EmitInputXorGate
assign xor1043 = (input_data[0664]^input_data[0660]^input_data[0663]^input_data[0658]); // EmitInputXorGate
assign xor1044 = (input_data[0667]^input_data[0670]^input_data[0673]^input_data[0669]); // EmitInputXorGate
assign xor1045 = (input_data[0676]^input_data[0679]^input_data[0674]^input_data[0680]); // EmitInputXorGate
assign xor1046 = (input_data[0688]^input_data[0685]^input_data[0686]^input_data[0683]); // EmitInputXorGate
assign xor1047 = (input_data[0694]^input_data[0697]^input_data[0691]^input_data[0693]); // EmitInputXorGate
assign xor1048 = (input_data[0698]^input_data[0705]^input_data[0700]^input_data[0703]); // EmitInputXorGate
assign xor1049 = (input_data[0708]^input_data[0711]^input_data[0706]^input_data[0712]); // EmitInputXorGate
assign xor1050 = (input_data[0718]^input_data[0715]^input_data[0717]^input_data[0720]); // EmitInputXorGate
assign xor1051 = (input_data[0725]^input_data[0726]^input_data[0723]^input_data[0729]); // EmitInputXorGate
assign xor1052 = (input_data[0735]^input_data[0736]^input_data[0730]^input_data[0732]); // EmitInputXorGate
assign xor1053 = (input_data[0741]^input_data[0742]^input_data[0745]^input_data[0739]); // EmitInputXorGate
assign xor1054 = (input_data[0753]^input_data[0748]^input_data[0751]^input_data[0746]); // EmitInputXorGate
assign xor1055 = (input_data[0759]^input_data[0754]^input_data[0760]^input_data[0756]); // EmitInputXorGate
assign xor1056 = (input_data[0768]^input_data[0765]^input_data[0766]^input_data[0763]); // EmitInputXorGate
assign xor1057 = (input_data[0774]^input_data[0777]^input_data[0771]^input_data[0773]); // EmitInputXorGate
assign xor1058 = (input_data[0785]^input_data[0778]^input_data[0780]^input_data[0783]); // EmitInputXorGate
assign xor1059 = (input_data[0788]^input_data[0791]^input_data[0786]^input_data[0792]); // EmitInputXorGate
assign xor1060 = (input_data[0795]^input_data[0797]^input_data[0801]^input_data[0798]); // EmitInputXorGate
assign xor1061 = (input_data[0802]^input_data[0808]^input_data[0804]^input_data[0807]); // EmitInputXorGate
assign xor1062 = (input_data[0814]^input_data[0816]^input_data[0811]^input_data[0813]); // EmitInputXorGate
assign xor1063 = (input_data[0819]^input_data[0825]^input_data[0821]^input_data[0822]); // EmitInputXorGate
assign xor1064 = (input_data[0828]^input_data[0831]^input_data[0826]^input_data[0833]); // EmitInputXorGate
assign xor1065 = (input_data[0839]^input_data[0834]^input_data[0840]^input_data[0836]); // EmitInputXorGate
assign xor1066 = (input_data[0845]^input_data[0846]^input_data[0843]^input_data[0848]); // EmitInputXorGate
assign xor1067 = (input_data[0857]^input_data[0851]^input_data[0853]^input_data[0854]); // EmitInputXorGate
assign xor1068 = (input_data[0860]^input_data[0863]^input_data[0858]^input_data[0864]); // EmitInputXorGate
assign xor1069 = (input_data[0870]^input_data[0873]^input_data[0869]^input_data[0867]); // EmitInputXorGate
assign xor1070 = (input_data[0879]^input_data[0881]^input_data[0874]^input_data[0876]); // EmitInputXorGate
assign xor1071 = (input_data[0888]^input_data[0884]^input_data[0887]^input_data[0882]); // EmitInputXorGate
assign xor1072 = (input_data[0894]^input_data[0897]^input_data[0891]^input_data[0893]); // EmitInputXorGate
assign xor1073 = (input_data[0898]^input_data[0904]^input_data[0900]^input_data[0903]); // EmitInputXorGate
assign xor1074 = (input_data[0907]^input_data[0910]^input_data[0912]^input_data[0909]); // EmitInputXorGate
assign xor1075 = (input_data[0915]^input_data[0917]^input_data[0921]^input_data[0918]); // EmitInputXorGate
assign xor1076 = (input_data[0924]^input_data[0927]^input_data[0922]^input_data[0928]); // EmitInputXorGate
assign xor1077 = (input_data[0934]^input_data[0937]^input_data[0931]^input_data[0933]); // EmitInputXorGate
assign xor1078 = (input_data[0943]^input_data[0945]^input_data[0938]^input_data[0940]); // EmitInputXorGate
assign xor1079 = (input_data[0952]^input_data[0948]^input_data[0951]^input_data[0946]); // EmitInputXorGate
assign xor1080 = (input_data[0958]^input_data[0955]^input_data[0957]^input_data[0960]); // EmitInputXorGate
assign xor1081 = (input_data[0969]^input_data[0965]^input_data[0966]^input_data[0963]); // EmitInputXorGate
assign xor1082 = (input_data[0975]^input_data[0977]^input_data[0970]^input_data[0972]); // EmitInputXorGate
assign xor1083 = (input_data[0978]^input_data[0984]^input_data[0980]^input_data[0983]); // EmitInputXorGate
assign xor1084 = (input_data[0987]^input_data[0990]^input_data[0993]^input_data[0989]); // EmitInputXorGate
assign xor1085 = (input_data[0994]^input_data[0996]^input_data[1000]^input_data[0999]); // EmitInputXorGate
assign xor1086 = (input_data[1008]^input_data[1005]^input_data[1006]^input_data[1003]); // EmitInputXorGate
assign xor1087 = (input_data[1014]^input_data[1017]^input_data[1011]^input_data[1013]); // EmitInputXorGate
assign xor1088 = (input_data[1020]^input_data[1023]^input_data[1018]); // EmitInputXorGate
assign xor1089 = (xor0964^xor0961^xor0962^xor0963); // MakeXorFrom
assign xor1090 = (xor0967^xor0968^xor0965^xor0966); // MakeXorFrom
assign xor1091 = (xor0971^xor0972^xor0969^xor0970); // MakeXorFrom
assign xor1092 = (xor0974^xor0975^xor0976^xor0973); // MakeXorFrom
assign xor1093 = (xor0979^xor0977^xor0980^xor0978); // MakeXorFrom
assign xor1094 = (xor0981^xor0982^xor0983^xor0984); // MakeXorFrom
assign xor1095 = (xor0987^xor0988^xor0985^xor0986); // MakeXorFrom
assign xor1096 = (xor0991^xor0992^xor0989^xor0990); // MakeXorFrom
assign xor1097 = (xor0995^xor0996^xor0993^xor0994); // MakeXorFrom
assign xor1098 = (xor0999^xor0997^xor0998^xor1000); // MakeXorFrom
assign xor1099 = (xor1003^xor1004^xor1001^xor1002); // MakeXorFrom
assign xor1100 = (xor1005^xor1006^xor1007^xor1008); // MakeXorFrom
assign xor1101 = (xor1011^xor1012^xor1009^xor1010); // MakeXorFrom
assign xor1102 = (xor1016^xor1013^xor1014^xor1015); // MakeXorFrom
assign xor1103 = (xor1019^xor1020^xor1017^xor1018); // MakeXorFrom
assign xor1104 = (xor1023^xor1024^xor1021^xor1022); // MakeXorFrom
assign xor1105 = (xor1026^xor1027^xor1028^xor1025); // MakeXorFrom
assign xor1106 = (xor1031^xor1032^xor1029^xor1030); // MakeXorFrom
assign xor1107 = (xor1036^xor1033^xor1034^xor1035); // MakeXorFrom
assign xor1108 = (xor1039^xor1040^xor1037^xor1038); // MakeXorFrom
assign xor1109 = (xor1043^xor1044^xor1041^xor1042); // MakeXorFrom
assign xor1110 = (xor1047^xor1048^xor1045^xor1046); // MakeXorFrom
assign xor1111 = (xor1051^xor1052^xor1049^xor1050); // MakeXorFrom
assign xor1112 = (xor1054^xor1055^xor1056^xor1053); // MakeXorFrom
assign xor1113 = (xor1059^xor1057^xor1060^xor1058); // MakeXorFrom
assign xor1114 = (xor1064^xor1061^xor1062^xor1063); // MakeXorFrom
assign xor1115 = (xor1067^xor1068^xor1065^xor1066); // MakeXorFrom
assign xor1116 = (xor1071^xor1072^xor1069^xor1070); // MakeXorFrom
assign xor1117 = (xor1075^xor1076^xor1073^xor1074); // MakeXorFrom
assign xor1118 = (xor1079^xor1077^xor1080^xor1078); // MakeXorFrom
assign xor1119 = (xor1081^xor1082^xor1083^xor1084); // MakeXorFrom
assign xor1120 = (xor1087^xor1088^xor1085^xor1086); // MakeXorFrom
assign xor1121 = (xor1092^xor1089^xor1090^xor1091); // MakeXorFrom
assign xor1122 = (xor1095^xor1096^xor1093^xor1094); // MakeXorFrom
assign xor1123 = (xor1099^xor1097^xor1098^xor1100); // MakeXorFrom
assign xor1124 = (xor1103^xor1104^xor1101^xor1102); // MakeXorFrom
assign xor1125 = (xor1106^xor1107^xor1108^xor1105); // MakeXorFrom
assign xor1126 = (xor1111^xor1109^xor1112^xor1110); // MakeXorFrom
assign xor1127 = (xor1116^xor1113^xor1114^xor1115); // MakeXorFrom
assign xor1128 = (xor1119^xor1120^xor1117^xor1118); // MakeXorFrom
assign xor1129 = (xor1123^xor1124^xor1121^xor1122); // MakeXorFrom
assign xor1130 = (xor1127^xor1128^xor1125^xor1126); // MakeXorFrom
assign xor1131 = (xor1129^xor1130); // MakeXorFrom
assign ecc_parity[-1] = xor1131;
assign ecc_parity[0] = xor0682;
assign ecc_parity[1] = xor0725;
assign ecc_parity[2] = xor0768;
assign ecc_parity[3] = xor0811;
assign ecc_parity[4] = xor0854;
assign ecc_parity[5] = xor0882;
assign ecc_parity[6] = xor0910;
assign ecc_parity[7] = xor0929;
assign ecc_parity[8] = xor0940;
assign ecc_parity[9] = xor0950;
assign input_data[0] = '0;
assign o_chk     [0] = ecc_parity[0-1];
assign input_data[1] = '0;
assign o_chk     [1] = ecc_parity[1-1];
assign input_data[2] = '0;
assign o_chk     [2] = ecc_parity[2-1];
assign input_data[3] = i_data   [0];
assign o_data    [0] = i_data   [0];
assign input_data[4] = '0;
assign o_chk     [3] = ecc_parity[3-1];
assign input_data[5] = i_data   [1];
assign o_data    [1] = i_data   [1];
assign input_data[6] = i_data   [2];
assign o_data    [2] = i_data   [2];
assign input_data[7] = i_data   [3];
assign o_data    [3] = i_data   [3];
assign input_data[8] = '0;
assign o_chk     [4] = ecc_parity[4-1];
assign input_data[9] = i_data   [4];
assign o_data    [4] = i_data   [4];
assign input_data[10] = i_data   [5];
assign o_data    [5] = i_data   [5];
assign input_data[11] = i_data   [6];
assign o_data    [6] = i_data   [6];
assign input_data[12] = i_data   [7];
assign o_data    [7] = i_data   [7];
assign input_data[13] = i_data   [8];
assign o_data    [8] = i_data   [8];
assign input_data[14] = i_data   [9];
assign o_data    [9] = i_data   [9];
assign input_data[15] = i_data   [10];
assign o_data    [10] = i_data   [10];
assign input_data[16] = '0;
assign o_chk     [5] = ecc_parity[5-1];
assign input_data[17] = i_data   [11];
assign o_data    [11] = i_data   [11];
assign input_data[18] = i_data   [12];
assign o_data    [12] = i_data   [12];
assign input_data[19] = i_data   [13];
assign o_data    [13] = i_data   [13];
assign input_data[20] = i_data   [14];
assign o_data    [14] = i_data   [14];
assign input_data[21] = i_data   [15];
assign o_data    [15] = i_data   [15];
assign input_data[22] = i_data   [16];
assign o_data    [16] = i_data   [16];
assign input_data[23] = i_data   [17];
assign o_data    [17] = i_data   [17];
assign input_data[24] = i_data   [18];
assign o_data    [18] = i_data   [18];
assign input_data[25] = i_data   [19];
assign o_data    [19] = i_data   [19];
assign input_data[26] = i_data   [20];
assign o_data    [20] = i_data   [20];
assign input_data[27] = i_data   [21];
assign o_data    [21] = i_data   [21];
assign input_data[28] = i_data   [22];
assign o_data    [22] = i_data   [22];
assign input_data[29] = i_data   [23];
assign o_data    [23] = i_data   [23];
assign input_data[30] = i_data   [24];
assign o_data    [24] = i_data   [24];
assign input_data[31] = i_data   [25];
assign o_data    [25] = i_data   [25];
assign input_data[32] = '0;
assign o_chk     [6] = ecc_parity[6-1];
assign input_data[33] = i_data   [26];
assign o_data    [26] = i_data   [26];
assign input_data[34] = i_data   [27];
assign o_data    [27] = i_data   [27];
assign input_data[35] = i_data   [28];
assign o_data    [28] = i_data   [28];
assign input_data[36] = i_data   [29];
assign o_data    [29] = i_data   [29];
assign input_data[37] = i_data   [30];
assign o_data    [30] = i_data   [30];
assign input_data[38] = i_data   [31];
assign o_data    [31] = i_data   [31];
assign input_data[39] = i_data   [32];
assign o_data    [32] = i_data   [32];
assign input_data[40] = i_data   [33];
assign o_data    [33] = i_data   [33];
assign input_data[41] = i_data   [34];
assign o_data    [34] = i_data   [34];
assign input_data[42] = i_data   [35];
assign o_data    [35] = i_data   [35];
assign input_data[43] = i_data   [36];
assign o_data    [36] = i_data   [36];
assign input_data[44] = i_data   [37];
assign o_data    [37] = i_data   [37];
assign input_data[45] = i_data   [38];
assign o_data    [38] = i_data   [38];
assign input_data[46] = i_data   [39];
assign o_data    [39] = i_data   [39];
assign input_data[47] = i_data   [40];
assign o_data    [40] = i_data   [40];
assign input_data[48] = i_data   [41];
assign o_data    [41] = i_data   [41];
assign input_data[49] = i_data   [42];
assign o_data    [42] = i_data   [42];
assign input_data[50] = i_data   [43];
assign o_data    [43] = i_data   [43];
assign input_data[51] = i_data   [44];
assign o_data    [44] = i_data   [44];
assign input_data[52] = i_data   [45];
assign o_data    [45] = i_data   [45];
assign input_data[53] = i_data   [46];
assign o_data    [46] = i_data   [46];
assign input_data[54] = i_data   [47];
assign o_data    [47] = i_data   [47];
assign input_data[55] = i_data   [48];
assign o_data    [48] = i_data   [48];
assign input_data[56] = i_data   [49];
assign o_data    [49] = i_data   [49];
assign input_data[57] = i_data   [50];
assign o_data    [50] = i_data   [50];
assign input_data[58] = i_data   [51];
assign o_data    [51] = i_data   [51];
assign input_data[59] = i_data   [52];
assign o_data    [52] = i_data   [52];
assign input_data[60] = i_data   [53];
assign o_data    [53] = i_data   [53];
assign input_data[61] = i_data   [54];
assign o_data    [54] = i_data   [54];
assign input_data[62] = i_data   [55];
assign o_data    [55] = i_data   [55];
assign input_data[63] = i_data   [56];
assign o_data    [56] = i_data   [56];
assign input_data[64] = '0;
assign o_chk     [7] = ecc_parity[7-1];
assign input_data[65] = i_data   [57];
assign o_data    [57] = i_data   [57];
assign input_data[66] = i_data   [58];
assign o_data    [58] = i_data   [58];
assign input_data[67] = i_data   [59];
assign o_data    [59] = i_data   [59];
assign input_data[68] = i_data   [60];
assign o_data    [60] = i_data   [60];
assign input_data[69] = i_data   [61];
assign o_data    [61] = i_data   [61];
assign input_data[70] = i_data   [62];
assign o_data    [62] = i_data   [62];
assign input_data[71] = i_data   [63];
assign o_data    [63] = i_data   [63];
assign input_data[72] = i_data   [64];
assign o_data    [64] = i_data   [64];
assign input_data[73] = i_data   [65];
assign o_data    [65] = i_data   [65];
assign input_data[74] = i_data   [66];
assign o_data    [66] = i_data   [66];
assign input_data[75] = i_data   [67];
assign o_data    [67] = i_data   [67];
assign input_data[76] = i_data   [68];
assign o_data    [68] = i_data   [68];
assign input_data[77] = i_data   [69];
assign o_data    [69] = i_data   [69];
assign input_data[78] = i_data   [70];
assign o_data    [70] = i_data   [70];
assign input_data[79] = i_data   [71];
assign o_data    [71] = i_data   [71];
assign input_data[80] = i_data   [72];
assign o_data    [72] = i_data   [72];
assign input_data[81] = i_data   [73];
assign o_data    [73] = i_data   [73];
assign input_data[82] = i_data   [74];
assign o_data    [74] = i_data   [74];
assign input_data[83] = i_data   [75];
assign o_data    [75] = i_data   [75];
assign input_data[84] = i_data   [76];
assign o_data    [76] = i_data   [76];
assign input_data[85] = i_data   [77];
assign o_data    [77] = i_data   [77];
assign input_data[86] = i_data   [78];
assign o_data    [78] = i_data   [78];
assign input_data[87] = i_data   [79];
assign o_data    [79] = i_data   [79];
assign input_data[88] = i_data   [80];
assign o_data    [80] = i_data   [80];
assign input_data[89] = i_data   [81];
assign o_data    [81] = i_data   [81];
assign input_data[90] = i_data   [82];
assign o_data    [82] = i_data   [82];
assign input_data[91] = i_data   [83];
assign o_data    [83] = i_data   [83];
assign input_data[92] = i_data   [84];
assign o_data    [84] = i_data   [84];
assign input_data[93] = i_data   [85];
assign o_data    [85] = i_data   [85];
assign input_data[94] = i_data   [86];
assign o_data    [86] = i_data   [86];
assign input_data[95] = i_data   [87];
assign o_data    [87] = i_data   [87];
assign input_data[96] = i_data   [88];
assign o_data    [88] = i_data   [88];
assign input_data[97] = i_data   [89];
assign o_data    [89] = i_data   [89];
assign input_data[98] = i_data   [90];
assign o_data    [90] = i_data   [90];
assign input_data[99] = i_data   [91];
assign o_data    [91] = i_data   [91];
assign input_data[100] = i_data   [92];
assign o_data    [92] = i_data   [92];
assign input_data[101] = i_data   [93];
assign o_data    [93] = i_data   [93];
assign input_data[102] = i_data   [94];
assign o_data    [94] = i_data   [94];
assign input_data[103] = i_data   [95];
assign o_data    [95] = i_data   [95];
assign input_data[104] = i_data   [96];
assign o_data    [96] = i_data   [96];
assign input_data[105] = i_data   [97];
assign o_data    [97] = i_data   [97];
assign input_data[106] = i_data   [98];
assign o_data    [98] = i_data   [98];
assign input_data[107] = i_data   [99];
assign o_data    [99] = i_data   [99];
assign input_data[108] = i_data   [100];
assign o_data    [100] = i_data   [100];
assign input_data[109] = i_data   [101];
assign o_data    [101] = i_data   [101];
assign input_data[110] = i_data   [102];
assign o_data    [102] = i_data   [102];
assign input_data[111] = i_data   [103];
assign o_data    [103] = i_data   [103];
assign input_data[112] = i_data   [104];
assign o_data    [104] = i_data   [104];
assign input_data[113] = i_data   [105];
assign o_data    [105] = i_data   [105];
assign input_data[114] = i_data   [106];
assign o_data    [106] = i_data   [106];
assign input_data[115] = i_data   [107];
assign o_data    [107] = i_data   [107];
assign input_data[116] = i_data   [108];
assign o_data    [108] = i_data   [108];
assign input_data[117] = i_data   [109];
assign o_data    [109] = i_data   [109];
assign input_data[118] = i_data   [110];
assign o_data    [110] = i_data   [110];
assign input_data[119] = i_data   [111];
assign o_data    [111] = i_data   [111];
assign input_data[120] = i_data   [112];
assign o_data    [112] = i_data   [112];
assign input_data[121] = i_data   [113];
assign o_data    [113] = i_data   [113];
assign input_data[122] = i_data   [114];
assign o_data    [114] = i_data   [114];
assign input_data[123] = i_data   [115];
assign o_data    [115] = i_data   [115];
assign input_data[124] = i_data   [116];
assign o_data    [116] = i_data   [116];
assign input_data[125] = i_data   [117];
assign o_data    [117] = i_data   [117];
assign input_data[126] = i_data   [118];
assign o_data    [118] = i_data   [118];
assign input_data[127] = i_data   [119];
assign o_data    [119] = i_data   [119];
assign input_data[128] = '0;
assign o_chk     [8] = ecc_parity[8-1];
assign input_data[129] = i_data   [120];
assign o_data    [120] = i_data   [120];
assign input_data[130] = i_data   [121];
assign o_data    [121] = i_data   [121];
assign input_data[131] = i_data   [122];
assign o_data    [122] = i_data   [122];
assign input_data[132] = i_data   [123];
assign o_data    [123] = i_data   [123];
assign input_data[133] = i_data   [124];
assign o_data    [124] = i_data   [124];
assign input_data[134] = i_data   [125];
assign o_data    [125] = i_data   [125];
assign input_data[135] = i_data   [126];
assign o_data    [126] = i_data   [126];
assign input_data[136] = i_data   [127];
assign o_data    [127] = i_data   [127];
assign input_data[137] = i_data   [128];
assign o_data    [128] = i_data   [128];
assign input_data[138] = i_data   [129];
assign o_data    [129] = i_data   [129];
assign input_data[139] = i_data   [130];
assign o_data    [130] = i_data   [130];
assign input_data[140] = i_data   [131];
assign o_data    [131] = i_data   [131];
assign input_data[141] = i_data   [132];
assign o_data    [132] = i_data   [132];
assign input_data[142] = i_data   [133];
assign o_data    [133] = i_data   [133];
assign input_data[143] = i_data   [134];
assign o_data    [134] = i_data   [134];
assign input_data[144] = i_data   [135];
assign o_data    [135] = i_data   [135];
assign input_data[145] = i_data   [136];
assign o_data    [136] = i_data   [136];
assign input_data[146] = i_data   [137];
assign o_data    [137] = i_data   [137];
assign input_data[147] = i_data   [138];
assign o_data    [138] = i_data   [138];
assign input_data[148] = i_data   [139];
assign o_data    [139] = i_data   [139];
assign input_data[149] = i_data   [140];
assign o_data    [140] = i_data   [140];
assign input_data[150] = i_data   [141];
assign o_data    [141] = i_data   [141];
assign input_data[151] = i_data   [142];
assign o_data    [142] = i_data   [142];
assign input_data[152] = i_data   [143];
assign o_data    [143] = i_data   [143];
assign input_data[153] = i_data   [144];
assign o_data    [144] = i_data   [144];
assign input_data[154] = i_data   [145];
assign o_data    [145] = i_data   [145];
assign input_data[155] = i_data   [146];
assign o_data    [146] = i_data   [146];
assign input_data[156] = i_data   [147];
assign o_data    [147] = i_data   [147];
assign input_data[157] = i_data   [148];
assign o_data    [148] = i_data   [148];
assign input_data[158] = i_data   [149];
assign o_data    [149] = i_data   [149];
assign input_data[159] = i_data   [150];
assign o_data    [150] = i_data   [150];
assign input_data[160] = i_data   [151];
assign o_data    [151] = i_data   [151];
assign input_data[161] = i_data   [152];
assign o_data    [152] = i_data   [152];
assign input_data[162] = i_data   [153];
assign o_data    [153] = i_data   [153];
assign input_data[163] = i_data   [154];
assign o_data    [154] = i_data   [154];
assign input_data[164] = i_data   [155];
assign o_data    [155] = i_data   [155];
assign input_data[165] = i_data   [156];
assign o_data    [156] = i_data   [156];
assign input_data[166] = i_data   [157];
assign o_data    [157] = i_data   [157];
assign input_data[167] = i_data   [158];
assign o_data    [158] = i_data   [158];
assign input_data[168] = i_data   [159];
assign o_data    [159] = i_data   [159];
assign input_data[169] = i_data   [160];
assign o_data    [160] = i_data   [160];
assign input_data[170] = i_data   [161];
assign o_data    [161] = i_data   [161];
assign input_data[171] = i_data   [162];
assign o_data    [162] = i_data   [162];
assign input_data[172] = i_data   [163];
assign o_data    [163] = i_data   [163];
assign input_data[173] = i_data   [164];
assign o_data    [164] = i_data   [164];
assign input_data[174] = i_data   [165];
assign o_data    [165] = i_data   [165];
assign input_data[175] = i_data   [166];
assign o_data    [166] = i_data   [166];
assign input_data[176] = i_data   [167];
assign o_data    [167] = i_data   [167];
assign input_data[177] = i_data   [168];
assign o_data    [168] = i_data   [168];
assign input_data[178] = i_data   [169];
assign o_data    [169] = i_data   [169];
assign input_data[179] = i_data   [170];
assign o_data    [170] = i_data   [170];
assign input_data[180] = i_data   [171];
assign o_data    [171] = i_data   [171];
assign input_data[181] = i_data   [172];
assign o_data    [172] = i_data   [172];
assign input_data[182] = i_data   [173];
assign o_data    [173] = i_data   [173];
assign input_data[183] = i_data   [174];
assign o_data    [174] = i_data   [174];
assign input_data[184] = i_data   [175];
assign o_data    [175] = i_data   [175];
assign input_data[185] = i_data   [176];
assign o_data    [176] = i_data   [176];
assign input_data[186] = i_data   [177];
assign o_data    [177] = i_data   [177];
assign input_data[187] = i_data   [178];
assign o_data    [178] = i_data   [178];
assign input_data[188] = i_data   [179];
assign o_data    [179] = i_data   [179];
assign input_data[189] = i_data   [180];
assign o_data    [180] = i_data   [180];
assign input_data[190] = i_data   [181];
assign o_data    [181] = i_data   [181];
assign input_data[191] = i_data   [182];
assign o_data    [182] = i_data   [182];
assign input_data[192] = i_data   [183];
assign o_data    [183] = i_data   [183];
assign input_data[193] = i_data   [184];
assign o_data    [184] = i_data   [184];
assign input_data[194] = i_data   [185];
assign o_data    [185] = i_data   [185];
assign input_data[195] = i_data   [186];
assign o_data    [186] = i_data   [186];
assign input_data[196] = i_data   [187];
assign o_data    [187] = i_data   [187];
assign input_data[197] = i_data   [188];
assign o_data    [188] = i_data   [188];
assign input_data[198] = i_data   [189];
assign o_data    [189] = i_data   [189];
assign input_data[199] = i_data   [190];
assign o_data    [190] = i_data   [190];
assign input_data[200] = i_data   [191];
assign o_data    [191] = i_data   [191];
assign input_data[201] = i_data   [192];
assign o_data    [192] = i_data   [192];
assign input_data[202] = i_data   [193];
assign o_data    [193] = i_data   [193];
assign input_data[203] = i_data   [194];
assign o_data    [194] = i_data   [194];
assign input_data[204] = i_data   [195];
assign o_data    [195] = i_data   [195];
assign input_data[205] = i_data   [196];
assign o_data    [196] = i_data   [196];
assign input_data[206] = i_data   [197];
assign o_data    [197] = i_data   [197];
assign input_data[207] = i_data   [198];
assign o_data    [198] = i_data   [198];
assign input_data[208] = i_data   [199];
assign o_data    [199] = i_data   [199];
assign input_data[209] = i_data   [200];
assign o_data    [200] = i_data   [200];
assign input_data[210] = i_data   [201];
assign o_data    [201] = i_data   [201];
assign input_data[211] = i_data   [202];
assign o_data    [202] = i_data   [202];
assign input_data[212] = i_data   [203];
assign o_data    [203] = i_data   [203];
assign input_data[213] = i_data   [204];
assign o_data    [204] = i_data   [204];
assign input_data[214] = i_data   [205];
assign o_data    [205] = i_data   [205];
assign input_data[215] = i_data   [206];
assign o_data    [206] = i_data   [206];
assign input_data[216] = i_data   [207];
assign o_data    [207] = i_data   [207];
assign input_data[217] = i_data   [208];
assign o_data    [208] = i_data   [208];
assign input_data[218] = i_data   [209];
assign o_data    [209] = i_data   [209];
assign input_data[219] = i_data   [210];
assign o_data    [210] = i_data   [210];
assign input_data[220] = i_data   [211];
assign o_data    [211] = i_data   [211];
assign input_data[221] = i_data   [212];
assign o_data    [212] = i_data   [212];
assign input_data[222] = i_data   [213];
assign o_data    [213] = i_data   [213];
assign input_data[223] = i_data   [214];
assign o_data    [214] = i_data   [214];
assign input_data[224] = i_data   [215];
assign o_data    [215] = i_data   [215];
assign input_data[225] = i_data   [216];
assign o_data    [216] = i_data   [216];
assign input_data[226] = i_data   [217];
assign o_data    [217] = i_data   [217];
assign input_data[227] = i_data   [218];
assign o_data    [218] = i_data   [218];
assign input_data[228] = i_data   [219];
assign o_data    [219] = i_data   [219];
assign input_data[229] = i_data   [220];
assign o_data    [220] = i_data   [220];
assign input_data[230] = i_data   [221];
assign o_data    [221] = i_data   [221];
assign input_data[231] = i_data   [222];
assign o_data    [222] = i_data   [222];
assign input_data[232] = i_data   [223];
assign o_data    [223] = i_data   [223];
assign input_data[233] = i_data   [224];
assign o_data    [224] = i_data   [224];
assign input_data[234] = i_data   [225];
assign o_data    [225] = i_data   [225];
assign input_data[235] = i_data   [226];
assign o_data    [226] = i_data   [226];
assign input_data[236] = i_data   [227];
assign o_data    [227] = i_data   [227];
assign input_data[237] = i_data   [228];
assign o_data    [228] = i_data   [228];
assign input_data[238] = i_data   [229];
assign o_data    [229] = i_data   [229];
assign input_data[239] = i_data   [230];
assign o_data    [230] = i_data   [230];
assign input_data[240] = i_data   [231];
assign o_data    [231] = i_data   [231];
assign input_data[241] = i_data   [232];
assign o_data    [232] = i_data   [232];
assign input_data[242] = i_data   [233];
assign o_data    [233] = i_data   [233];
assign input_data[243] = i_data   [234];
assign o_data    [234] = i_data   [234];
assign input_data[244] = i_data   [235];
assign o_data    [235] = i_data   [235];
assign input_data[245] = i_data   [236];
assign o_data    [236] = i_data   [236];
assign input_data[246] = i_data   [237];
assign o_data    [237] = i_data   [237];
assign input_data[247] = i_data   [238];
assign o_data    [238] = i_data   [238];
assign input_data[248] = i_data   [239];
assign o_data    [239] = i_data   [239];
assign input_data[249] = i_data   [240];
assign o_data    [240] = i_data   [240];
assign input_data[250] = i_data   [241];
assign o_data    [241] = i_data   [241];
assign input_data[251] = i_data   [242];
assign o_data    [242] = i_data   [242];
assign input_data[252] = i_data   [243];
assign o_data    [243] = i_data   [243];
assign input_data[253] = i_data   [244];
assign o_data    [244] = i_data   [244];
assign input_data[254] = i_data   [245];
assign o_data    [245] = i_data   [245];
assign input_data[255] = i_data   [246];
assign o_data    [246] = i_data   [246];
assign input_data[256] = '0;
assign o_chk     [9] = ecc_parity[9-1];
assign input_data[257] = i_data   [247];
assign o_data    [247] = i_data   [247];
assign input_data[258] = i_data   [248];
assign o_data    [248] = i_data   [248];
assign input_data[259] = i_data   [249];
assign o_data    [249] = i_data   [249];
assign input_data[260] = i_data   [250];
assign o_data    [250] = i_data   [250];
assign input_data[261] = i_data   [251];
assign o_data    [251] = i_data   [251];
assign input_data[262] = i_data   [252];
assign o_data    [252] = i_data   [252];
assign input_data[263] = i_data   [253];
assign o_data    [253] = i_data   [253];
assign input_data[264] = i_data   [254];
assign o_data    [254] = i_data   [254];
assign input_data[265] = i_data   [255];
assign o_data    [255] = i_data   [255];
assign input_data[266] = i_data   [256];
assign o_data    [256] = i_data   [256];
assign input_data[267] = i_data   [257];
assign o_data    [257] = i_data   [257];
assign input_data[268] = i_data   [258];
assign o_data    [258] = i_data   [258];
assign input_data[269] = i_data   [259];
assign o_data    [259] = i_data   [259];
assign input_data[270] = i_data   [260];
assign o_data    [260] = i_data   [260];
assign input_data[271] = i_data   [261];
assign o_data    [261] = i_data   [261];
assign input_data[272] = i_data   [262];
assign o_data    [262] = i_data   [262];
assign input_data[273] = i_data   [263];
assign o_data    [263] = i_data   [263];
assign input_data[274] = i_data   [264];
assign o_data    [264] = i_data   [264];
assign input_data[275] = i_data   [265];
assign o_data    [265] = i_data   [265];
assign input_data[276] = i_data   [266];
assign o_data    [266] = i_data   [266];
assign input_data[277] = i_data   [267];
assign o_data    [267] = i_data   [267];
assign input_data[278] = i_data   [268];
assign o_data    [268] = i_data   [268];
assign input_data[279] = i_data   [269];
assign o_data    [269] = i_data   [269];
assign input_data[280] = i_data   [270];
assign o_data    [270] = i_data   [270];
assign input_data[281] = i_data   [271];
assign o_data    [271] = i_data   [271];
assign input_data[282] = i_data   [272];
assign o_data    [272] = i_data   [272];
assign input_data[283] = i_data   [273];
assign o_data    [273] = i_data   [273];
assign input_data[284] = i_data   [274];
assign o_data    [274] = i_data   [274];
assign input_data[285] = i_data   [275];
assign o_data    [275] = i_data   [275];
assign input_data[286] = i_data   [276];
assign o_data    [276] = i_data   [276];
assign input_data[287] = i_data   [277];
assign o_data    [277] = i_data   [277];
assign input_data[288] = i_data   [278];
assign o_data    [278] = i_data   [278];
assign input_data[289] = i_data   [279];
assign o_data    [279] = i_data   [279];
assign input_data[290] = i_data   [280];
assign o_data    [280] = i_data   [280];
assign input_data[291] = i_data   [281];
assign o_data    [281] = i_data   [281];
assign input_data[292] = i_data   [282];
assign o_data    [282] = i_data   [282];
assign input_data[293] = i_data   [283];
assign o_data    [283] = i_data   [283];
assign input_data[294] = i_data   [284];
assign o_data    [284] = i_data   [284];
assign input_data[295] = i_data   [285];
assign o_data    [285] = i_data   [285];
assign input_data[296] = i_data   [286];
assign o_data    [286] = i_data   [286];
assign input_data[297] = i_data   [287];
assign o_data    [287] = i_data   [287];
assign input_data[298] = i_data   [288];
assign o_data    [288] = i_data   [288];
assign input_data[299] = i_data   [289];
assign o_data    [289] = i_data   [289];
assign input_data[300] = i_data   [290];
assign o_data    [290] = i_data   [290];
assign input_data[301] = i_data   [291];
assign o_data    [291] = i_data   [291];
assign input_data[302] = i_data   [292];
assign o_data    [292] = i_data   [292];
assign input_data[303] = i_data   [293];
assign o_data    [293] = i_data   [293];
assign input_data[304] = i_data   [294];
assign o_data    [294] = i_data   [294];
assign input_data[305] = i_data   [295];
assign o_data    [295] = i_data   [295];
assign input_data[306] = i_data   [296];
assign o_data    [296] = i_data   [296];
assign input_data[307] = i_data   [297];
assign o_data    [297] = i_data   [297];
assign input_data[308] = i_data   [298];
assign o_data    [298] = i_data   [298];
assign input_data[309] = i_data   [299];
assign o_data    [299] = i_data   [299];
assign input_data[310] = i_data   [300];
assign o_data    [300] = i_data   [300];
assign input_data[311] = i_data   [301];
assign o_data    [301] = i_data   [301];
assign input_data[312] = i_data   [302];
assign o_data    [302] = i_data   [302];
assign input_data[313] = i_data   [303];
assign o_data    [303] = i_data   [303];
assign input_data[314] = i_data   [304];
assign o_data    [304] = i_data   [304];
assign input_data[315] = i_data   [305];
assign o_data    [305] = i_data   [305];
assign input_data[316] = i_data   [306];
assign o_data    [306] = i_data   [306];
assign input_data[317] = i_data   [307];
assign o_data    [307] = i_data   [307];
assign input_data[318] = i_data   [308];
assign o_data    [308] = i_data   [308];
assign input_data[319] = i_data   [309];
assign o_data    [309] = i_data   [309];
assign input_data[320] = i_data   [310];
assign o_data    [310] = i_data   [310];
assign input_data[321] = i_data   [311];
assign o_data    [311] = i_data   [311];
assign input_data[322] = i_data   [312];
assign o_data    [312] = i_data   [312];
assign input_data[323] = i_data   [313];
assign o_data    [313] = i_data   [313];
assign input_data[324] = i_data   [314];
assign o_data    [314] = i_data   [314];
assign input_data[325] = i_data   [315];
assign o_data    [315] = i_data   [315];
assign input_data[326] = i_data   [316];
assign o_data    [316] = i_data   [316];
assign input_data[327] = i_data   [317];
assign o_data    [317] = i_data   [317];
assign input_data[328] = i_data   [318];
assign o_data    [318] = i_data   [318];
assign input_data[329] = i_data   [319];
assign o_data    [319] = i_data   [319];
assign input_data[330] = i_data   [320];
assign o_data    [320] = i_data   [320];
assign input_data[331] = i_data   [321];
assign o_data    [321] = i_data   [321];
assign input_data[332] = i_data   [322];
assign o_data    [322] = i_data   [322];
assign input_data[333] = i_data   [323];
assign o_data    [323] = i_data   [323];
assign input_data[334] = i_data   [324];
assign o_data    [324] = i_data   [324];
assign input_data[335] = i_data   [325];
assign o_data    [325] = i_data   [325];
assign input_data[336] = i_data   [326];
assign o_data    [326] = i_data   [326];
assign input_data[337] = i_data   [327];
assign o_data    [327] = i_data   [327];
assign input_data[338] = i_data   [328];
assign o_data    [328] = i_data   [328];
assign input_data[339] = i_data   [329];
assign o_data    [329] = i_data   [329];
assign input_data[340] = i_data   [330];
assign o_data    [330] = i_data   [330];
assign input_data[341] = i_data   [331];
assign o_data    [331] = i_data   [331];
assign input_data[342] = i_data   [332];
assign o_data    [332] = i_data   [332];
assign input_data[343] = i_data   [333];
assign o_data    [333] = i_data   [333];
assign input_data[344] = i_data   [334];
assign o_data    [334] = i_data   [334];
assign input_data[345] = i_data   [335];
assign o_data    [335] = i_data   [335];
assign input_data[346] = i_data   [336];
assign o_data    [336] = i_data   [336];
assign input_data[347] = i_data   [337];
assign o_data    [337] = i_data   [337];
assign input_data[348] = i_data   [338];
assign o_data    [338] = i_data   [338];
assign input_data[349] = i_data   [339];
assign o_data    [339] = i_data   [339];
assign input_data[350] = i_data   [340];
assign o_data    [340] = i_data   [340];
assign input_data[351] = i_data   [341];
assign o_data    [341] = i_data   [341];
assign input_data[352] = i_data   [342];
assign o_data    [342] = i_data   [342];
assign input_data[353] = i_data   [343];
assign o_data    [343] = i_data   [343];
assign input_data[354] = i_data   [344];
assign o_data    [344] = i_data   [344];
assign input_data[355] = i_data   [345];
assign o_data    [345] = i_data   [345];
assign input_data[356] = i_data   [346];
assign o_data    [346] = i_data   [346];
assign input_data[357] = i_data   [347];
assign o_data    [347] = i_data   [347];
assign input_data[358] = i_data   [348];
assign o_data    [348] = i_data   [348];
assign input_data[359] = i_data   [349];
assign o_data    [349] = i_data   [349];
assign input_data[360] = i_data   [350];
assign o_data    [350] = i_data   [350];
assign input_data[361] = i_data   [351];
assign o_data    [351] = i_data   [351];
assign input_data[362] = i_data   [352];
assign o_data    [352] = i_data   [352];
assign input_data[363] = i_data   [353];
assign o_data    [353] = i_data   [353];
assign input_data[364] = i_data   [354];
assign o_data    [354] = i_data   [354];
assign input_data[365] = i_data   [355];
assign o_data    [355] = i_data   [355];
assign input_data[366] = i_data   [356];
assign o_data    [356] = i_data   [356];
assign input_data[367] = i_data   [357];
assign o_data    [357] = i_data   [357];
assign input_data[368] = i_data   [358];
assign o_data    [358] = i_data   [358];
assign input_data[369] = i_data   [359];
assign o_data    [359] = i_data   [359];
assign input_data[370] = i_data   [360];
assign o_data    [360] = i_data   [360];
assign input_data[371] = i_data   [361];
assign o_data    [361] = i_data   [361];
assign input_data[372] = i_data   [362];
assign o_data    [362] = i_data   [362];
assign input_data[373] = i_data   [363];
assign o_data    [363] = i_data   [363];
assign input_data[374] = i_data   [364];
assign o_data    [364] = i_data   [364];
assign input_data[375] = i_data   [365];
assign o_data    [365] = i_data   [365];
assign input_data[376] = i_data   [366];
assign o_data    [366] = i_data   [366];
assign input_data[377] = i_data   [367];
assign o_data    [367] = i_data   [367];
assign input_data[378] = i_data   [368];
assign o_data    [368] = i_data   [368];
assign input_data[379] = i_data   [369];
assign o_data    [369] = i_data   [369];
assign input_data[380] = i_data   [370];
assign o_data    [370] = i_data   [370];
assign input_data[381] = i_data   [371];
assign o_data    [371] = i_data   [371];
assign input_data[382] = i_data   [372];
assign o_data    [372] = i_data   [372];
assign input_data[383] = i_data   [373];
assign o_data    [373] = i_data   [373];
assign input_data[384] = i_data   [374];
assign o_data    [374] = i_data   [374];
assign input_data[385] = i_data   [375];
assign o_data    [375] = i_data   [375];
assign input_data[386] = i_data   [376];
assign o_data    [376] = i_data   [376];
assign input_data[387] = i_data   [377];
assign o_data    [377] = i_data   [377];
assign input_data[388] = i_data   [378];
assign o_data    [378] = i_data   [378];
assign input_data[389] = i_data   [379];
assign o_data    [379] = i_data   [379];
assign input_data[390] = i_data   [380];
assign o_data    [380] = i_data   [380];
assign input_data[391] = i_data   [381];
assign o_data    [381] = i_data   [381];
assign input_data[392] = i_data   [382];
assign o_data    [382] = i_data   [382];
assign input_data[393] = i_data   [383];
assign o_data    [383] = i_data   [383];
assign input_data[394] = i_data   [384];
assign o_data    [384] = i_data   [384];
assign input_data[395] = i_data   [385];
assign o_data    [385] = i_data   [385];
assign input_data[396] = i_data   [386];
assign o_data    [386] = i_data   [386];
assign input_data[397] = i_data   [387];
assign o_data    [387] = i_data   [387];
assign input_data[398] = i_data   [388];
assign o_data    [388] = i_data   [388];
assign input_data[399] = i_data   [389];
assign o_data    [389] = i_data   [389];
assign input_data[400] = i_data   [390];
assign o_data    [390] = i_data   [390];
assign input_data[401] = i_data   [391];
assign o_data    [391] = i_data   [391];
assign input_data[402] = i_data   [392];
assign o_data    [392] = i_data   [392];
assign input_data[403] = i_data   [393];
assign o_data    [393] = i_data   [393];
assign input_data[404] = i_data   [394];
assign o_data    [394] = i_data   [394];
assign input_data[405] = i_data   [395];
assign o_data    [395] = i_data   [395];
assign input_data[406] = i_data   [396];
assign o_data    [396] = i_data   [396];
assign input_data[407] = i_data   [397];
assign o_data    [397] = i_data   [397];
assign input_data[408] = i_data   [398];
assign o_data    [398] = i_data   [398];
assign input_data[409] = i_data   [399];
assign o_data    [399] = i_data   [399];
assign input_data[410] = i_data   [400];
assign o_data    [400] = i_data   [400];
assign input_data[411] = i_data   [401];
assign o_data    [401] = i_data   [401];
assign input_data[412] = i_data   [402];
assign o_data    [402] = i_data   [402];
assign input_data[413] = i_data   [403];
assign o_data    [403] = i_data   [403];
assign input_data[414] = i_data   [404];
assign o_data    [404] = i_data   [404];
assign input_data[415] = i_data   [405];
assign o_data    [405] = i_data   [405];
assign input_data[416] = i_data   [406];
assign o_data    [406] = i_data   [406];
assign input_data[417] = i_data   [407];
assign o_data    [407] = i_data   [407];
assign input_data[418] = i_data   [408];
assign o_data    [408] = i_data   [408];
assign input_data[419] = i_data   [409];
assign o_data    [409] = i_data   [409];
assign input_data[420] = i_data   [410];
assign o_data    [410] = i_data   [410];
assign input_data[421] = i_data   [411];
assign o_data    [411] = i_data   [411];
assign input_data[422] = i_data   [412];
assign o_data    [412] = i_data   [412];
assign input_data[423] = i_data   [413];
assign o_data    [413] = i_data   [413];
assign input_data[424] = i_data   [414];
assign o_data    [414] = i_data   [414];
assign input_data[425] = i_data   [415];
assign o_data    [415] = i_data   [415];
assign input_data[426] = i_data   [416];
assign o_data    [416] = i_data   [416];
assign input_data[427] = i_data   [417];
assign o_data    [417] = i_data   [417];
assign input_data[428] = i_data   [418];
assign o_data    [418] = i_data   [418];
assign input_data[429] = i_data   [419];
assign o_data    [419] = i_data   [419];
assign input_data[430] = i_data   [420];
assign o_data    [420] = i_data   [420];
assign input_data[431] = i_data   [421];
assign o_data    [421] = i_data   [421];
assign input_data[432] = i_data   [422];
assign o_data    [422] = i_data   [422];
assign input_data[433] = i_data   [423];
assign o_data    [423] = i_data   [423];
assign input_data[434] = i_data   [424];
assign o_data    [424] = i_data   [424];
assign input_data[435] = i_data   [425];
assign o_data    [425] = i_data   [425];
assign input_data[436] = i_data   [426];
assign o_data    [426] = i_data   [426];
assign input_data[437] = i_data   [427];
assign o_data    [427] = i_data   [427];
assign input_data[438] = i_data   [428];
assign o_data    [428] = i_data   [428];
assign input_data[439] = i_data   [429];
assign o_data    [429] = i_data   [429];
assign input_data[440] = i_data   [430];
assign o_data    [430] = i_data   [430];
assign input_data[441] = i_data   [431];
assign o_data    [431] = i_data   [431];
assign input_data[442] = i_data   [432];
assign o_data    [432] = i_data   [432];
assign input_data[443] = i_data   [433];
assign o_data    [433] = i_data   [433];
assign input_data[444] = i_data   [434];
assign o_data    [434] = i_data   [434];
assign input_data[445] = i_data   [435];
assign o_data    [435] = i_data   [435];
assign input_data[446] = i_data   [436];
assign o_data    [436] = i_data   [436];
assign input_data[447] = i_data   [437];
assign o_data    [437] = i_data   [437];
assign input_data[448] = i_data   [438];
assign o_data    [438] = i_data   [438];
assign input_data[449] = i_data   [439];
assign o_data    [439] = i_data   [439];
assign input_data[450] = i_data   [440];
assign o_data    [440] = i_data   [440];
assign input_data[451] = i_data   [441];
assign o_data    [441] = i_data   [441];
assign input_data[452] = i_data   [442];
assign o_data    [442] = i_data   [442];
assign input_data[453] = i_data   [443];
assign o_data    [443] = i_data   [443];
assign input_data[454] = i_data   [444];
assign o_data    [444] = i_data   [444];
assign input_data[455] = i_data   [445];
assign o_data    [445] = i_data   [445];
assign input_data[456] = i_data   [446];
assign o_data    [446] = i_data   [446];
assign input_data[457] = i_data   [447];
assign o_data    [447] = i_data   [447];
assign input_data[458] = i_data   [448];
assign o_data    [448] = i_data   [448];
assign input_data[459] = i_data   [449];
assign o_data    [449] = i_data   [449];
assign input_data[460] = i_data   [450];
assign o_data    [450] = i_data   [450];
assign input_data[461] = i_data   [451];
assign o_data    [451] = i_data   [451];
assign input_data[462] = i_data   [452];
assign o_data    [452] = i_data   [452];
assign input_data[463] = i_data   [453];
assign o_data    [453] = i_data   [453];
assign input_data[464] = i_data   [454];
assign o_data    [454] = i_data   [454];
assign input_data[465] = i_data   [455];
assign o_data    [455] = i_data   [455];
assign input_data[466] = i_data   [456];
assign o_data    [456] = i_data   [456];
assign input_data[467] = i_data   [457];
assign o_data    [457] = i_data   [457];
assign input_data[468] = i_data   [458];
assign o_data    [458] = i_data   [458];
assign input_data[469] = i_data   [459];
assign o_data    [459] = i_data   [459];
assign input_data[470] = i_data   [460];
assign o_data    [460] = i_data   [460];
assign input_data[471] = i_data   [461];
assign o_data    [461] = i_data   [461];
assign input_data[472] = i_data   [462];
assign o_data    [462] = i_data   [462];
assign input_data[473] = i_data   [463];
assign o_data    [463] = i_data   [463];
assign input_data[474] = i_data   [464];
assign o_data    [464] = i_data   [464];
assign input_data[475] = i_data   [465];
assign o_data    [465] = i_data   [465];
assign input_data[476] = i_data   [466];
assign o_data    [466] = i_data   [466];
assign input_data[477] = i_data   [467];
assign o_data    [467] = i_data   [467];
assign input_data[478] = i_data   [468];
assign o_data    [468] = i_data   [468];
assign input_data[479] = i_data   [469];
assign o_data    [469] = i_data   [469];
assign input_data[480] = i_data   [470];
assign o_data    [470] = i_data   [470];
assign input_data[481] = i_data   [471];
assign o_data    [471] = i_data   [471];
assign input_data[482] = i_data   [472];
assign o_data    [472] = i_data   [472];
assign input_data[483] = i_data   [473];
assign o_data    [473] = i_data   [473];
assign input_data[484] = i_data   [474];
assign o_data    [474] = i_data   [474];
assign input_data[485] = i_data   [475];
assign o_data    [475] = i_data   [475];
assign input_data[486] = i_data   [476];
assign o_data    [476] = i_data   [476];
assign input_data[487] = i_data   [477];
assign o_data    [477] = i_data   [477];
assign input_data[488] = i_data   [478];
assign o_data    [478] = i_data   [478];
assign input_data[489] = i_data   [479];
assign o_data    [479] = i_data   [479];
assign input_data[490] = i_data   [480];
assign o_data    [480] = i_data   [480];
assign input_data[491] = i_data   [481];
assign o_data    [481] = i_data   [481];
assign input_data[492] = i_data   [482];
assign o_data    [482] = i_data   [482];
assign input_data[493] = i_data   [483];
assign o_data    [483] = i_data   [483];
assign input_data[494] = i_data   [484];
assign o_data    [484] = i_data   [484];
assign input_data[495] = i_data   [485];
assign o_data    [485] = i_data   [485];
assign input_data[496] = i_data   [486];
assign o_data    [486] = i_data   [486];
assign input_data[497] = i_data   [487];
assign o_data    [487] = i_data   [487];
assign input_data[498] = i_data   [488];
assign o_data    [488] = i_data   [488];
assign input_data[499] = i_data   [489];
assign o_data    [489] = i_data   [489];
assign input_data[500] = i_data   [490];
assign o_data    [490] = i_data   [490];
assign input_data[501] = i_data   [491];
assign o_data    [491] = i_data   [491];
assign input_data[502] = i_data   [492];
assign o_data    [492] = i_data   [492];
assign input_data[503] = i_data   [493];
assign o_data    [493] = i_data   [493];
assign input_data[504] = i_data   [494];
assign o_data    [494] = i_data   [494];
assign input_data[505] = i_data   [495];
assign o_data    [495] = i_data   [495];
assign input_data[506] = i_data   [496];
assign o_data    [496] = i_data   [496];
assign input_data[507] = i_data   [497];
assign o_data    [497] = i_data   [497];
assign input_data[508] = i_data   [498];
assign o_data    [498] = i_data   [498];
assign input_data[509] = i_data   [499];
assign o_data    [499] = i_data   [499];
assign input_data[510] = i_data   [500];
assign o_data    [500] = i_data   [500];
assign input_data[511] = i_data   [501];
assign o_data    [501] = i_data   [501];
assign input_data[512] = '0;
assign o_chk     [10] = ecc_parity[10-1];
assign input_data[513] = i_data   [502];
assign o_data    [502] = i_data   [502];
assign input_data[514] = i_data   [503];
assign o_data    [503] = i_data   [503];
assign input_data[515] = i_data   [504];
assign o_data    [504] = i_data   [504];
assign input_data[516] = i_data   [505];
assign o_data    [505] = i_data   [505];
assign input_data[517] = i_data   [506];
assign o_data    [506] = i_data   [506];
assign input_data[518] = i_data   [507];
assign o_data    [507] = i_data   [507];
assign input_data[519] = i_data   [508];
assign o_data    [508] = i_data   [508];
assign input_data[520] = i_data   [509];
assign o_data    [509] = i_data   [509];
assign input_data[521] = i_data   [510];
assign o_data    [510] = i_data   [510];
assign input_data[522] = i_data   [511];
assign o_data    [511] = i_data   [511];
assign input_data[523] = i_data   [512];
assign o_data    [512] = i_data   [512];
assign input_data[524] = i_data   [513];
assign o_data    [513] = i_data   [513];
assign input_data[525] = i_data   [514];
assign o_data    [514] = i_data   [514];
assign input_data[526] = i_data   [515];
assign o_data    [515] = i_data   [515];
assign input_data[527] = i_data   [516];
assign o_data    [516] = i_data   [516];
assign input_data[528] = i_data   [517];
assign o_data    [517] = i_data   [517];
assign input_data[529] = i_data   [518];
assign o_data    [518] = i_data   [518];
assign input_data[530] = i_data   [519];
assign o_data    [519] = i_data   [519];
assign input_data[531] = i_data   [520];
assign o_data    [520] = i_data   [520];
assign input_data[532] = i_data   [521];
assign o_data    [521] = i_data   [521];
assign input_data[533] = i_data   [522];
assign o_data    [522] = i_data   [522];
assign input_data[534] = i_data   [523];
assign o_data    [523] = i_data   [523];
assign input_data[535] = i_data   [524];
assign o_data    [524] = i_data   [524];
assign input_data[536] = i_data   [525];
assign o_data    [525] = i_data   [525];
assign input_data[537] = i_data   [526];
assign o_data    [526] = i_data   [526];
assign input_data[538] = i_data   [527];
assign o_data    [527] = i_data   [527];
assign input_data[539] = i_data   [528];
assign o_data    [528] = i_data   [528];
assign input_data[540] = i_data   [529];
assign o_data    [529] = i_data   [529];
assign input_data[541] = i_data   [530];
assign o_data    [530] = i_data   [530];
assign input_data[542] = i_data   [531];
assign o_data    [531] = i_data   [531];
assign input_data[543] = i_data   [532];
assign o_data    [532] = i_data   [532];
assign input_data[544] = i_data   [533];
assign o_data    [533] = i_data   [533];
assign input_data[545] = i_data   [534];
assign o_data    [534] = i_data   [534];
assign input_data[546] = i_data   [535];
assign o_data    [535] = i_data   [535];
assign input_data[547] = i_data   [536];
assign o_data    [536] = i_data   [536];
assign input_data[548] = i_data   [537];
assign o_data    [537] = i_data   [537];
assign input_data[549] = i_data   [538];
assign o_data    [538] = i_data   [538];
assign input_data[550] = i_data   [539];
assign o_data    [539] = i_data   [539];
assign input_data[551] = i_data   [540];
assign o_data    [540] = i_data   [540];
assign input_data[552] = i_data   [541];
assign o_data    [541] = i_data   [541];
assign input_data[553] = i_data   [542];
assign o_data    [542] = i_data   [542];
assign input_data[554] = i_data   [543];
assign o_data    [543] = i_data   [543];
assign input_data[555] = i_data   [544];
assign o_data    [544] = i_data   [544];
assign input_data[556] = i_data   [545];
assign o_data    [545] = i_data   [545];
assign input_data[557] = i_data   [546];
assign o_data    [546] = i_data   [546];
assign input_data[558] = i_data   [547];
assign o_data    [547] = i_data   [547];
assign input_data[559] = i_data   [548];
assign o_data    [548] = i_data   [548];
assign input_data[560] = i_data   [549];
assign o_data    [549] = i_data   [549];
assign input_data[561] = i_data   [550];
assign o_data    [550] = i_data   [550];
assign input_data[562] = i_data   [551];
assign o_data    [551] = i_data   [551];
assign input_data[563] = i_data   [552];
assign o_data    [552] = i_data   [552];
assign input_data[564] = i_data   [553];
assign o_data    [553] = i_data   [553];
assign input_data[565] = i_data   [554];
assign o_data    [554] = i_data   [554];
assign input_data[566] = i_data   [555];
assign o_data    [555] = i_data   [555];
assign input_data[567] = i_data   [556];
assign o_data    [556] = i_data   [556];
assign input_data[568] = i_data   [557];
assign o_data    [557] = i_data   [557];
assign input_data[569] = i_data   [558];
assign o_data    [558] = i_data   [558];
assign input_data[570] = i_data   [559];
assign o_data    [559] = i_data   [559];
assign input_data[571] = i_data   [560];
assign o_data    [560] = i_data   [560];
assign input_data[572] = i_data   [561];
assign o_data    [561] = i_data   [561];
assign input_data[573] = i_data   [562];
assign o_data    [562] = i_data   [562];
assign input_data[574] = i_data   [563];
assign o_data    [563] = i_data   [563];
assign input_data[575] = i_data   [564];
assign o_data    [564] = i_data   [564];
assign input_data[576] = i_data   [565];
assign o_data    [565] = i_data   [565];
assign input_data[577] = i_data   [566];
assign o_data    [566] = i_data   [566];
assign input_data[578] = i_data   [567];
assign o_data    [567] = i_data   [567];
assign input_data[579] = i_data   [568];
assign o_data    [568] = i_data   [568];
assign input_data[580] = i_data   [569];
assign o_data    [569] = i_data   [569];
assign input_data[581] = i_data   [570];
assign o_data    [570] = i_data   [570];
assign input_data[582] = i_data   [571];
assign o_data    [571] = i_data   [571];
assign input_data[583] = i_data   [572];
assign o_data    [572] = i_data   [572];
assign input_data[584] = i_data   [573];
assign o_data    [573] = i_data   [573];
assign input_data[585] = i_data   [574];
assign o_data    [574] = i_data   [574];
assign input_data[586] = i_data   [575];
assign o_data    [575] = i_data   [575];
assign input_data[587] = i_data   [576];
assign o_data    [576] = i_data   [576];
assign input_data[588] = i_data   [577];
assign o_data    [577] = i_data   [577];
assign input_data[589] = i_data   [578];
assign o_data    [578] = i_data   [578];
assign input_data[590] = i_data   [579];
assign o_data    [579] = i_data   [579];
assign input_data[591] = i_data   [580];
assign o_data    [580] = i_data   [580];
assign input_data[592] = i_data   [581];
assign o_data    [581] = i_data   [581];
assign input_data[593] = i_data   [582];
assign o_data    [582] = i_data   [582];
assign input_data[594] = i_data   [583];
assign o_data    [583] = i_data   [583];
assign input_data[595] = i_data   [584];
assign o_data    [584] = i_data   [584];
assign input_data[596] = i_data   [585];
assign o_data    [585] = i_data   [585];
assign input_data[597] = i_data   [586];
assign o_data    [586] = i_data   [586];
assign input_data[598] = i_data   [587];
assign o_data    [587] = i_data   [587];
assign input_data[599] = i_data   [588];
assign o_data    [588] = i_data   [588];
assign input_data[600] = i_data   [589];
assign o_data    [589] = i_data   [589];
assign input_data[601] = i_data   [590];
assign o_data    [590] = i_data   [590];
assign input_data[602] = i_data   [591];
assign o_data    [591] = i_data   [591];
assign input_data[603] = i_data   [592];
assign o_data    [592] = i_data   [592];
assign input_data[604] = i_data   [593];
assign o_data    [593] = i_data   [593];
assign input_data[605] = i_data   [594];
assign o_data    [594] = i_data   [594];
assign input_data[606] = i_data   [595];
assign o_data    [595] = i_data   [595];
assign input_data[607] = i_data   [596];
assign o_data    [596] = i_data   [596];
assign input_data[608] = i_data   [597];
assign o_data    [597] = i_data   [597];
assign input_data[609] = i_data   [598];
assign o_data    [598] = i_data   [598];
assign input_data[610] = i_data   [599];
assign o_data    [599] = i_data   [599];
assign input_data[611] = i_data   [600];
assign o_data    [600] = i_data   [600];
assign input_data[612] = i_data   [601];
assign o_data    [601] = i_data   [601];
assign input_data[613] = i_data   [602];
assign o_data    [602] = i_data   [602];
assign input_data[614] = i_data   [603];
assign o_data    [603] = i_data   [603];
assign input_data[615] = i_data   [604];
assign o_data    [604] = i_data   [604];
assign input_data[616] = i_data   [605];
assign o_data    [605] = i_data   [605];
assign input_data[617] = i_data   [606];
assign o_data    [606] = i_data   [606];
assign input_data[618] = i_data   [607];
assign o_data    [607] = i_data   [607];
assign input_data[619] = i_data   [608];
assign o_data    [608] = i_data   [608];
assign input_data[620] = i_data   [609];
assign o_data    [609] = i_data   [609];
assign input_data[621] = i_data   [610];
assign o_data    [610] = i_data   [610];
assign input_data[622] = i_data   [611];
assign o_data    [611] = i_data   [611];
assign input_data[623] = i_data   [612];
assign o_data    [612] = i_data   [612];
assign input_data[624] = i_data   [613];
assign o_data    [613] = i_data   [613];
assign input_data[625] = i_data   [614];
assign o_data    [614] = i_data   [614];
assign input_data[626] = i_data   [615];
assign o_data    [615] = i_data   [615];
assign input_data[627] = i_data   [616];
assign o_data    [616] = i_data   [616];
assign input_data[628] = i_data   [617];
assign o_data    [617] = i_data   [617];
assign input_data[629] = i_data   [618];
assign o_data    [618] = i_data   [618];
assign input_data[630] = i_data   [619];
assign o_data    [619] = i_data   [619];
assign input_data[631] = i_data   [620];
assign o_data    [620] = i_data   [620];
assign input_data[632] = i_data   [621];
assign o_data    [621] = i_data   [621];
assign input_data[633] = i_data   [622];
assign o_data    [622] = i_data   [622];
assign input_data[634] = i_data   [623];
assign o_data    [623] = i_data   [623];
assign input_data[635] = i_data   [624];
assign o_data    [624] = i_data   [624];
assign input_data[636] = i_data   [625];
assign o_data    [625] = i_data   [625];
assign input_data[637] = i_data   [626];
assign o_data    [626] = i_data   [626];
assign input_data[638] = i_data   [627];
assign o_data    [627] = i_data   [627];
assign input_data[639] = i_data   [628];
assign o_data    [628] = i_data   [628];
assign input_data[640] = i_data   [629];
assign o_data    [629] = i_data   [629];
assign input_data[641] = i_data   [630];
assign o_data    [630] = i_data   [630];
assign input_data[642] = i_data   [631];
assign o_data    [631] = i_data   [631];
assign input_data[643] = i_data   [632];
assign o_data    [632] = i_data   [632];
assign input_data[644] = i_data   [633];
assign o_data    [633] = i_data   [633];
assign input_data[645] = i_data   [634];
assign o_data    [634] = i_data   [634];
assign input_data[646] = i_data   [635];
assign o_data    [635] = i_data   [635];
assign input_data[647] = i_data   [636];
assign o_data    [636] = i_data   [636];
assign input_data[648] = i_data   [637];
assign o_data    [637] = i_data   [637];
assign input_data[649] = i_data   [638];
assign o_data    [638] = i_data   [638];
assign input_data[650] = i_data   [639];
assign o_data    [639] = i_data   [639];
assign input_data[651] = i_data   [640];
assign o_data    [640] = i_data   [640];
assign input_data[652] = i_data   [641];
assign o_data    [641] = i_data   [641];
assign input_data[653] = i_data   [642];
assign o_data    [642] = i_data   [642];
assign input_data[654] = i_data   [643];
assign o_data    [643] = i_data   [643];
assign input_data[655] = i_data   [644];
assign o_data    [644] = i_data   [644];
assign input_data[656] = i_data   [645];
assign o_data    [645] = i_data   [645];
assign input_data[657] = i_data   [646];
assign o_data    [646] = i_data   [646];
assign input_data[658] = i_data   [647];
assign o_data    [647] = i_data   [647];
assign input_data[659] = i_data   [648];
assign o_data    [648] = i_data   [648];
assign input_data[660] = i_data   [649];
assign o_data    [649] = i_data   [649];
assign input_data[661] = i_data   [650];
assign o_data    [650] = i_data   [650];
assign input_data[662] = i_data   [651];
assign o_data    [651] = i_data   [651];
assign input_data[663] = i_data   [652];
assign o_data    [652] = i_data   [652];
assign input_data[664] = i_data   [653];
assign o_data    [653] = i_data   [653];
assign input_data[665] = i_data   [654];
assign o_data    [654] = i_data   [654];
assign input_data[666] = i_data   [655];
assign o_data    [655] = i_data   [655];
assign input_data[667] = i_data   [656];
assign o_data    [656] = i_data   [656];
assign input_data[668] = i_data   [657];
assign o_data    [657] = i_data   [657];
assign input_data[669] = i_data   [658];
assign o_data    [658] = i_data   [658];
assign input_data[670] = i_data   [659];
assign o_data    [659] = i_data   [659];
assign input_data[671] = i_data   [660];
assign o_data    [660] = i_data   [660];
assign input_data[672] = i_data   [661];
assign o_data    [661] = i_data   [661];
assign input_data[673] = i_data   [662];
assign o_data    [662] = i_data   [662];
assign input_data[674] = i_data   [663];
assign o_data    [663] = i_data   [663];
assign input_data[675] = i_data   [664];
assign o_data    [664] = i_data   [664];
assign input_data[676] = i_data   [665];
assign o_data    [665] = i_data   [665];
assign input_data[677] = i_data   [666];
assign o_data    [666] = i_data   [666];
assign input_data[678] = i_data   [667];
assign o_data    [667] = i_data   [667];
assign input_data[679] = i_data   [668];
assign o_data    [668] = i_data   [668];
assign input_data[680] = i_data   [669];
assign o_data    [669] = i_data   [669];
assign input_data[681] = i_data   [670];
assign o_data    [670] = i_data   [670];
assign input_data[682] = i_data   [671];
assign o_data    [671] = i_data   [671];
assign input_data[683] = i_data   [672];
assign o_data    [672] = i_data   [672];
assign input_data[684] = i_data   [673];
assign o_data    [673] = i_data   [673];
assign input_data[685] = i_data   [674];
assign o_data    [674] = i_data   [674];
assign input_data[686] = i_data   [675];
assign o_data    [675] = i_data   [675];
assign input_data[687] = i_data   [676];
assign o_data    [676] = i_data   [676];
assign input_data[688] = i_data   [677];
assign o_data    [677] = i_data   [677];
assign input_data[689] = i_data   [678];
assign o_data    [678] = i_data   [678];
assign input_data[690] = i_data   [679];
assign o_data    [679] = i_data   [679];
assign input_data[691] = i_data   [680];
assign o_data    [680] = i_data   [680];
assign input_data[692] = i_data   [681];
assign o_data    [681] = i_data   [681];
assign input_data[693] = i_data   [682];
assign o_data    [682] = i_data   [682];
assign input_data[694] = i_data   [683];
assign o_data    [683] = i_data   [683];
assign input_data[695] = i_data   [684];
assign o_data    [684] = i_data   [684];
assign input_data[696] = i_data   [685];
assign o_data    [685] = i_data   [685];
assign input_data[697] = i_data   [686];
assign o_data    [686] = i_data   [686];
assign input_data[698] = i_data   [687];
assign o_data    [687] = i_data   [687];
assign input_data[699] = i_data   [688];
assign o_data    [688] = i_data   [688];
assign input_data[700] = i_data   [689];
assign o_data    [689] = i_data   [689];
assign input_data[701] = i_data   [690];
assign o_data    [690] = i_data   [690];
assign input_data[702] = i_data   [691];
assign o_data    [691] = i_data   [691];
assign input_data[703] = i_data   [692];
assign o_data    [692] = i_data   [692];
assign input_data[704] = i_data   [693];
assign o_data    [693] = i_data   [693];
assign input_data[705] = i_data   [694];
assign o_data    [694] = i_data   [694];
assign input_data[706] = i_data   [695];
assign o_data    [695] = i_data   [695];
assign input_data[707] = i_data   [696];
assign o_data    [696] = i_data   [696];
assign input_data[708] = i_data   [697];
assign o_data    [697] = i_data   [697];
assign input_data[709] = i_data   [698];
assign o_data    [698] = i_data   [698];
assign input_data[710] = i_data   [699];
assign o_data    [699] = i_data   [699];
assign input_data[711] = i_data   [700];
assign o_data    [700] = i_data   [700];
assign input_data[712] = i_data   [701];
assign o_data    [701] = i_data   [701];
assign input_data[713] = i_data   [702];
assign o_data    [702] = i_data   [702];
assign input_data[714] = i_data   [703];
assign o_data    [703] = i_data   [703];
assign input_data[715] = i_data   [704];
assign o_data    [704] = i_data   [704];
assign input_data[716] = i_data   [705];
assign o_data    [705] = i_data   [705];
assign input_data[717] = i_data   [706];
assign o_data    [706] = i_data   [706];
assign input_data[718] = i_data   [707];
assign o_data    [707] = i_data   [707];
assign input_data[719] = i_data   [708];
assign o_data    [708] = i_data   [708];
assign input_data[720] = i_data   [709];
assign o_data    [709] = i_data   [709];
assign input_data[721] = i_data   [710];
assign o_data    [710] = i_data   [710];
assign input_data[722] = i_data   [711];
assign o_data    [711] = i_data   [711];
assign input_data[723] = i_data   [712];
assign o_data    [712] = i_data   [712];
assign input_data[724] = i_data   [713];
assign o_data    [713] = i_data   [713];
assign input_data[725] = i_data   [714];
assign o_data    [714] = i_data   [714];
assign input_data[726] = i_data   [715];
assign o_data    [715] = i_data   [715];
assign input_data[727] = i_data   [716];
assign o_data    [716] = i_data   [716];
assign input_data[728] = i_data   [717];
assign o_data    [717] = i_data   [717];
assign input_data[729] = i_data   [718];
assign o_data    [718] = i_data   [718];
assign input_data[730] = i_data   [719];
assign o_data    [719] = i_data   [719];
assign input_data[731] = i_data   [720];
assign o_data    [720] = i_data   [720];
assign input_data[732] = i_data   [721];
assign o_data    [721] = i_data   [721];
assign input_data[733] = i_data   [722];
assign o_data    [722] = i_data   [722];
assign input_data[734] = i_data   [723];
assign o_data    [723] = i_data   [723];
assign input_data[735] = i_data   [724];
assign o_data    [724] = i_data   [724];
assign input_data[736] = i_data   [725];
assign o_data    [725] = i_data   [725];
assign input_data[737] = i_data   [726];
assign o_data    [726] = i_data   [726];
assign input_data[738] = i_data   [727];
assign o_data    [727] = i_data   [727];
assign input_data[739] = i_data   [728];
assign o_data    [728] = i_data   [728];
assign input_data[740] = i_data   [729];
assign o_data    [729] = i_data   [729];
assign input_data[741] = i_data   [730];
assign o_data    [730] = i_data   [730];
assign input_data[742] = i_data   [731];
assign o_data    [731] = i_data   [731];
assign input_data[743] = i_data   [732];
assign o_data    [732] = i_data   [732];
assign input_data[744] = i_data   [733];
assign o_data    [733] = i_data   [733];
assign input_data[745] = i_data   [734];
assign o_data    [734] = i_data   [734];
assign input_data[746] = i_data   [735];
assign o_data    [735] = i_data   [735];
assign input_data[747] = i_data   [736];
assign o_data    [736] = i_data   [736];
assign input_data[748] = i_data   [737];
assign o_data    [737] = i_data   [737];
assign input_data[749] = i_data   [738];
assign o_data    [738] = i_data   [738];
assign input_data[750] = i_data   [739];
assign o_data    [739] = i_data   [739];
assign input_data[751] = i_data   [740];
assign o_data    [740] = i_data   [740];
assign input_data[752] = i_data   [741];
assign o_data    [741] = i_data   [741];
assign input_data[753] = i_data   [742];
assign o_data    [742] = i_data   [742];
assign input_data[754] = i_data   [743];
assign o_data    [743] = i_data   [743];
assign input_data[755] = i_data   [744];
assign o_data    [744] = i_data   [744];
assign input_data[756] = i_data   [745];
assign o_data    [745] = i_data   [745];
assign input_data[757] = i_data   [746];
assign o_data    [746] = i_data   [746];
assign input_data[758] = i_data   [747];
assign o_data    [747] = i_data   [747];
assign input_data[759] = i_data   [748];
assign o_data    [748] = i_data   [748];
assign input_data[760] = i_data   [749];
assign o_data    [749] = i_data   [749];
assign input_data[761] = i_data   [750];
assign o_data    [750] = i_data   [750];
assign input_data[762] = i_data   [751];
assign o_data    [751] = i_data   [751];
assign input_data[763] = i_data   [752];
assign o_data    [752] = i_data   [752];
assign input_data[764] = i_data   [753];
assign o_data    [753] = i_data   [753];
assign input_data[765] = i_data   [754];
assign o_data    [754] = i_data   [754];
assign input_data[766] = i_data   [755];
assign o_data    [755] = i_data   [755];
assign input_data[767] = i_data   [756];
assign o_data    [756] = i_data   [756];
assign input_data[768] = i_data   [757];
assign o_data    [757] = i_data   [757];
assign input_data[769] = i_data   [758];
assign o_data    [758] = i_data   [758];
assign input_data[770] = i_data   [759];
assign o_data    [759] = i_data   [759];
assign input_data[771] = i_data   [760];
assign o_data    [760] = i_data   [760];
assign input_data[772] = i_data   [761];
assign o_data    [761] = i_data   [761];
assign input_data[773] = i_data   [762];
assign o_data    [762] = i_data   [762];
assign input_data[774] = i_data   [763];
assign o_data    [763] = i_data   [763];
assign input_data[775] = i_data   [764];
assign o_data    [764] = i_data   [764];
assign input_data[776] = i_data   [765];
assign o_data    [765] = i_data   [765];
assign input_data[777] = i_data   [766];
assign o_data    [766] = i_data   [766];
assign input_data[778] = i_data   [767];
assign o_data    [767] = i_data   [767];
assign input_data[779] = i_data   [768];
assign o_data    [768] = i_data   [768];
assign input_data[780] = i_data   [769];
assign o_data    [769] = i_data   [769];
assign input_data[781] = i_data   [770];
assign o_data    [770] = i_data   [770];
assign input_data[782] = i_data   [771];
assign o_data    [771] = i_data   [771];
assign input_data[783] = i_data   [772];
assign o_data    [772] = i_data   [772];
assign input_data[784] = i_data   [773];
assign o_data    [773] = i_data   [773];
assign input_data[785] = i_data   [774];
assign o_data    [774] = i_data   [774];
assign input_data[786] = i_data   [775];
assign o_data    [775] = i_data   [775];
assign input_data[787] = i_data   [776];
assign o_data    [776] = i_data   [776];
assign input_data[788] = i_data   [777];
assign o_data    [777] = i_data   [777];
assign input_data[789] = i_data   [778];
assign o_data    [778] = i_data   [778];
assign input_data[790] = i_data   [779];
assign o_data    [779] = i_data   [779];
assign input_data[791] = i_data   [780];
assign o_data    [780] = i_data   [780];
assign input_data[792] = i_data   [781];
assign o_data    [781] = i_data   [781];
assign input_data[793] = i_data   [782];
assign o_data    [782] = i_data   [782];
assign input_data[794] = i_data   [783];
assign o_data    [783] = i_data   [783];
assign input_data[795] = i_data   [784];
assign o_data    [784] = i_data   [784];
assign input_data[796] = i_data   [785];
assign o_data    [785] = i_data   [785];
assign input_data[797] = i_data   [786];
assign o_data    [786] = i_data   [786];
assign input_data[798] = i_data   [787];
assign o_data    [787] = i_data   [787];
assign input_data[799] = i_data   [788];
assign o_data    [788] = i_data   [788];
assign input_data[800] = i_data   [789];
assign o_data    [789] = i_data   [789];
assign input_data[801] = i_data   [790];
assign o_data    [790] = i_data   [790];
assign input_data[802] = i_data   [791];
assign o_data    [791] = i_data   [791];
assign input_data[803] = i_data   [792];
assign o_data    [792] = i_data   [792];
assign input_data[804] = i_data   [793];
assign o_data    [793] = i_data   [793];
assign input_data[805] = i_data   [794];
assign o_data    [794] = i_data   [794];
assign input_data[806] = i_data   [795];
assign o_data    [795] = i_data   [795];
assign input_data[807] = i_data   [796];
assign o_data    [796] = i_data   [796];
assign input_data[808] = i_data   [797];
assign o_data    [797] = i_data   [797];
assign input_data[809] = i_data   [798];
assign o_data    [798] = i_data   [798];
assign input_data[810] = i_data   [799];
assign o_data    [799] = i_data   [799];
assign input_data[811] = i_data   [800];
assign o_data    [800] = i_data   [800];
assign input_data[812] = i_data   [801];
assign o_data    [801] = i_data   [801];
assign input_data[813] = i_data   [802];
assign o_data    [802] = i_data   [802];
assign input_data[814] = i_data   [803];
assign o_data    [803] = i_data   [803];
assign input_data[815] = i_data   [804];
assign o_data    [804] = i_data   [804];
assign input_data[816] = i_data   [805];
assign o_data    [805] = i_data   [805];
assign input_data[817] = i_data   [806];
assign o_data    [806] = i_data   [806];
assign input_data[818] = i_data   [807];
assign o_data    [807] = i_data   [807];
assign input_data[819] = i_data   [808];
assign o_data    [808] = i_data   [808];
assign input_data[820] = i_data   [809];
assign o_data    [809] = i_data   [809];
assign input_data[821] = i_data   [810];
assign o_data    [810] = i_data   [810];
assign input_data[822] = i_data   [811];
assign o_data    [811] = i_data   [811];
assign input_data[823] = i_data   [812];
assign o_data    [812] = i_data   [812];
assign input_data[824] = i_data   [813];
assign o_data    [813] = i_data   [813];
assign input_data[825] = i_data   [814];
assign o_data    [814] = i_data   [814];
assign input_data[826] = i_data   [815];
assign o_data    [815] = i_data   [815];
assign input_data[827] = i_data   [816];
assign o_data    [816] = i_data   [816];
assign input_data[828] = i_data   [817];
assign o_data    [817] = i_data   [817];
assign input_data[829] = i_data   [818];
assign o_data    [818] = i_data   [818];
assign input_data[830] = i_data   [819];
assign o_data    [819] = i_data   [819];
assign input_data[831] = i_data   [820];
assign o_data    [820] = i_data   [820];
assign input_data[832] = i_data   [821];
assign o_data    [821] = i_data   [821];
assign input_data[833] = i_data   [822];
assign o_data    [822] = i_data   [822];
assign input_data[834] = i_data   [823];
assign o_data    [823] = i_data   [823];
assign input_data[835] = i_data   [824];
assign o_data    [824] = i_data   [824];
assign input_data[836] = i_data   [825];
assign o_data    [825] = i_data   [825];
assign input_data[837] = i_data   [826];
assign o_data    [826] = i_data   [826];
assign input_data[838] = i_data   [827];
assign o_data    [827] = i_data   [827];
assign input_data[839] = i_data   [828];
assign o_data    [828] = i_data   [828];
assign input_data[840] = i_data   [829];
assign o_data    [829] = i_data   [829];
assign input_data[841] = i_data   [830];
assign o_data    [830] = i_data   [830];
assign input_data[842] = i_data   [831];
assign o_data    [831] = i_data   [831];
assign input_data[843] = i_data   [832];
assign o_data    [832] = i_data   [832];
assign input_data[844] = i_data   [833];
assign o_data    [833] = i_data   [833];
assign input_data[845] = i_data   [834];
assign o_data    [834] = i_data   [834];
assign input_data[846] = i_data   [835];
assign o_data    [835] = i_data   [835];
assign input_data[847] = i_data   [836];
assign o_data    [836] = i_data   [836];
assign input_data[848] = i_data   [837];
assign o_data    [837] = i_data   [837];
assign input_data[849] = i_data   [838];
assign o_data    [838] = i_data   [838];
assign input_data[850] = i_data   [839];
assign o_data    [839] = i_data   [839];
assign input_data[851] = i_data   [840];
assign o_data    [840] = i_data   [840];
assign input_data[852] = i_data   [841];
assign o_data    [841] = i_data   [841];
assign input_data[853] = i_data   [842];
assign o_data    [842] = i_data   [842];
assign input_data[854] = i_data   [843];
assign o_data    [843] = i_data   [843];
assign input_data[855] = i_data   [844];
assign o_data    [844] = i_data   [844];
assign input_data[856] = i_data   [845];
assign o_data    [845] = i_data   [845];
assign input_data[857] = i_data   [846];
assign o_data    [846] = i_data   [846];
assign input_data[858] = i_data   [847];
assign o_data    [847] = i_data   [847];
assign input_data[859] = i_data   [848];
assign o_data    [848] = i_data   [848];
assign input_data[860] = i_data   [849];
assign o_data    [849] = i_data   [849];
assign input_data[861] = i_data   [850];
assign o_data    [850] = i_data   [850];
assign input_data[862] = i_data   [851];
assign o_data    [851] = i_data   [851];
assign input_data[863] = i_data   [852];
assign o_data    [852] = i_data   [852];
assign input_data[864] = i_data   [853];
assign o_data    [853] = i_data   [853];
assign input_data[865] = i_data   [854];
assign o_data    [854] = i_data   [854];
assign input_data[866] = i_data   [855];
assign o_data    [855] = i_data   [855];
assign input_data[867] = i_data   [856];
assign o_data    [856] = i_data   [856];
assign input_data[868] = i_data   [857];
assign o_data    [857] = i_data   [857];
assign input_data[869] = i_data   [858];
assign o_data    [858] = i_data   [858];
assign input_data[870] = i_data   [859];
assign o_data    [859] = i_data   [859];
assign input_data[871] = i_data   [860];
assign o_data    [860] = i_data   [860];
assign input_data[872] = i_data   [861];
assign o_data    [861] = i_data   [861];
assign input_data[873] = i_data   [862];
assign o_data    [862] = i_data   [862];
assign input_data[874] = i_data   [863];
assign o_data    [863] = i_data   [863];
assign input_data[875] = i_data   [864];
assign o_data    [864] = i_data   [864];
assign input_data[876] = i_data   [865];
assign o_data    [865] = i_data   [865];
assign input_data[877] = i_data   [866];
assign o_data    [866] = i_data   [866];
assign input_data[878] = i_data   [867];
assign o_data    [867] = i_data   [867];
assign input_data[879] = i_data   [868];
assign o_data    [868] = i_data   [868];
assign input_data[880] = i_data   [869];
assign o_data    [869] = i_data   [869];
assign input_data[881] = i_data   [870];
assign o_data    [870] = i_data   [870];
assign input_data[882] = i_data   [871];
assign o_data    [871] = i_data   [871];
assign input_data[883] = i_data   [872];
assign o_data    [872] = i_data   [872];
assign input_data[884] = i_data   [873];
assign o_data    [873] = i_data   [873];
assign input_data[885] = i_data   [874];
assign o_data    [874] = i_data   [874];
assign input_data[886] = i_data   [875];
assign o_data    [875] = i_data   [875];
assign input_data[887] = i_data   [876];
assign o_data    [876] = i_data   [876];
assign input_data[888] = i_data   [877];
assign o_data    [877] = i_data   [877];
assign input_data[889] = i_data   [878];
assign o_data    [878] = i_data   [878];
assign input_data[890] = i_data   [879];
assign o_data    [879] = i_data   [879];
assign input_data[891] = i_data   [880];
assign o_data    [880] = i_data   [880];
assign input_data[892] = i_data   [881];
assign o_data    [881] = i_data   [881];
assign input_data[893] = i_data   [882];
assign o_data    [882] = i_data   [882];
assign input_data[894] = i_data   [883];
assign o_data    [883] = i_data   [883];
assign input_data[895] = i_data   [884];
assign o_data    [884] = i_data   [884];
assign input_data[896] = i_data   [885];
assign o_data    [885] = i_data   [885];
assign input_data[897] = i_data   [886];
assign o_data    [886] = i_data   [886];
assign input_data[898] = i_data   [887];
assign o_data    [887] = i_data   [887];
assign input_data[899] = i_data   [888];
assign o_data    [888] = i_data   [888];
assign input_data[900] = i_data   [889];
assign o_data    [889] = i_data   [889];
assign input_data[901] = i_data   [890];
assign o_data    [890] = i_data   [890];
assign input_data[902] = i_data   [891];
assign o_data    [891] = i_data   [891];
assign input_data[903] = i_data   [892];
assign o_data    [892] = i_data   [892];
assign input_data[904] = i_data   [893];
assign o_data    [893] = i_data   [893];
assign input_data[905] = i_data   [894];
assign o_data    [894] = i_data   [894];
assign input_data[906] = i_data   [895];
assign o_data    [895] = i_data   [895];
assign input_data[907] = i_data   [896];
assign o_data    [896] = i_data   [896];
assign input_data[908] = i_data   [897];
assign o_data    [897] = i_data   [897];
assign input_data[909] = i_data   [898];
assign o_data    [898] = i_data   [898];
assign input_data[910] = i_data   [899];
assign o_data    [899] = i_data   [899];
assign input_data[911] = i_data   [900];
assign o_data    [900] = i_data   [900];
assign input_data[912] = i_data   [901];
assign o_data    [901] = i_data   [901];
assign input_data[913] = i_data   [902];
assign o_data    [902] = i_data   [902];
assign input_data[914] = i_data   [903];
assign o_data    [903] = i_data   [903];
assign input_data[915] = i_data   [904];
assign o_data    [904] = i_data   [904];
assign input_data[916] = i_data   [905];
assign o_data    [905] = i_data   [905];
assign input_data[917] = i_data   [906];
assign o_data    [906] = i_data   [906];
assign input_data[918] = i_data   [907];
assign o_data    [907] = i_data   [907];
assign input_data[919] = i_data   [908];
assign o_data    [908] = i_data   [908];
assign input_data[920] = i_data   [909];
assign o_data    [909] = i_data   [909];
assign input_data[921] = i_data   [910];
assign o_data    [910] = i_data   [910];
assign input_data[922] = i_data   [911];
assign o_data    [911] = i_data   [911];
assign input_data[923] = i_data   [912];
assign o_data    [912] = i_data   [912];
assign input_data[924] = i_data   [913];
assign o_data    [913] = i_data   [913];
assign input_data[925] = i_data   [914];
assign o_data    [914] = i_data   [914];
assign input_data[926] = i_data   [915];
assign o_data    [915] = i_data   [915];
assign input_data[927] = i_data   [916];
assign o_data    [916] = i_data   [916];
assign input_data[928] = i_data   [917];
assign o_data    [917] = i_data   [917];
assign input_data[929] = i_data   [918];
assign o_data    [918] = i_data   [918];
assign input_data[930] = i_data   [919];
assign o_data    [919] = i_data   [919];
assign input_data[931] = i_data   [920];
assign o_data    [920] = i_data   [920];
assign input_data[932] = i_data   [921];
assign o_data    [921] = i_data   [921];
assign input_data[933] = i_data   [922];
assign o_data    [922] = i_data   [922];
assign input_data[934] = i_data   [923];
assign o_data    [923] = i_data   [923];
assign input_data[935] = i_data   [924];
assign o_data    [924] = i_data   [924];
assign input_data[936] = i_data   [925];
assign o_data    [925] = i_data   [925];
assign input_data[937] = i_data   [926];
assign o_data    [926] = i_data   [926];
assign input_data[938] = i_data   [927];
assign o_data    [927] = i_data   [927];
assign input_data[939] = i_data   [928];
assign o_data    [928] = i_data   [928];
assign input_data[940] = i_data   [929];
assign o_data    [929] = i_data   [929];
assign input_data[941] = i_data   [930];
assign o_data    [930] = i_data   [930];
assign input_data[942] = i_data   [931];
assign o_data    [931] = i_data   [931];
assign input_data[943] = i_data   [932];
assign o_data    [932] = i_data   [932];
assign input_data[944] = i_data   [933];
assign o_data    [933] = i_data   [933];
assign input_data[945] = i_data   [934];
assign o_data    [934] = i_data   [934];
assign input_data[946] = i_data   [935];
assign o_data    [935] = i_data   [935];
assign input_data[947] = i_data   [936];
assign o_data    [936] = i_data   [936];
assign input_data[948] = i_data   [937];
assign o_data    [937] = i_data   [937];
assign input_data[949] = i_data   [938];
assign o_data    [938] = i_data   [938];
assign input_data[950] = i_data   [939];
assign o_data    [939] = i_data   [939];
assign input_data[951] = i_data   [940];
assign o_data    [940] = i_data   [940];
assign input_data[952] = i_data   [941];
assign o_data    [941] = i_data   [941];
assign input_data[953] = i_data   [942];
assign o_data    [942] = i_data   [942];
assign input_data[954] = i_data   [943];
assign o_data    [943] = i_data   [943];
assign input_data[955] = i_data   [944];
assign o_data    [944] = i_data   [944];
assign input_data[956] = i_data   [945];
assign o_data    [945] = i_data   [945];
assign input_data[957] = i_data   [946];
assign o_data    [946] = i_data   [946];
assign input_data[958] = i_data   [947];
assign o_data    [947] = i_data   [947];
assign input_data[959] = i_data   [948];
assign o_data    [948] = i_data   [948];
assign input_data[960] = i_data   [949];
assign o_data    [949] = i_data   [949];
assign input_data[961] = i_data   [950];
assign o_data    [950] = i_data   [950];
assign input_data[962] = i_data   [951];
assign o_data    [951] = i_data   [951];
assign input_data[963] = i_data   [952];
assign o_data    [952] = i_data   [952];
assign input_data[964] = i_data   [953];
assign o_data    [953] = i_data   [953];
assign input_data[965] = i_data   [954];
assign o_data    [954] = i_data   [954];
assign input_data[966] = i_data   [955];
assign o_data    [955] = i_data   [955];
assign input_data[967] = i_data   [956];
assign o_data    [956] = i_data   [956];
assign input_data[968] = i_data   [957];
assign o_data    [957] = i_data   [957];
assign input_data[969] = i_data   [958];
assign o_data    [958] = i_data   [958];
assign input_data[970] = i_data   [959];
assign o_data    [959] = i_data   [959];
assign input_data[971] = i_data   [960];
assign o_data    [960] = i_data   [960];
assign input_data[972] = i_data   [961];
assign o_data    [961] = i_data   [961];
assign input_data[973] = i_data   [962];
assign o_data    [962] = i_data   [962];
assign input_data[974] = i_data   [963];
assign o_data    [963] = i_data   [963];
assign input_data[975] = i_data   [964];
assign o_data    [964] = i_data   [964];
assign input_data[976] = i_data   [965];
assign o_data    [965] = i_data   [965];
assign input_data[977] = i_data   [966];
assign o_data    [966] = i_data   [966];
assign input_data[978] = i_data   [967];
assign o_data    [967] = i_data   [967];
assign input_data[979] = i_data   [968];
assign o_data    [968] = i_data   [968];
assign input_data[980] = i_data   [969];
assign o_data    [969] = i_data   [969];
assign input_data[981] = i_data   [970];
assign o_data    [970] = i_data   [970];
assign input_data[982] = i_data   [971];
assign o_data    [971] = i_data   [971];
assign input_data[983] = i_data   [972];
assign o_data    [972] = i_data   [972];
assign input_data[984] = i_data   [973];
assign o_data    [973] = i_data   [973];
assign input_data[985] = i_data   [974];
assign o_data    [974] = i_data   [974];
assign input_data[986] = i_data   [975];
assign o_data    [975] = i_data   [975];
assign input_data[987] = i_data   [976];
assign o_data    [976] = i_data   [976];
assign input_data[988] = i_data   [977];
assign o_data    [977] = i_data   [977];
assign input_data[989] = i_data   [978];
assign o_data    [978] = i_data   [978];
assign input_data[990] = i_data   [979];
assign o_data    [979] = i_data   [979];
assign input_data[991] = i_data   [980];
assign o_data    [980] = i_data   [980];
assign input_data[992] = i_data   [981];
assign o_data    [981] = i_data   [981];
assign input_data[993] = i_data   [982];
assign o_data    [982] = i_data   [982];
assign input_data[994] = i_data   [983];
assign o_data    [983] = i_data   [983];
assign input_data[995] = i_data   [984];
assign o_data    [984] = i_data   [984];
assign input_data[996] = i_data   [985];
assign o_data    [985] = i_data   [985];
assign input_data[997] = i_data   [986];
assign o_data    [986] = i_data   [986];
assign input_data[998] = i_data   [987];
assign o_data    [987] = i_data   [987];
assign input_data[999] = i_data   [988];
assign o_data    [988] = i_data   [988];
assign input_data[1000] = i_data   [989];
assign o_data    [989] = i_data   [989];
assign input_data[1001] = i_data   [990];
assign o_data    [990] = i_data   [990];
assign input_data[1002] = i_data   [991];
assign o_data    [991] = i_data   [991];
assign input_data[1003] = i_data   [992];
assign o_data    [992] = i_data   [992];
assign input_data[1004] = i_data   [993];
assign o_data    [993] = i_data   [993];
assign input_data[1005] = i_data   [994];
assign o_data    [994] = i_data   [994];
assign input_data[1006] = i_data   [995];
assign o_data    [995] = i_data   [995];
assign input_data[1007] = i_data   [996];
assign o_data    [996] = i_data   [996];
assign input_data[1008] = i_data   [997];
assign o_data    [997] = i_data   [997];
assign input_data[1009] = i_data   [998];
assign o_data    [998] = i_data   [998];
assign input_data[1010] = i_data   [999];
assign o_data    [999] = i_data   [999];
assign input_data[1011] = i_data   [1000];
assign o_data    [1000] = i_data   [1000];
assign input_data[1012] = i_data   [1001];
assign o_data    [1001] = i_data   [1001];
assign input_data[1013] = i_data   [1002];
assign o_data    [1002] = i_data   [1002];
assign input_data[1014] = i_data   [1003];
assign o_data    [1003] = i_data   [1003];
assign input_data[1015] = i_data   [1004];
assign o_data    [1004] = i_data   [1004];
assign input_data[1016] = i_data   [1005];
assign o_data    [1005] = i_data   [1005];
assign input_data[1017] = i_data   [1006];
assign o_data    [1006] = i_data   [1006];
assign input_data[1018] = i_data   [1007];
assign o_data    [1007] = i_data   [1007];
assign input_data[1019] = i_data   [1008];
assign o_data    [1008] = i_data   [1008];
assign input_data[1020] = i_data   [1009];
assign o_data    [1009] = i_data   [1009];
assign input_data[1021] = i_data   [1010];
assign o_data    [1010] = i_data   [1010];
assign input_data[1022] = i_data   [1011];
assign o_data    [1011] = i_data   [1011];
assign input_data[1023] = i_data   [1012];
assign o_data    [1012] = i_data   [1012];
endmodule
