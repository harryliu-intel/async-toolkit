//                                                                             
// File:       mby_fuse_regs.svh                                               
// Creator:    kmoses1                                                         
// Time:       Sunday Feb 2, 2014 [8:21:51 am]                                 
//                                                                             
// Path:       /tmp/kmoses1/nebulon_run/20231                                  
// Arguments:  /p/com/eda/denali/blueprint/3.7.4/Linux/blueprint -fuse -html -I
//             /p/com/eda/intel/nebulon/2.07p2/include/ -ovm                   
//             mby_fusegen_nebulon.rdl                                         
//                                                                             
// Sources:    /nfs/iil/proj/mpg/kmoses1_wa1/ip_template-nhdk-x0_new/source/rdl/mby_fusegen_nebulon.rdl:5b3e806ef7d09a39437507f3cfbd0ecb
//             /p/com/eda/intel/nebulon/2.07p2/generators/generator_common.pm:4973c402c43f97e18c4aba02585df570
//             /p/com/eda/intel/nebulon/2.07p2/generators/html.pm:a408055bdb3ba8a9656d793e9472104f
//             /p/com/eda/intel/nebulon/2.07p2/generators/ovm.pm:e21c7be001887ff41e17c43b43b1fcdc
//             /p/com/eda/intel/nebulon/2.07p2/include/fuse_udp.rdl:c11891ce81c95bc748bf1f2bdbde2f6f
//             /usr/intel/pkgs/perl/5.8.7/lib64/5.8.7/Digest/base.pm:54bebd0439900c1d44d212cba39747b5
//             /usr/intel/pkgs/perl/5.8.7/lib64/site_perl/Devel/StackTrace.pm:3b99e973435e2dea00aa3a8d6f1b9ddd
//                                                                             
// Blueprint:   3.7.4 (Tue Jun 23 00:17:01 PDT 2009)                           
// Machine:    icsl0104                                                        
// OS:         Linux 2.6.16.60-0.58.1.3835.0.PTF.638363-smp                    
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2014 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY DENALI BLUEPRINT, DO NOT EDIT       
//                                                                             


//RAL code compatible with Saola versions: v20131113 and newer 

`ifndef RAL_MBY_FUSE_FILE
`define RAL_MBY_FUSE_FILE

class mby_fuse_mby_fuse_reg extends sla_ral_reg;

  // --------------------------
  sla_ral_field fuse_1;
  sla_ral_field fuse_2;
  sla_ral_field fuse_3;
  sla_ral_field fuse_4;

  // --------------------------
  `ovm_object_utils(mby_fuse_mby_fuse_reg)

  // --------------------------
  function new(
                string         name = "",
                `ifdef SLA_RAL_COVERAGE
                sla_ral_coverage_t cov_t = COVERAGE_OFF,
                `endif
                int            bus_num=0,
                int            dev_num=0,
                int            func_num=0,
                int            offset=0,
                int            size=0,
                sla_ral_data_t reset_val=0,
                boolean_t      mon_enabled = SLA_FALSE
             );
      super.new();
      set_space_addr("CFG",undef);
      set_space_addr("MEM",undef);
      set_space_addr("IO",undef);
      set_space_addr("MSG",undef);
      set_space_addr("CREG",undef); 
      set_space_addr("LT_MEM",undef);     

      build();

      `ifdef SLA_RAL_COVERAGE
      `CONFIG_RAL_COVERAGE(regname, , )
      if(_coverage_type != COVERAGE_OFF) begin
        if(_sample_type inside {FD_RO_SAMPLE, RO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_WRITE)
        else if(_sample_type inside {FD_WO_SAMPLE, WO_SAMPLE})
        `CREATE_OP_SAMPLE_COV(RAL_READ)
        else
        `CREATE_OP_SAMPLE_COV(RAL_NONE)
        `CREATE_DESIRED_COV
        `CREATE_ACTUAL_COV
      end
      `endif

  endfunction

  `ifdef SLA_RAL_COVERAGE
  `CREATE_RAL_OP_COVERGROUP
  covergroup desired_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(fuse_1, fuse_1.desired)
     `RAL_FIELD_CP_1(fuse_1, fuse_1.desired, 0)
     `RAL_FIELD_CP(fuse_2, fuse_2.desired)
     `RAL_FIELD_CP_1(fuse_2, fuse_2.desired, 0)
     `RAL_FIELD_CP(fuse_3, fuse_3.desired)
     `RAL_FIELD_CP_1(fuse_3, fuse_3.desired, 0)
     `RAL_FIELD_CP(fuse_4, fuse_4.desired)
     `RAL_FIELD_CP_1(fuse_4, fuse_4.desired, 0)
  endgroup

  covergroup actual_cg @(cov_ev);
     option.per_instance = 1;
     `RAL_FIELD_CP(fuse_1, fuse_1.actual)
     `RAL_FIELD_CP_1(fuse_1, fuse_1.actual, 0)
     `RAL_FIELD_CP(fuse_2, fuse_2.actual)
     `RAL_FIELD_CP_1(fuse_2, fuse_2.actual, 0)
     `RAL_FIELD_CP(fuse_3, fuse_3.actual)
     `RAL_FIELD_CP_1(fuse_3, fuse_3.actual, 0)
     `RAL_FIELD_CP(fuse_4, fuse_4.actual)
     `RAL_FIELD_CP_1(fuse_4, fuse_4.actual, 0)
  endgroup
  `endif

  // --------------------------
  // add constraint based on database legal values
  // --------------------------
  function void build();
    fuse_1 = new("fuse_1", "RW", 1, 0, {""});
    fuse_1.set_rand_mode(0);
    void'(add_field( fuse_1 ));

    fuse_2 = new("fuse_2", "RW", 1, 1, {""});
    fuse_2.set_rand_mode(0);
    void'(add_field( fuse_2 ));

    fuse_3 = new("fuse_3", "RW", 1, 2, {""});
    fuse_3.set_rand_mode(0);
    void'(add_field( fuse_3 ));

    fuse_4 = new("fuse_4", "RW", 1, 3, {""});
    fuse_4.set_rand_mode(0);
    void'(add_field( fuse_4 ));

  endfunction

`DEFINE_NONE_SCOPE_REG_API(mby_fuse_mby_fuse_reg) 
endclass : mby_fuse_mby_fuse_reg

// ================================================

class mby_fuse_file extends sla_ral_file;

  rand mby_fuse_mby_fuse_reg mby_fuse;

  bit mby_fuse_create;

  `ovm_component_utils(mby_fuse_file)

  function new(string n, ovm_component p);
    super.new(n,p);
  endfunction

  function void instance_regs();
    if(instanceALL) begin
      mby_fuse_create = 1;
    end
    else begin
      mby_fuse.rand_mode(0);
    end
  endfunction

  // --------------------------
  function void build();
    `ifdef SLA_RAL_COVERAGE
    regfilename = this.get_name();
    `endif

    // call the function above before the register instantiation to determine which one to instance
    instance_regs();

    if(mby_fuse_create) begin
    `ifdef SLA_RAL_COVERAGE
      sla_ral_reg::regname = "mby_fuse";
    `endif
      mby_fuse = mby_fuse_mby_fuse_reg::type_id::create("mby_fuse", this);
      mby_fuse.set_cfg(16'h0, 16'h0, 16'h0, 4'h0, 32, 32'b00000000000000000000000000000000);
      if ( $test$plusargs("mby_fuse:dont_test") ) mby_fuse.set_test_reg(1'b0);
      if (!add_reg( mby_fuse )) begin
        `sla_error(get_name(), ("Could not add register mby_fuse"));
      end
    end

  endfunction

 virtual function void print_sv_ral_file();  
    $display("RAL File Type [%s], RAL File Instance [%s], SV File ---> %s", get_type_name(), get_name(), `__FILE__); 
 endfunction 
endclass : mby_fuse_file

// ================================================


`endif
