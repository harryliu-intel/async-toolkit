// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

//-----------------------------------------------------------------------------
// Title         : Egress hard reset sequence
// Project       : Madison Bay
//-----------------------------------------------------------------------------
// File          : mby_egr_hard_reset_seq.sv
// Author        : jose.j.godinez.carrillo  <jjgodine@ichips.intel.com>
// Created       : 22.08.2018
// Last modified : 22.08.2018
//-----------------------------------------------------------------------------
// Description :
//
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by Intel Corporation This model is the confidential and
// proprietary property of Intel Corporation and the possession or use of this
// file requires a written license from Intel Corporation.
//-----------------------------------------------------------------------------
// Modification history :
// 22.08.2018 : created
//-----------------------------------------------------------------------------

//-----------------------------------------------------------------------------
// Class: mby_egr_hard_reset_seq
//-----------------------------------------------------------------------------
import shdv_reset_pkg::*;
class mby_egr_mid_reset_seq extends mby_egr_extended_base_seq;

   shdv_reset_event        reset_event;
   shdv_reset_manager      reset_manager;
   shdv_reset_data         reset_data;

   `uvm_object_utils(mby_egr_mid_reset_seq)

   typedef enum {
      HARD_RESET,
      SOFT_RESET,
      POWER_GOOD
   }reset_type;

   rand int delay, duration;
   rand reset_type rst_type;

   constraint reset_select{
      soft rst_type == POWER_GOOD;
      soft duration  inside {[80:100]};
      soft delay     inside {[0:5]};
   }
   //--------------------------------------------------------------------------
   // Task: body()
   //--------------------------------------------------------------------------
   task body();

      virtual mby_egr_env_if  env_if;

      reset_data              = shdv_reset_data::type_id::create("reset_data");
      reset_data.rst_domain   = "egr";

      `uvm_info(get_name(), $sformatf("[RST_DBG]: reset scenario type = %s, delay = %0d, duration = %0d", rst_type.name(),delay,duration), UVM_NONE)
      case (rst_type)
         POWER_GOOD  : begin
            reset_data.rst_type  = "power_good";
            reset_event          = reset_manager.get_global("egr_power_good");
         end
         HARD_RESET  : begin
            reset_data.rst_type   = "hard";
            reset_event          = reset_manager.get_global("egr_reset");
         end
         SOFT_RESET  : reset_data.rst_type   = "soft";
         default  :  ;
      endcase

      wait_n(delay);
      `uvm_info(get_name(), "[RST_DBG]: Reset event triggered", UVM_LOW)
      reset_event.set(reset_data);

      wait_n(duration);
      `uvm_info(get_name(), "[RST_DBG]: Reset event cleared", UVM_LOW)
      reset_event.clear();


   endtask : body

endclass : mby_egr_mid_reset_seq
