magic
tech scmos
timestamp 962518978
<< ndiffusion >>
rect -220 -727 -214 -726
rect -220 -733 -214 -729
rect -220 -739 -214 -735
rect -220 -745 -214 -741
rect -220 -751 -214 -747
rect -220 -754 -214 -753
rect -220 -758 -218 -754
rect -220 -759 -214 -758
rect -220 -765 -214 -761
rect -220 -771 -214 -767
rect -220 -777 -214 -773
rect -220 -783 -214 -779
rect -220 -786 -214 -785
<< pdiffusion >>
rect -195 -717 -187 -714
rect -199 -718 -187 -717
rect -199 -722 -187 -720
rect -199 -726 -193 -722
rect -199 -727 -187 -726
rect -199 -730 -187 -729
rect -189 -734 -187 -730
rect -199 -735 -187 -734
rect -199 -738 -187 -737
rect -199 -742 -193 -738
rect -199 -743 -187 -742
rect -199 -746 -187 -745
rect -189 -750 -187 -746
rect -199 -751 -187 -750
rect -199 -754 -187 -753
rect -199 -758 -193 -754
rect -199 -759 -187 -758
rect -199 -762 -187 -761
rect -189 -766 -187 -762
rect -199 -767 -187 -766
rect -199 -770 -187 -769
rect -199 -774 -193 -770
rect -199 -775 -187 -774
rect -199 -778 -187 -777
rect -189 -782 -187 -778
rect -199 -783 -187 -782
rect -199 -786 -187 -785
<< ntransistor >>
rect -220 -729 -214 -727
rect -220 -735 -214 -733
rect -220 -741 -214 -739
rect -220 -747 -214 -745
rect -220 -753 -214 -751
rect -220 -761 -214 -759
rect -220 -767 -214 -765
rect -220 -773 -214 -771
rect -220 -779 -214 -777
rect -220 -785 -214 -783
<< ptransistor >>
rect -199 -720 -187 -718
rect -199 -729 -187 -727
rect -199 -737 -187 -735
rect -199 -745 -187 -743
rect -199 -753 -187 -751
rect -199 -761 -187 -759
rect -199 -769 -187 -767
rect -199 -777 -187 -775
rect -199 -785 -187 -783
<< polysilicon >>
rect -202 -720 -199 -718
rect -187 -720 -184 -718
rect -223 -729 -220 -727
rect -214 -729 -211 -727
rect -203 -729 -199 -727
rect -187 -729 -184 -727
rect -203 -733 -201 -729
rect -223 -735 -220 -733
rect -214 -735 -201 -733
rect -203 -737 -199 -735
rect -187 -737 -184 -735
rect -223 -741 -220 -739
rect -214 -741 -206 -739
rect -208 -743 -206 -741
rect -208 -745 -199 -743
rect -187 -745 -184 -743
rect -223 -747 -220 -745
rect -214 -747 -211 -745
rect -203 -751 -201 -745
rect -223 -753 -220 -751
rect -214 -753 -211 -751
rect -203 -753 -199 -751
rect -187 -753 -184 -751
rect -223 -761 -220 -759
rect -214 -761 -211 -759
rect -203 -761 -199 -759
rect -187 -761 -184 -759
rect -223 -767 -220 -765
rect -214 -767 -211 -765
rect -203 -767 -201 -761
rect -208 -769 -199 -767
rect -187 -769 -184 -767
rect -208 -771 -206 -769
rect -223 -773 -220 -771
rect -214 -773 -206 -771
rect -203 -777 -199 -775
rect -187 -777 -184 -775
rect -223 -779 -220 -777
rect -214 -779 -201 -777
rect -203 -783 -201 -779
rect -223 -785 -220 -783
rect -214 -785 -211 -783
rect -203 -785 -199 -783
rect -187 -785 -184 -783
<< ndcontact >>
rect -220 -726 -214 -722
rect -218 -758 -214 -754
rect -220 -790 -214 -786
<< pdcontact >>
rect -199 -717 -195 -713
rect -193 -726 -187 -722
rect -199 -734 -189 -730
rect -193 -742 -187 -738
rect -199 -750 -189 -746
rect -193 -758 -187 -754
rect -199 -766 -189 -762
rect -193 -774 -187 -770
rect -199 -782 -189 -778
rect -199 -790 -187 -786
<< metal1 >>
rect -199 -717 -195 -713
rect -220 -726 -214 -722
rect -199 -730 -196 -717
rect -193 -726 -187 -722
rect -199 -734 -189 -730
rect -199 -746 -196 -734
rect -193 -742 -187 -738
rect -199 -750 -189 -746
rect -199 -754 -196 -750
rect -218 -758 -196 -754
rect -193 -758 -187 -754
rect -199 -762 -196 -758
rect -199 -766 -189 -762
rect -199 -778 -196 -766
rect -193 -774 -187 -770
rect -199 -782 -189 -778
rect -220 -790 -214 -786
rect -199 -790 -187 -786
<< labels >>
rlabel polysilicon -186 -784 -186 -784 7 a
rlabel polysilicon -186 -776 -186 -776 7 a
rlabel polysilicon -186 -768 -186 -768 7 b
rlabel polysilicon -186 -760 -186 -760 7 b
rlabel polysilicon -186 -752 -186 -752 7 c
rlabel polysilicon -186 -744 -186 -744 7 c
rlabel polysilicon -186 -736 -186 -736 7 d
rlabel polysilicon -186 -728 -186 -728 7 d
rlabel space -191 -791 -184 -723 3 ^p
rlabel polysilicon -221 -734 -221 -734 3 d
rlabel polysilicon -221 -740 -221 -740 3 c
rlabel polysilicon -221 -746 -221 -746 3 b
rlabel polysilicon -221 -752 -221 -752 3 a
rlabel polysilicon -221 -760 -221 -760 3 d
rlabel polysilicon -221 -766 -221 -766 3 c
rlabel polysilicon -221 -772 -221 -772 3 b
rlabel polysilicon -221 -778 -221 -778 3 a
rlabel polysilicon -221 -784 -221 -784 3 _SReset!
rlabel polysilicon -221 -728 -221 -728 3 _SReset!
rlabel space -223 -791 -217 -721 7 ^n
rlabel polysilicon -186 -719 -186 -719 1 _PReset!
rlabel pdcontact -197 -732 -197 -732 1 x
rlabel pdcontact -197 -748 -197 -748 1 x
rlabel pdcontact -197 -764 -197 -764 1 x
rlabel pdcontact -197 -780 -197 -780 1 x
rlabel pdcontact -190 -772 -190 -772 1 Vdd!
rlabel pdcontact -190 -756 -190 -756 1 Vdd!
rlabel pdcontact -190 -740 -190 -740 1 Vdd!
rlabel pdcontact -190 -724 -190 -724 1 Vdd!
rlabel pdcontact -190 -788 -190 -788 1 Vdd!
rlabel ndcontact -216 -756 -216 -756 1 x
rlabel ndcontact -216 -724 -216 -724 5 GND!
rlabel ndcontact -216 -788 -216 -788 1 GND!
rlabel pdcontact -197 -715 -197 -715 5 x
<< end >>
