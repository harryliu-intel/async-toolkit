///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_mst_glort_map.sv                                   
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_mst_glort_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_FF
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_FF

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_RSTD


module rtlgen_mby_ppe_mst_glort_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_mst_glort_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_PH2_FF
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_MST_GLORT_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_MST_GLORT_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_mst_glort_map ( //lintra s-2096
    // Clocks


    // Resets



    // Register Inputs
    handcode_reg_rdata_CGRP_USED_TABLE,
    handcode_reg_rdata_EGRESS_MST_TABLE,
    handcode_reg_rdata_EGRESS_VID_CFG,
    handcode_reg_rdata_EGRESS_VID_TABLE,
    handcode_reg_rdata_GLORT_CAM,
    handcode_reg_rdata_GLORT_DIRECT_MAP_CTRL,
    handcode_reg_rdata_GLORT_DIRECT_MAP_DST0,
    handcode_reg_rdata_GLORT_DIRECT_MAP_DST1,
    handcode_reg_rdata_GLORT_DIRECT_MAP_DST2,
    handcode_reg_rdata_GLORT_DIRECT_MAP_DST3,
    handcode_reg_rdata_GLORT_DIRECT_MAP_DST4,
    handcode_reg_rdata_GLORT_RAM,
    handcode_reg_rdata_INGRESS_MST_TABLE,

    handcode_rvalid_CGRP_USED_TABLE,
    handcode_rvalid_EGRESS_MST_TABLE,
    handcode_rvalid_EGRESS_VID_CFG,
    handcode_rvalid_EGRESS_VID_TABLE,
    handcode_rvalid_GLORT_CAM,
    handcode_rvalid_GLORT_DIRECT_MAP_CTRL,
    handcode_rvalid_GLORT_DIRECT_MAP_DST0,
    handcode_rvalid_GLORT_DIRECT_MAP_DST1,
    handcode_rvalid_GLORT_DIRECT_MAP_DST2,
    handcode_rvalid_GLORT_DIRECT_MAP_DST3,
    handcode_rvalid_GLORT_DIRECT_MAP_DST4,
    handcode_rvalid_GLORT_RAM,
    handcode_rvalid_INGRESS_MST_TABLE,

    handcode_wvalid_CGRP_USED_TABLE,
    handcode_wvalid_EGRESS_MST_TABLE,
    handcode_wvalid_EGRESS_VID_CFG,
    handcode_wvalid_EGRESS_VID_TABLE,
    handcode_wvalid_GLORT_CAM,
    handcode_wvalid_GLORT_DIRECT_MAP_CTRL,
    handcode_wvalid_GLORT_DIRECT_MAP_DST0,
    handcode_wvalid_GLORT_DIRECT_MAP_DST1,
    handcode_wvalid_GLORT_DIRECT_MAP_DST2,
    handcode_wvalid_GLORT_DIRECT_MAP_DST3,
    handcode_wvalid_GLORT_DIRECT_MAP_DST4,
    handcode_wvalid_GLORT_RAM,
    handcode_wvalid_INGRESS_MST_TABLE,

    handcode_error_CGRP_USED_TABLE,
    handcode_error_EGRESS_MST_TABLE,
    handcode_error_EGRESS_VID_CFG,
    handcode_error_EGRESS_VID_TABLE,
    handcode_error_GLORT_CAM,
    handcode_error_GLORT_DIRECT_MAP_CTRL,
    handcode_error_GLORT_DIRECT_MAP_DST0,
    handcode_error_GLORT_DIRECT_MAP_DST1,
    handcode_error_GLORT_DIRECT_MAP_DST2,
    handcode_error_GLORT_DIRECT_MAP_DST3,
    handcode_error_GLORT_DIRECT_MAP_DST4,
    handcode_error_GLORT_RAM,
    handcode_error_INGRESS_MST_TABLE,


    // Register Outputs

    // Register signals for HandCoded registers
    handcode_reg_wdata_CGRP_USED_TABLE,
    handcode_reg_wdata_EGRESS_MST_TABLE,
    handcode_reg_wdata_EGRESS_VID_CFG,
    handcode_reg_wdata_EGRESS_VID_TABLE,
    handcode_reg_wdata_GLORT_CAM,
    handcode_reg_wdata_GLORT_DIRECT_MAP_CTRL,
    handcode_reg_wdata_GLORT_DIRECT_MAP_DST0,
    handcode_reg_wdata_GLORT_DIRECT_MAP_DST1,
    handcode_reg_wdata_GLORT_DIRECT_MAP_DST2,
    handcode_reg_wdata_GLORT_DIRECT_MAP_DST3,
    handcode_reg_wdata_GLORT_DIRECT_MAP_DST4,
    handcode_reg_wdata_GLORT_RAM,
    handcode_reg_wdata_INGRESS_MST_TABLE,

    we_CGRP_USED_TABLE,
    we_EGRESS_MST_TABLE,
    we_EGRESS_VID_CFG,
    we_EGRESS_VID_TABLE,
    we_GLORT_CAM,
    we_GLORT_DIRECT_MAP_CTRL,
    we_GLORT_DIRECT_MAP_DST0,
    we_GLORT_DIRECT_MAP_DST1,
    we_GLORT_DIRECT_MAP_DST2,
    we_GLORT_DIRECT_MAP_DST3,
    we_GLORT_DIRECT_MAP_DST4,
    we_GLORT_RAM,
    we_INGRESS_MST_TABLE,

    re_CGRP_USED_TABLE,
    re_EGRESS_MST_TABLE,
    re_EGRESS_VID_CFG,
    re_EGRESS_VID_TABLE,
    re_GLORT_CAM,
    re_GLORT_DIRECT_MAP_CTRL,
    re_GLORT_DIRECT_MAP_DST0,
    re_GLORT_DIRECT_MAP_DST1,
    re_GLORT_DIRECT_MAP_DST2,
    re_GLORT_DIRECT_MAP_DST3,
    re_GLORT_DIRECT_MAP_DST4,
    re_GLORT_RAM,
    re_INGRESS_MST_TABLE,




    // Config Access
    req,
    ack
    

);

import mby_ppe_mst_glort_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:0] MBY_PPE_MST_GLORT_MAP_OFFSET = {MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] MST_GLORT_SB_BAR = 3'b0;
parameter [7:0] MST_GLORT_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;

    // Clocks


    // Resets



    // Register Inputs
input CGRP_USED_TABLE_t  handcode_reg_rdata_CGRP_USED_TABLE;
input EGRESS_MST_TABLE_t  handcode_reg_rdata_EGRESS_MST_TABLE;
input EGRESS_VID_CFG_t  handcode_reg_rdata_EGRESS_VID_CFG;
input EGRESS_VID_TABLE_t  handcode_reg_rdata_EGRESS_VID_TABLE;
input GLORT_CAM_t  handcode_reg_rdata_GLORT_CAM;
input GLORT_DIRECT_MAP_CTRL_t  handcode_reg_rdata_GLORT_DIRECT_MAP_CTRL;
input GLORT_DIRECT_MAP_DST0_t  handcode_reg_rdata_GLORT_DIRECT_MAP_DST0;
input GLORT_DIRECT_MAP_DST1_t  handcode_reg_rdata_GLORT_DIRECT_MAP_DST1;
input GLORT_DIRECT_MAP_DST2_t  handcode_reg_rdata_GLORT_DIRECT_MAP_DST2;
input GLORT_DIRECT_MAP_DST3_t  handcode_reg_rdata_GLORT_DIRECT_MAP_DST3;
input GLORT_DIRECT_MAP_DST4_t  handcode_reg_rdata_GLORT_DIRECT_MAP_DST4;
input GLORT_RAM_t  handcode_reg_rdata_GLORT_RAM;
input INGRESS_MST_TABLE_t  handcode_reg_rdata_INGRESS_MST_TABLE;

input handcode_rvalid_CGRP_USED_TABLE_t  handcode_rvalid_CGRP_USED_TABLE;
input handcode_rvalid_EGRESS_MST_TABLE_t  handcode_rvalid_EGRESS_MST_TABLE;
input handcode_rvalid_EGRESS_VID_CFG_t  handcode_rvalid_EGRESS_VID_CFG;
input handcode_rvalid_EGRESS_VID_TABLE_t  handcode_rvalid_EGRESS_VID_TABLE;
input handcode_rvalid_GLORT_CAM_t  handcode_rvalid_GLORT_CAM;
input handcode_rvalid_GLORT_DIRECT_MAP_CTRL_t  handcode_rvalid_GLORT_DIRECT_MAP_CTRL;
input handcode_rvalid_GLORT_DIRECT_MAP_DST0_t  handcode_rvalid_GLORT_DIRECT_MAP_DST0;
input handcode_rvalid_GLORT_DIRECT_MAP_DST1_t  handcode_rvalid_GLORT_DIRECT_MAP_DST1;
input handcode_rvalid_GLORT_DIRECT_MAP_DST2_t  handcode_rvalid_GLORT_DIRECT_MAP_DST2;
input handcode_rvalid_GLORT_DIRECT_MAP_DST3_t  handcode_rvalid_GLORT_DIRECT_MAP_DST3;
input handcode_rvalid_GLORT_DIRECT_MAP_DST4_t  handcode_rvalid_GLORT_DIRECT_MAP_DST4;
input handcode_rvalid_GLORT_RAM_t  handcode_rvalid_GLORT_RAM;
input handcode_rvalid_INGRESS_MST_TABLE_t  handcode_rvalid_INGRESS_MST_TABLE;

input handcode_wvalid_CGRP_USED_TABLE_t  handcode_wvalid_CGRP_USED_TABLE;
input handcode_wvalid_EGRESS_MST_TABLE_t  handcode_wvalid_EGRESS_MST_TABLE;
input handcode_wvalid_EGRESS_VID_CFG_t  handcode_wvalid_EGRESS_VID_CFG;
input handcode_wvalid_EGRESS_VID_TABLE_t  handcode_wvalid_EGRESS_VID_TABLE;
input handcode_wvalid_GLORT_CAM_t  handcode_wvalid_GLORT_CAM;
input handcode_wvalid_GLORT_DIRECT_MAP_CTRL_t  handcode_wvalid_GLORT_DIRECT_MAP_CTRL;
input handcode_wvalid_GLORT_DIRECT_MAP_DST0_t  handcode_wvalid_GLORT_DIRECT_MAP_DST0;
input handcode_wvalid_GLORT_DIRECT_MAP_DST1_t  handcode_wvalid_GLORT_DIRECT_MAP_DST1;
input handcode_wvalid_GLORT_DIRECT_MAP_DST2_t  handcode_wvalid_GLORT_DIRECT_MAP_DST2;
input handcode_wvalid_GLORT_DIRECT_MAP_DST3_t  handcode_wvalid_GLORT_DIRECT_MAP_DST3;
input handcode_wvalid_GLORT_DIRECT_MAP_DST4_t  handcode_wvalid_GLORT_DIRECT_MAP_DST4;
input handcode_wvalid_GLORT_RAM_t  handcode_wvalid_GLORT_RAM;
input handcode_wvalid_INGRESS_MST_TABLE_t  handcode_wvalid_INGRESS_MST_TABLE;

input handcode_error_CGRP_USED_TABLE_t  handcode_error_CGRP_USED_TABLE;
input handcode_error_EGRESS_MST_TABLE_t  handcode_error_EGRESS_MST_TABLE;
input handcode_error_EGRESS_VID_CFG_t  handcode_error_EGRESS_VID_CFG;
input handcode_error_EGRESS_VID_TABLE_t  handcode_error_EGRESS_VID_TABLE;
input handcode_error_GLORT_CAM_t  handcode_error_GLORT_CAM;
input handcode_error_GLORT_DIRECT_MAP_CTRL_t  handcode_error_GLORT_DIRECT_MAP_CTRL;
input handcode_error_GLORT_DIRECT_MAP_DST0_t  handcode_error_GLORT_DIRECT_MAP_DST0;
input handcode_error_GLORT_DIRECT_MAP_DST1_t  handcode_error_GLORT_DIRECT_MAP_DST1;
input handcode_error_GLORT_DIRECT_MAP_DST2_t  handcode_error_GLORT_DIRECT_MAP_DST2;
input handcode_error_GLORT_DIRECT_MAP_DST3_t  handcode_error_GLORT_DIRECT_MAP_DST3;
input handcode_error_GLORT_DIRECT_MAP_DST4_t  handcode_error_GLORT_DIRECT_MAP_DST4;
input handcode_error_GLORT_RAM_t  handcode_error_GLORT_RAM;
input handcode_error_INGRESS_MST_TABLE_t  handcode_error_INGRESS_MST_TABLE;


    // Register Outputs

    // Register signals for HandCoded registers
output CGRP_USED_TABLE_t  handcode_reg_wdata_CGRP_USED_TABLE;
output EGRESS_MST_TABLE_t  handcode_reg_wdata_EGRESS_MST_TABLE;
output EGRESS_VID_CFG_t  handcode_reg_wdata_EGRESS_VID_CFG;
output EGRESS_VID_TABLE_t  handcode_reg_wdata_EGRESS_VID_TABLE;
output GLORT_CAM_t  handcode_reg_wdata_GLORT_CAM;
output GLORT_DIRECT_MAP_CTRL_t  handcode_reg_wdata_GLORT_DIRECT_MAP_CTRL;
output GLORT_DIRECT_MAP_DST0_t  handcode_reg_wdata_GLORT_DIRECT_MAP_DST0;
output GLORT_DIRECT_MAP_DST1_t  handcode_reg_wdata_GLORT_DIRECT_MAP_DST1;
output GLORT_DIRECT_MAP_DST2_t  handcode_reg_wdata_GLORT_DIRECT_MAP_DST2;
output GLORT_DIRECT_MAP_DST3_t  handcode_reg_wdata_GLORT_DIRECT_MAP_DST3;
output GLORT_DIRECT_MAP_DST4_t  handcode_reg_wdata_GLORT_DIRECT_MAP_DST4;
output GLORT_RAM_t  handcode_reg_wdata_GLORT_RAM;
output INGRESS_MST_TABLE_t  handcode_reg_wdata_INGRESS_MST_TABLE;

output we_CGRP_USED_TABLE_t  we_CGRP_USED_TABLE;
output we_EGRESS_MST_TABLE_t  we_EGRESS_MST_TABLE;
output we_EGRESS_VID_CFG_t  we_EGRESS_VID_CFG;
output we_EGRESS_VID_TABLE_t  we_EGRESS_VID_TABLE;
output we_GLORT_CAM_t  we_GLORT_CAM;
output we_GLORT_DIRECT_MAP_CTRL_t  we_GLORT_DIRECT_MAP_CTRL;
output we_GLORT_DIRECT_MAP_DST0_t  we_GLORT_DIRECT_MAP_DST0;
output we_GLORT_DIRECT_MAP_DST1_t  we_GLORT_DIRECT_MAP_DST1;
output we_GLORT_DIRECT_MAP_DST2_t  we_GLORT_DIRECT_MAP_DST2;
output we_GLORT_DIRECT_MAP_DST3_t  we_GLORT_DIRECT_MAP_DST3;
output we_GLORT_DIRECT_MAP_DST4_t  we_GLORT_DIRECT_MAP_DST4;
output we_GLORT_RAM_t  we_GLORT_RAM;
output we_INGRESS_MST_TABLE_t  we_INGRESS_MST_TABLE;

output re_CGRP_USED_TABLE_t  re_CGRP_USED_TABLE;
output re_EGRESS_MST_TABLE_t  re_EGRESS_MST_TABLE;
output re_EGRESS_VID_CFG_t  re_EGRESS_VID_CFG;
output re_EGRESS_VID_TABLE_t  re_EGRESS_VID_TABLE;
output re_GLORT_CAM_t  re_GLORT_CAM;
output re_GLORT_DIRECT_MAP_CTRL_t  re_GLORT_DIRECT_MAP_CTRL;
output re_GLORT_DIRECT_MAP_DST0_t  re_GLORT_DIRECT_MAP_DST0;
output re_GLORT_DIRECT_MAP_DST1_t  re_GLORT_DIRECT_MAP_DST1;
output re_GLORT_DIRECT_MAP_DST2_t  re_GLORT_DIRECT_MAP_DST2;
output re_GLORT_DIRECT_MAP_DST3_t  re_GLORT_DIRECT_MAP_DST3;
output re_GLORT_DIRECT_MAP_DST4_t  re_GLORT_DIRECT_MAP_DST4;
output re_GLORT_RAM_t  re_GLORT_RAM;
output re_INGRESS_MST_TABLE_t  re_INGRESS_MST_TABLE;




    // Config Access
input mby_ppe_mst_glort_map_cr_req_t  req;
output mby_ppe_mst_glort_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_mst_glort_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_MST_GLORT_MAP_MEM;
assign case_req_addr_MBY_PPE_MST_GLORT_MAP_MEM = req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_mst_glort;
always_comb begin : sb_fid_cond_mst_glort_BLOCK
    unique casez (req_fid) 
		MST_GLORT_SB_FID: sb_fid_cond_mst_glort = 1;
		default: sb_fid_cond_mst_glort = 0;
    endcase 
end


logic sb_bar_cond_mst_glort;
always_comb begin : sb_bar_cond_mst_glort_BLOCK
    unique casez (req_bar) 
		MST_GLORT_SB_BAR: sb_bar_cond_mst_glort = 1;
		default: sb_bar_cond_mst_glort = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// EGRESS_VID_TABLE using HANDCODED_REG template.
logic addr_decode_EGRESS_VID_TABLE;
logic write_req_EGRESS_VID_TABLE;
logic read_req_EGRESS_VID_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b0??,8'h??,4'b??0?,1'b?},
      {32'b0??,8'h??,4'b??10,1'b0}:
          addr_decode_EGRESS_VID_TABLE = req.valid;
      default: 
         addr_decode_EGRESS_VID_TABLE = 1'b0; 
   endcase
end

always_comb write_req_EGRESS_VID_TABLE = f_IsMEMWr(req_opcode) && addr_decode_EGRESS_VID_TABLE ;
always_comb read_req_EGRESS_VID_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_EGRESS_VID_TABLE ;

always_comb we_EGRESS_VID_TABLE = {8{write_req_EGRESS_VID_TABLE}} & be;
always_comb re_EGRESS_VID_TABLE = {8{read_req_EGRESS_VID_TABLE}} & be;
always_comb handcode_reg_wdata_EGRESS_VID_TABLE = write_data;


// ----------------------------------------------------------------------
// EGRESS_VID_CFG using HANDCODED_REG template.
logic addr_decode_EGRESS_VID_CFG;
logic write_req_EGRESS_VID_CFG;
logic read_req_EGRESS_VID_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h4,4'b0???,8'h??,1'b?}: 
         addr_decode_EGRESS_VID_CFG = req.valid;
      default: 
         addr_decode_EGRESS_VID_CFG = 1'b0; 
   endcase
end

always_comb write_req_EGRESS_VID_CFG = f_IsMEMWr(req_opcode) && addr_decode_EGRESS_VID_CFG ;
always_comb read_req_EGRESS_VID_CFG  = f_IsMEMRd(req_opcode) && addr_decode_EGRESS_VID_CFG ;

always_comb we_EGRESS_VID_CFG = {8{write_req_EGRESS_VID_CFG}} & be;
always_comb re_EGRESS_VID_CFG = {8{read_req_EGRESS_VID_CFG}} & be;
always_comb handcode_reg_wdata_EGRESS_VID_CFG = write_data;


// ----------------------------------------------------------------------
// INGRESS_MST_TABLE using HANDCODED_REG template.
logic addr_decode_INGRESS_MST_TABLE;
logic write_req_INGRESS_MST_TABLE;
logic read_req_INGRESS_MST_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h4,4'b1???,8'h??,1'b?}: 
         addr_decode_INGRESS_MST_TABLE = req.valid;
      default: 
         addr_decode_INGRESS_MST_TABLE = 1'b0; 
   endcase
end

always_comb write_req_INGRESS_MST_TABLE = f_IsMEMWr(req_opcode) && addr_decode_INGRESS_MST_TABLE ;
always_comb read_req_INGRESS_MST_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_INGRESS_MST_TABLE ;

always_comb we_INGRESS_MST_TABLE = {8{write_req_INGRESS_MST_TABLE}} & be;
always_comb re_INGRESS_MST_TABLE = {8{read_req_INGRESS_MST_TABLE}} & be;
always_comb handcode_reg_wdata_INGRESS_MST_TABLE = write_data;


// ----------------------------------------------------------------------
// EGRESS_MST_TABLE using HANDCODED_REG template.
logic addr_decode_EGRESS_MST_TABLE;
logic write_req_EGRESS_MST_TABLE;
logic read_req_EGRESS_MST_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b10??,8'h??,4'b??0?,1'b?},
      {32'b10??,8'h??,4'b??10,1'b0}:
          addr_decode_EGRESS_MST_TABLE = req.valid;
      default: 
         addr_decode_EGRESS_MST_TABLE = 1'b0; 
   endcase
end

always_comb write_req_EGRESS_MST_TABLE = f_IsMEMWr(req_opcode) && addr_decode_EGRESS_MST_TABLE ;
always_comb read_req_EGRESS_MST_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_EGRESS_MST_TABLE ;

always_comb we_EGRESS_MST_TABLE = {8{write_req_EGRESS_MST_TABLE}} & be;
always_comb re_EGRESS_MST_TABLE = {8{read_req_EGRESS_MST_TABLE}} & be;
always_comb handcode_reg_wdata_EGRESS_MST_TABLE = write_data;


// ----------------------------------------------------------------------
// GLORT_DIRECT_MAP_CTRL using HANDCODED_REG template.
logic addr_decode_GLORT_DIRECT_MAP_CTRL;
logic write_req_GLORT_DIRECT_MAP_CTRL;
logic read_req_GLORT_DIRECT_MAP_CTRL;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'hC000,1'b0}: 
         addr_decode_GLORT_DIRECT_MAP_CTRL = req.valid;
      default: 
         addr_decode_GLORT_DIRECT_MAP_CTRL = 1'b0; 
   endcase
end

always_comb write_req_GLORT_DIRECT_MAP_CTRL = f_IsMEMWr(req_opcode) && addr_decode_GLORT_DIRECT_MAP_CTRL ;
always_comb read_req_GLORT_DIRECT_MAP_CTRL  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_DIRECT_MAP_CTRL ;

always_comb we_GLORT_DIRECT_MAP_CTRL = {8{write_req_GLORT_DIRECT_MAP_CTRL}} & be;
always_comb re_GLORT_DIRECT_MAP_CTRL = {8{read_req_GLORT_DIRECT_MAP_CTRL}} & be;
always_comb handcode_reg_wdata_GLORT_DIRECT_MAP_CTRL = write_data;


// ----------------------------------------------------------------------
// GLORT_DIRECT_MAP_DST0 using HANDCODED_REG template.
logic addr_decode_GLORT_DIRECT_MAP_DST0;
logic write_req_GLORT_DIRECT_MAP_DST0;
logic read_req_GLORT_DIRECT_MAP_DST0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'hC000,1'b1}: 
         addr_decode_GLORT_DIRECT_MAP_DST0 = req.valid;
      default: 
         addr_decode_GLORT_DIRECT_MAP_DST0 = 1'b0; 
   endcase
end

always_comb write_req_GLORT_DIRECT_MAP_DST0 = f_IsMEMWr(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST0 ;
always_comb read_req_GLORT_DIRECT_MAP_DST0  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST0 ;

always_comb we_GLORT_DIRECT_MAP_DST0 = {8{write_req_GLORT_DIRECT_MAP_DST0}} & be;
always_comb re_GLORT_DIRECT_MAP_DST0 = {8{read_req_GLORT_DIRECT_MAP_DST0}} & be;
always_comb handcode_reg_wdata_GLORT_DIRECT_MAP_DST0 = write_data;


// ----------------------------------------------------------------------
// GLORT_DIRECT_MAP_DST1 using HANDCODED_REG template.
logic addr_decode_GLORT_DIRECT_MAP_DST1;
logic write_req_GLORT_DIRECT_MAP_DST1;
logic read_req_GLORT_DIRECT_MAP_DST1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'hC001,1'b0}: 
         addr_decode_GLORT_DIRECT_MAP_DST1 = req.valid;
      default: 
         addr_decode_GLORT_DIRECT_MAP_DST1 = 1'b0; 
   endcase
end

always_comb write_req_GLORT_DIRECT_MAP_DST1 = f_IsMEMWr(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST1 ;
always_comb read_req_GLORT_DIRECT_MAP_DST1  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST1 ;

always_comb we_GLORT_DIRECT_MAP_DST1 = {8{write_req_GLORT_DIRECT_MAP_DST1}} & be;
always_comb re_GLORT_DIRECT_MAP_DST1 = {8{read_req_GLORT_DIRECT_MAP_DST1}} & be;
always_comb handcode_reg_wdata_GLORT_DIRECT_MAP_DST1 = write_data;


// ----------------------------------------------------------------------
// GLORT_DIRECT_MAP_DST2 using HANDCODED_REG template.
logic addr_decode_GLORT_DIRECT_MAP_DST2;
logic write_req_GLORT_DIRECT_MAP_DST2;
logic read_req_GLORT_DIRECT_MAP_DST2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'hC001,1'b1}: 
         addr_decode_GLORT_DIRECT_MAP_DST2 = req.valid;
      default: 
         addr_decode_GLORT_DIRECT_MAP_DST2 = 1'b0; 
   endcase
end

always_comb write_req_GLORT_DIRECT_MAP_DST2 = f_IsMEMWr(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST2 ;
always_comb read_req_GLORT_DIRECT_MAP_DST2  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST2 ;

always_comb we_GLORT_DIRECT_MAP_DST2 = {8{write_req_GLORT_DIRECT_MAP_DST2}} & be;
always_comb re_GLORT_DIRECT_MAP_DST2 = {8{read_req_GLORT_DIRECT_MAP_DST2}} & be;
always_comb handcode_reg_wdata_GLORT_DIRECT_MAP_DST2 = write_data;


// ----------------------------------------------------------------------
// GLORT_DIRECT_MAP_DST3 using HANDCODED_REG template.
logic addr_decode_GLORT_DIRECT_MAP_DST3;
logic write_req_GLORT_DIRECT_MAP_DST3;
logic read_req_GLORT_DIRECT_MAP_DST3;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'hC002,1'b0}: 
         addr_decode_GLORT_DIRECT_MAP_DST3 = req.valid;
      default: 
         addr_decode_GLORT_DIRECT_MAP_DST3 = 1'b0; 
   endcase
end

always_comb write_req_GLORT_DIRECT_MAP_DST3 = f_IsMEMWr(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST3 ;
always_comb read_req_GLORT_DIRECT_MAP_DST3  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST3 ;

always_comb we_GLORT_DIRECT_MAP_DST3 = {8{write_req_GLORT_DIRECT_MAP_DST3}} & be;
always_comb re_GLORT_DIRECT_MAP_DST3 = {8{read_req_GLORT_DIRECT_MAP_DST3}} & be;
always_comb handcode_reg_wdata_GLORT_DIRECT_MAP_DST3 = write_data;


// ----------------------------------------------------------------------
// GLORT_DIRECT_MAP_DST4 using HANDCODED_REG template.
logic addr_decode_GLORT_DIRECT_MAP_DST4;
logic write_req_GLORT_DIRECT_MAP_DST4;
logic read_req_GLORT_DIRECT_MAP_DST4;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'hC002,1'b1}: 
         addr_decode_GLORT_DIRECT_MAP_DST4 = req.valid;
      default: 
         addr_decode_GLORT_DIRECT_MAP_DST4 = 1'b0; 
   endcase
end

always_comb write_req_GLORT_DIRECT_MAP_DST4 = f_IsMEMWr(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST4 ;
always_comb read_req_GLORT_DIRECT_MAP_DST4  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_DIRECT_MAP_DST4 ;

always_comb we_GLORT_DIRECT_MAP_DST4 = {8{write_req_GLORT_DIRECT_MAP_DST4}} & be;
always_comb re_GLORT_DIRECT_MAP_DST4 = {8{read_req_GLORT_DIRECT_MAP_DST4}} & be;
always_comb handcode_reg_wdata_GLORT_DIRECT_MAP_DST4 = write_data;


// ----------------------------------------------------------------------
// GLORT_RAM using HANDCODED_REG template.
logic addr_decode_GLORT_RAM;
logic write_req_GLORT_RAM;
logic read_req_GLORT_RAM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'hC0,4'b001?,4'h?,1'b?}: 
         addr_decode_GLORT_RAM = req.valid;
      default: 
         addr_decode_GLORT_RAM = 1'b0; 
   endcase
end

always_comb write_req_GLORT_RAM = f_IsMEMWr(req_opcode) && addr_decode_GLORT_RAM ;
always_comb read_req_GLORT_RAM  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_RAM ;

always_comb we_GLORT_RAM = {8{write_req_GLORT_RAM}} & be;
always_comb re_GLORT_RAM = {8{read_req_GLORT_RAM}} & be;
always_comb handcode_reg_wdata_GLORT_RAM = write_data;


// ----------------------------------------------------------------------
// GLORT_CAM using HANDCODED_REG template.
logic addr_decode_GLORT_CAM;
logic write_req_GLORT_CAM;
logic read_req_GLORT_CAM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'hC0,4'b010?,4'h?,1'b?}: 
         addr_decode_GLORT_CAM = req.valid;
      default: 
         addr_decode_GLORT_CAM = 1'b0; 
   endcase
end

always_comb write_req_GLORT_CAM = f_IsMEMWr(req_opcode) && addr_decode_GLORT_CAM ;
always_comb read_req_GLORT_CAM  = f_IsMEMRd(req_opcode) && addr_decode_GLORT_CAM ;

always_comb we_GLORT_CAM = {8{write_req_GLORT_CAM}} & be;
always_comb re_GLORT_CAM = {8{read_req_GLORT_CAM}} & be;
always_comb handcode_reg_wdata_GLORT_CAM = write_data;


// ----------------------------------------------------------------------
// CGRP_USED_TABLE using HANDCODED_REG template.
logic addr_decode_CGRP_USED_TABLE;
logic write_req_CGRP_USED_TABLE;
logic read_req_CGRP_USED_TABLE;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MST_GLORT_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'hC07,4'b011?,1'b?},
      {40'hC07,4'b1???,1'b?},
      {44'hC08?,1'b?},
      {40'hC09,4'b00??,1'b?},
      {40'hC09,4'b010?,1'b?},
      {44'hC096,1'b0}:
          addr_decode_CGRP_USED_TABLE = req.valid;
      default: 
         addr_decode_CGRP_USED_TABLE = 1'b0; 
   endcase
end

always_comb write_req_CGRP_USED_TABLE = f_IsMEMWr(req_opcode) && addr_decode_CGRP_USED_TABLE ;
always_comb read_req_CGRP_USED_TABLE  = f_IsMEMRd(req_opcode) && addr_decode_CGRP_USED_TABLE ;

always_comb we_CGRP_USED_TABLE = {8{write_req_CGRP_USED_TABLE}} & be;
always_comb re_CGRP_USED_TABLE = {8{read_req_CGRP_USED_TABLE}} & be;
always_comb handcode_reg_wdata_CGRP_USED_TABLE = write_data;


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_MST_GLORT_MAP_MEM) 
           {32'b0??,8'h??,4'b??0?,1'b?},
           {32'b0??,8'h??,4'b??10,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_EGRESS_VID_TABLE;
                    ack.read_miss = handcode_error_EGRESS_VID_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h4,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_EGRESS_VID_CFG;
                    ack.read_miss = handcode_error_EGRESS_VID_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h4,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_INGRESS_MST_TABLE;
                    ack.read_miss = handcode_error_INGRESS_MST_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b10??,8'h??,4'b??0?,1'b?},
           {32'b10??,8'h??,4'b??10,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_EGRESS_MST_TABLE;
                    ack.read_miss = handcode_error_EGRESS_MST_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'hC000,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_DIRECT_MAP_CTRL;
                    ack.read_miss = handcode_error_GLORT_DIRECT_MAP_CTRL;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'hC000,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_DIRECT_MAP_DST0;
                    ack.read_miss = handcode_error_GLORT_DIRECT_MAP_DST0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'hC001,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_DIRECT_MAP_DST1;
                    ack.read_miss = handcode_error_GLORT_DIRECT_MAP_DST1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'hC001,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_DIRECT_MAP_DST2;
                    ack.read_miss = handcode_error_GLORT_DIRECT_MAP_DST2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'hC002,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_DIRECT_MAP_DST3;
                    ack.read_miss = handcode_error_GLORT_DIRECT_MAP_DST3;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'hC002,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_DIRECT_MAP_DST4;
                    ack.read_miss = handcode_error_GLORT_DIRECT_MAP_DST4;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'hC0,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_RAM;
                    ack.read_miss = handcode_error_GLORT_RAM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'hC0,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_GLORT_CAM;
                    ack.read_miss = handcode_error_GLORT_CAM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'hC07,4'b011?,1'b?},
           {40'hC07,4'b1???,1'b?},
           {44'hC08?,1'b?},
           {40'hC09,4'b00??,1'b?},
           {40'hC09,4'b010?,1'b?},
           {44'hC096,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_CGRP_USED_TABLE;
                    ack.read_miss = handcode_error_CGRP_USED_TABLE;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_MST_GLORT_MAP_MEM) 
           {32'b0??,8'h??,4'b??0?,1'b?},
           {32'b0??,8'h??,4'b??10,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_EGRESS_VID_TABLE;
                    ack.write_miss = handcode_error_EGRESS_VID_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h4,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_EGRESS_VID_CFG;
                    ack.write_miss = handcode_error_EGRESS_VID_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h4,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_INGRESS_MST_TABLE;
                    ack.write_miss = handcode_error_INGRESS_MST_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b10??,8'h??,4'b??0?,1'b?},
           {32'b10??,8'h??,4'b??10,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_EGRESS_MST_TABLE;
                    ack.write_miss = handcode_error_EGRESS_MST_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'hC000,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_DIRECT_MAP_CTRL;
                    ack.write_miss = handcode_error_GLORT_DIRECT_MAP_CTRL;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'hC000,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_DIRECT_MAP_DST0;
                    ack.write_miss = handcode_error_GLORT_DIRECT_MAP_DST0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'hC001,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_DIRECT_MAP_DST1;
                    ack.write_miss = handcode_error_GLORT_DIRECT_MAP_DST1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'hC001,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_DIRECT_MAP_DST2;
                    ack.write_miss = handcode_error_GLORT_DIRECT_MAP_DST2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'hC002,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_DIRECT_MAP_DST3;
                    ack.write_miss = handcode_error_GLORT_DIRECT_MAP_DST3;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'hC002,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_DIRECT_MAP_DST4;
                    ack.write_miss = handcode_error_GLORT_DIRECT_MAP_DST4;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'hC0,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_RAM;
                    ack.write_miss = handcode_error_GLORT_RAM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'hC0,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_GLORT_CAM;
                    ack.write_miss = handcode_error_GLORT_CAM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'hC07,4'b011?,1'b?},
           {40'hC07,4'b1???,1'b?},
           {44'hC08?,1'b?},
           {40'hC09,4'b00??,1'b?},
           {40'hC09,4'b010?,1'b?},
           {44'hC096,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_CGRP_USED_TABLE;
                    ack.write_miss = handcode_error_CGRP_USED_TABLE;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_MST_GLORT_MAP_MEM) 
           {32'b0??,8'h??,4'b??0?,1'b?},
           {32'b0??,8'h??,4'b??10,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_EGRESS_VID_TABLE;
                 default: read_data = '0;
              endcase
           end
           {32'h4,4'b0???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_EGRESS_VID_CFG;
                 default: read_data = '0;
              endcase
           end
           {32'h4,4'b1???,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_INGRESS_MST_TABLE;
                 default: read_data = '0;
              endcase
           end
           {32'b10??,8'h??,4'b??0?,1'b?},
           {32'b10??,8'h??,4'b??10,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_EGRESS_MST_TABLE;
                 default: read_data = '0;
              endcase
           end
           {44'hC000,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_DIRECT_MAP_CTRL;
                 default: read_data = '0;
              endcase
           end
           {44'hC000,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_DIRECT_MAP_DST0;
                 default: read_data = '0;
              endcase
           end
           {44'hC001,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_DIRECT_MAP_DST1;
                 default: read_data = '0;
              endcase
           end
           {44'hC001,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_DIRECT_MAP_DST2;
                 default: read_data = '0;
              endcase
           end
           {44'hC002,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_DIRECT_MAP_DST3;
                 default: read_data = '0;
              endcase
           end
           {44'hC002,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_DIRECT_MAP_DST4;
                 default: read_data = '0;
              endcase
           end
           {36'hC0,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_RAM;
                 default: read_data = '0;
              endcase
           end
           {36'hC0,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_GLORT_CAM;
                 default: read_data = '0;
              endcase
           end
           {40'hC07,4'b011?,1'b?},
           {40'hC07,4'b1???,1'b?},
           {44'hC08?,1'b?},
           {40'hC09,4'b00??,1'b?},
           {40'hC09,4'b010?,1'b?},
           {44'hC096,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MST_GLORT_SB_FID,MST_GLORT_SB_BAR}: read_data = handcode_reg_rdata_CGRP_USED_TABLE;
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {


// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
