///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Jon Bagge <jon.bagge.com> 
// -- Project Name : MBY 
// -- Description  : classifier netlist. 
// ------------------------------------------------------------------- 

module classifier_top (
input reset, 
par_class_if.classifier par_class_if, 
//Input List
input                   cclk                                      
);

logic  [266:0] classifier_em_a_delay_fifo_0_from_mem;
logic  [285:0] classifier_em_a_delay_fifo_0_to_mem;
logic  [266:0] classifier_em_a_delay_fifo_1_from_mem;
logic  [285:0] classifier_em_a_delay_fifo_1_to_mem;
logic  [266:0] classifier_em_a_delay_fifo_2_from_mem;
logic  [285:0] classifier_em_a_delay_fifo_2_to_mem;
logic  [266:0] classifier_em_a_delay_fifo_3_from_mem;
logic  [285:0] classifier_em_a_delay_fifo_3_to_mem;
logic   [60:0] classifier_em_a_hash_cfg_from_mem;
logic   [79:0] classifier_em_a_hash_cfg_to_mem;
logic   [80:0] classifier_em_a_hash_lookup_from_mem;
logic  [104:0] classifier_em_a_hash_lookup_to_mem;
logic  [137:0] classifier_em_a_hash_miss_from_mem;
logic  [156:0] classifier_em_a_hash_miss_to_mem;
logic   [72:0] classifier_em_a_key_mask_0_from_mem;
logic   [91:0] classifier_em_a_key_mask_0_to_mem;
logic   [72:0] classifier_em_a_key_mask_1_from_mem;
logic   [91:0] classifier_em_a_key_mask_1_to_mem;
logic   [72:0] classifier_em_a_key_mask_2_from_mem;
logic   [91:0] classifier_em_a_key_mask_2_to_mem;
logic   [60:0] classifier_em_b_hash_cfg_from_mem;
logic   [79:0] classifier_em_b_hash_cfg_to_mem;
logic   [80:0] classifier_em_b_hash_lookup_from_mem;
logic  [101:0] classifier_em_b_hash_lookup_to_mem;
logic  [137:0] classifier_em_b_hash_miss_from_mem;
logic  [156:0] classifier_em_b_hash_miss_to_mem;
logic   [72:0] classifier_em_b_key_mask_from_mem;
logic   [91:0] classifier_em_b_key_mask_to_mem;
logic  [326:0] classifier_lpm_key_cam_from_tcam;
logic  [485:0] classifier_lpm_key_cam_to_tcam; 
logic  [306:0] classifier_lpm_tree_state_0_from_mem;
logic  [323:0] classifier_lpm_tree_state_0_to_mem;
logic  [306:0] classifier_lpm_tree_state_10_from_mem;
logic  [323:0] classifier_lpm_tree_state_10_to_mem;
logic  [306:0] classifier_lpm_tree_state_11_from_mem;
logic  [323:0] classifier_lpm_tree_state_11_to_mem;
logic  [306:0] classifier_lpm_tree_state_12_from_mem;
logic  [323:0] classifier_lpm_tree_state_12_to_mem;
logic  [306:0] classifier_lpm_tree_state_13_from_mem;
logic  [323:0] classifier_lpm_tree_state_13_to_mem;
logic  [306:0] classifier_lpm_tree_state_14_from_mem;
logic  [323:0] classifier_lpm_tree_state_14_to_mem;
logic  [306:0] classifier_lpm_tree_state_15_from_mem;
logic  [323:0] classifier_lpm_tree_state_15_to_mem;
logic  [306:0] classifier_lpm_tree_state_16_from_mem;
logic  [323:0] classifier_lpm_tree_state_16_to_mem;
logic  [306:0] classifier_lpm_tree_state_17_from_mem;
logic  [323:0] classifier_lpm_tree_state_17_to_mem;
logic  [306:0] classifier_lpm_tree_state_18_from_mem;
logic  [323:0] classifier_lpm_tree_state_18_to_mem;
logic  [306:0] classifier_lpm_tree_state_19_from_mem;
logic  [323:0] classifier_lpm_tree_state_19_to_mem;
logic  [306:0] classifier_lpm_tree_state_1_from_mem;
logic  [323:0] classifier_lpm_tree_state_1_to_mem;
logic  [306:0] classifier_lpm_tree_state_20_from_mem;
logic  [323:0] classifier_lpm_tree_state_20_to_mem;
logic  [306:0] classifier_lpm_tree_state_21_from_mem;
logic  [323:0] classifier_lpm_tree_state_21_to_mem;
logic  [306:0] classifier_lpm_tree_state_22_from_mem;
logic  [323:0] classifier_lpm_tree_state_22_to_mem;
logic  [306:0] classifier_lpm_tree_state_23_from_mem;
logic  [323:0] classifier_lpm_tree_state_23_to_mem;
logic  [306:0] classifier_lpm_tree_state_24_from_mem;
logic  [323:0] classifier_lpm_tree_state_24_to_mem;
logic  [306:0] classifier_lpm_tree_state_25_from_mem;
logic  [323:0] classifier_lpm_tree_state_25_to_mem;
logic  [306:0] classifier_lpm_tree_state_26_from_mem;
logic  [323:0] classifier_lpm_tree_state_26_to_mem;
logic  [306:0] classifier_lpm_tree_state_27_from_mem;
logic  [323:0] classifier_lpm_tree_state_27_to_mem;
logic  [306:0] classifier_lpm_tree_state_28_from_mem;
logic  [323:0] classifier_lpm_tree_state_28_to_mem;
logic  [306:0] classifier_lpm_tree_state_29_from_mem;
logic  [323:0] classifier_lpm_tree_state_29_to_mem;
logic  [306:0] classifier_lpm_tree_state_2_from_mem;
logic  [323:0] classifier_lpm_tree_state_2_to_mem;
logic  [306:0] classifier_lpm_tree_state_30_from_mem;
logic  [323:0] classifier_lpm_tree_state_30_to_mem;
logic  [306:0] classifier_lpm_tree_state_31_from_mem;
logic  [323:0] classifier_lpm_tree_state_31_to_mem;
logic  [306:0] classifier_lpm_tree_state_32_from_mem;
logic  [323:0] classifier_lpm_tree_state_32_to_mem;
logic  [306:0] classifier_lpm_tree_state_33_from_mem;
logic  [323:0] classifier_lpm_tree_state_33_to_mem;
logic  [306:0] classifier_lpm_tree_state_34_from_mem;
logic  [323:0] classifier_lpm_tree_state_34_to_mem;
logic  [306:0] classifier_lpm_tree_state_35_from_mem;
logic  [323:0] classifier_lpm_tree_state_35_to_mem;
logic  [306:0] classifier_lpm_tree_state_36_from_mem;
logic  [323:0] classifier_lpm_tree_state_36_to_mem;
logic  [306:0] classifier_lpm_tree_state_37_from_mem;
logic  [323:0] classifier_lpm_tree_state_37_to_mem;
logic  [306:0] classifier_lpm_tree_state_38_from_mem;
logic  [323:0] classifier_lpm_tree_state_38_to_mem;
logic  [306:0] classifier_lpm_tree_state_39_from_mem;
logic  [323:0] classifier_lpm_tree_state_39_to_mem;
logic  [306:0] classifier_lpm_tree_state_3_from_mem;
logic  [323:0] classifier_lpm_tree_state_3_to_mem;
logic  [306:0] classifier_lpm_tree_state_40_from_mem;
logic  [323:0] classifier_lpm_tree_state_40_to_mem;
logic  [306:0] classifier_lpm_tree_state_41_from_mem;
logic  [323:0] classifier_lpm_tree_state_41_to_mem;
logic  [306:0] classifier_lpm_tree_state_42_from_mem;
logic  [323:0] classifier_lpm_tree_state_42_to_mem;
logic  [306:0] classifier_lpm_tree_state_43_from_mem;
logic  [323:0] classifier_lpm_tree_state_43_to_mem;
logic  [306:0] classifier_lpm_tree_state_44_from_mem;
logic  [323:0] classifier_lpm_tree_state_44_to_mem;
logic  [306:0] classifier_lpm_tree_state_45_from_mem;
logic  [323:0] classifier_lpm_tree_state_45_to_mem;
logic  [306:0] classifier_lpm_tree_state_46_from_mem;
logic  [323:0] classifier_lpm_tree_state_46_to_mem;
logic  [306:0] classifier_lpm_tree_state_47_from_mem;
logic  [323:0] classifier_lpm_tree_state_47_to_mem;
logic  [306:0] classifier_lpm_tree_state_48_from_mem;
logic  [323:0] classifier_lpm_tree_state_48_to_mem;
logic  [306:0] classifier_lpm_tree_state_49_from_mem;
logic  [323:0] classifier_lpm_tree_state_49_to_mem;
logic  [306:0] classifier_lpm_tree_state_4_from_mem;
logic  [323:0] classifier_lpm_tree_state_4_to_mem;
logic  [306:0] classifier_lpm_tree_state_50_from_mem;
logic  [323:0] classifier_lpm_tree_state_50_to_mem;
logic  [306:0] classifier_lpm_tree_state_51_from_mem;
logic  [323:0] classifier_lpm_tree_state_51_to_mem;
logic  [306:0] classifier_lpm_tree_state_52_from_mem;
logic  [323:0] classifier_lpm_tree_state_52_to_mem;
logic  [306:0] classifier_lpm_tree_state_53_from_mem;
logic  [323:0] classifier_lpm_tree_state_53_to_mem;
logic  [306:0] classifier_lpm_tree_state_54_from_mem;
logic  [323:0] classifier_lpm_tree_state_54_to_mem;
logic  [306:0] classifier_lpm_tree_state_55_from_mem;
logic  [323:0] classifier_lpm_tree_state_55_to_mem;
logic  [306:0] classifier_lpm_tree_state_56_from_mem;
logic  [323:0] classifier_lpm_tree_state_56_to_mem;
logic  [306:0] classifier_lpm_tree_state_57_from_mem;
logic  [323:0] classifier_lpm_tree_state_57_to_mem;
logic  [306:0] classifier_lpm_tree_state_58_from_mem;
logic  [323:0] classifier_lpm_tree_state_58_to_mem;
logic  [306:0] classifier_lpm_tree_state_59_from_mem;
logic  [323:0] classifier_lpm_tree_state_59_to_mem;
logic  [306:0] classifier_lpm_tree_state_5_from_mem;
logic  [323:0] classifier_lpm_tree_state_5_to_mem;
logic  [306:0] classifier_lpm_tree_state_60_from_mem;
logic  [323:0] classifier_lpm_tree_state_60_to_mem;
logic  [306:0] classifier_lpm_tree_state_61_from_mem;
logic  [323:0] classifier_lpm_tree_state_61_to_mem;
logic  [306:0] classifier_lpm_tree_state_62_from_mem;
logic  [323:0] classifier_lpm_tree_state_62_to_mem;
logic  [306:0] classifier_lpm_tree_state_63_from_mem;
logic  [323:0] classifier_lpm_tree_state_63_to_mem;
logic  [306:0] classifier_lpm_tree_state_64_from_mem;
logic  [323:0] classifier_lpm_tree_state_64_to_mem;
logic  [306:0] classifier_lpm_tree_state_65_from_mem;
logic  [323:0] classifier_lpm_tree_state_65_to_mem;
logic  [306:0] classifier_lpm_tree_state_66_from_mem;
logic  [323:0] classifier_lpm_tree_state_66_to_mem;
logic  [306:0] classifier_lpm_tree_state_67_from_mem;
logic  [323:0] classifier_lpm_tree_state_67_to_mem;
logic  [306:0] classifier_lpm_tree_state_68_from_mem;
logic  [323:0] classifier_lpm_tree_state_68_to_mem;
logic  [306:0] classifier_lpm_tree_state_69_from_mem;
logic  [323:0] classifier_lpm_tree_state_69_to_mem;
logic  [306:0] classifier_lpm_tree_state_6_from_mem;
logic  [323:0] classifier_lpm_tree_state_6_to_mem;
logic  [306:0] classifier_lpm_tree_state_70_from_mem;
logic  [323:0] classifier_lpm_tree_state_70_to_mem;
logic  [306:0] classifier_lpm_tree_state_71_from_mem;
logic  [323:0] classifier_lpm_tree_state_71_to_mem;
logic  [306:0] classifier_lpm_tree_state_72_from_mem;
logic  [323:0] classifier_lpm_tree_state_72_to_mem;
logic  [306:0] classifier_lpm_tree_state_73_from_mem;
logic  [323:0] classifier_lpm_tree_state_73_to_mem;
logic  [306:0] classifier_lpm_tree_state_74_from_mem;
logic  [323:0] classifier_lpm_tree_state_74_to_mem;
logic  [306:0] classifier_lpm_tree_state_75_from_mem;
logic  [323:0] classifier_lpm_tree_state_75_to_mem;
logic  [306:0] classifier_lpm_tree_state_76_from_mem;
logic  [323:0] classifier_lpm_tree_state_76_to_mem;
logic  [306:0] classifier_lpm_tree_state_77_from_mem;
logic  [323:0] classifier_lpm_tree_state_77_to_mem;
logic  [306:0] classifier_lpm_tree_state_78_from_mem;
logic  [323:0] classifier_lpm_tree_state_78_to_mem;
logic  [306:0] classifier_lpm_tree_state_79_from_mem;
logic  [323:0] classifier_lpm_tree_state_79_to_mem;
logic  [306:0] classifier_lpm_tree_state_7_from_mem;
logic  [323:0] classifier_lpm_tree_state_7_to_mem;
logic  [306:0] classifier_lpm_tree_state_80_from_mem;
logic  [323:0] classifier_lpm_tree_state_80_to_mem;
logic  [306:0] classifier_lpm_tree_state_81_from_mem;
logic  [323:0] classifier_lpm_tree_state_81_to_mem;
logic  [306:0] classifier_lpm_tree_state_82_from_mem;
logic  [323:0] classifier_lpm_tree_state_82_to_mem;
logic  [306:0] classifier_lpm_tree_state_83_from_mem;
logic  [323:0] classifier_lpm_tree_state_83_to_mem;
logic  [306:0] classifier_lpm_tree_state_84_from_mem;
logic  [323:0] classifier_lpm_tree_state_84_to_mem;
logic  [306:0] classifier_lpm_tree_state_85_from_mem;
logic  [323:0] classifier_lpm_tree_state_85_to_mem;
logic  [306:0] classifier_lpm_tree_state_86_from_mem;
logic  [323:0] classifier_lpm_tree_state_86_to_mem;
logic  [306:0] classifier_lpm_tree_state_87_from_mem;
logic  [323:0] classifier_lpm_tree_state_87_to_mem;
logic  [306:0] classifier_lpm_tree_state_88_from_mem;
logic  [323:0] classifier_lpm_tree_state_88_to_mem;
logic  [306:0] classifier_lpm_tree_state_89_from_mem;
logic  [323:0] classifier_lpm_tree_state_89_to_mem;
logic  [306:0] classifier_lpm_tree_state_8_from_mem;
logic  [323:0] classifier_lpm_tree_state_8_to_mem;
logic  [306:0] classifier_lpm_tree_state_90_from_mem;
logic  [323:0] classifier_lpm_tree_state_90_to_mem;
logic  [306:0] classifier_lpm_tree_state_91_from_mem;
logic  [323:0] classifier_lpm_tree_state_91_to_mem;
logic  [306:0] classifier_lpm_tree_state_92_from_mem;
logic  [323:0] classifier_lpm_tree_state_92_to_mem;
logic  [306:0] classifier_lpm_tree_state_93_from_mem;
logic  [323:0] classifier_lpm_tree_state_93_to_mem;
logic  [306:0] classifier_lpm_tree_state_94_from_mem;
logic  [323:0] classifier_lpm_tree_state_94_to_mem;
logic  [306:0] classifier_lpm_tree_state_95_from_mem;
logic  [323:0] classifier_lpm_tree_state_95_to_mem;
logic  [306:0] classifier_lpm_tree_state_9_from_mem;
logic  [323:0] classifier_lpm_tree_state_9_to_mem;
logic   [72:0] classifier_map_domain_action0_from_mem;
logic   [92:0] classifier_map_domain_action0_to_mem;
logic   [72:0] classifier_map_domain_action1_from_mem;
logic   [92:0] classifier_map_domain_action1_to_mem;
logic   [72:0] classifier_map_domain_pol_cfg_from_mem;
logic   [81:0] classifier_map_domain_pol_cfg_to_mem;
logic   [72:0] classifier_map_domain_profile_from_mem;
logic   [89:0] classifier_map_domain_profile_to_mem;
logic [4181:0] classifier_map_domain_tcam_from_tcam;
logic [4434:0] classifier_map_domain_tcam_to_tcam;
logic   [72:0] classifier_map_dscp_tc_from_mem;
logic   [91:0] classifier_map_dscp_tc_to_mem;  
logic   [72:0] classifier_map_exp_tc_from_mem; 
logic   [89:0] classifier_map_exp_tc_to_mem;   
logic   [72:0] classifier_map_extract_0_from_mem;
logic   [87:0] classifier_map_extract_0_to_mem;
logic   [72:0] classifier_map_extract_1_from_mem;
logic   [87:0] classifier_map_extract_1_to_mem;
logic   [72:0] classifier_map_extract_2_from_mem;
logic   [87:0] classifier_map_extract_2_to_mem;
logic   [72:0] classifier_map_ip_cfg_from_mem; 
logic   [87:0] classifier_map_ip_cfg_to_mem;   
logic   [72:0] classifier_map_ip_hi_from_mem;  
logic   [87:0] classifier_map_ip_hi_to_mem;    
logic   [72:0] classifier_map_ip_lo_from_mem;  
logic   [87:0] classifier_map_ip_lo_to_mem;    
logic   [72:0] classifier_map_l4_dst_from_mem; 
logic   [86:0] classifier_map_l4_dst_to_mem;   
logic   [72:0] classifier_map_l4_src_from_mem; 
logic   [86:0] classifier_map_l4_src_to_mem;   
logic   [72:0] classifier_map_len_limit_from_mem;
logic   [91:0] classifier_map_len_limit_to_mem;
logic  [137:0] classifier_map_mac_from_mem;    
logic  [152:0] classifier_map_mac_to_mem;      
logic   [72:0] classifier_map_port_cfg_from_mem;
logic   [91:0] classifier_map_port_cfg_to_mem; 
logic   [72:0] classifier_map_port_default_0_from_mem;
logic   [85:0] classifier_map_port_default_0_to_mem;
logic   [72:0] classifier_map_port_default_10_from_mem;
logic   [85:0] classifier_map_port_default_10_to_mem;
logic   [72:0] classifier_map_port_default_11_from_mem;
logic   [85:0] classifier_map_port_default_11_to_mem;
logic   [72:0] classifier_map_port_default_12_from_mem;
logic   [85:0] classifier_map_port_default_12_to_mem;
logic   [72:0] classifier_map_port_default_13_from_mem;
logic   [85:0] classifier_map_port_default_13_to_mem;
logic   [72:0] classifier_map_port_default_14_from_mem;
logic   [85:0] classifier_map_port_default_14_to_mem;
logic   [72:0] classifier_map_port_default_15_from_mem;
logic   [85:0] classifier_map_port_default_15_to_mem;
logic   [72:0] classifier_map_port_default_16_from_mem;
logic   [85:0] classifier_map_port_default_16_to_mem;
logic   [72:0] classifier_map_port_default_17_from_mem;
logic   [85:0] classifier_map_port_default_17_to_mem;
logic   [72:0] classifier_map_port_default_18_from_mem;
logic   [85:0] classifier_map_port_default_18_to_mem;
logic   [72:0] classifier_map_port_default_19_from_mem;
logic   [85:0] classifier_map_port_default_19_to_mem;
logic   [72:0] classifier_map_port_default_1_from_mem;
logic   [85:0] classifier_map_port_default_1_to_mem;
logic   [72:0] classifier_map_port_default_20_from_mem;
logic   [85:0] classifier_map_port_default_20_to_mem;
logic   [72:0] classifier_map_port_default_21_from_mem;
logic   [85:0] classifier_map_port_default_21_to_mem;
logic   [72:0] classifier_map_port_default_22_from_mem;
logic   [85:0] classifier_map_port_default_22_to_mem;
logic   [72:0] classifier_map_port_default_23_from_mem;
logic   [85:0] classifier_map_port_default_23_to_mem;
logic   [72:0] classifier_map_port_default_24_from_mem;
logic   [85:0] classifier_map_port_default_24_to_mem;
logic   [72:0] classifier_map_port_default_25_from_mem;
logic   [85:0] classifier_map_port_default_25_to_mem;
logic   [72:0] classifier_map_port_default_26_from_mem;
logic   [85:0] classifier_map_port_default_26_to_mem;
logic   [72:0] classifier_map_port_default_27_from_mem;
logic   [85:0] classifier_map_port_default_27_to_mem;
logic   [72:0] classifier_map_port_default_28_from_mem;
logic   [85:0] classifier_map_port_default_28_to_mem;
logic   [72:0] classifier_map_port_default_29_from_mem;
logic   [85:0] classifier_map_port_default_29_to_mem;
logic   [72:0] classifier_map_port_default_2_from_mem;
logic   [85:0] classifier_map_port_default_2_to_mem;
logic   [72:0] classifier_map_port_default_30_from_mem;
logic   [85:0] classifier_map_port_default_30_to_mem;
logic   [72:0] classifier_map_port_default_31_from_mem;
logic   [85:0] classifier_map_port_default_31_to_mem;
logic   [72:0] classifier_map_port_default_32_from_mem;
logic   [85:0] classifier_map_port_default_32_to_mem;
logic   [72:0] classifier_map_port_default_3_from_mem;
logic   [85:0] classifier_map_port_default_3_to_mem;
logic   [72:0] classifier_map_port_default_4_from_mem;
logic   [85:0] classifier_map_port_default_4_to_mem;
logic   [72:0] classifier_map_port_default_5_from_mem;
logic   [85:0] classifier_map_port_default_5_to_mem;
logic   [72:0] classifier_map_port_default_6_from_mem;
logic   [85:0] classifier_map_port_default_6_to_mem;
logic   [72:0] classifier_map_port_default_7_from_mem;
logic   [85:0] classifier_map_port_default_7_to_mem;
logic   [72:0] classifier_map_port_default_8_from_mem;
logic   [85:0] classifier_map_port_default_8_to_mem;
logic   [72:0] classifier_map_port_default_9_from_mem;
logic   [85:0] classifier_map_port_default_9_to_mem;
logic   [72:0] classifier_map_port_from_mem;   
logic   [91:0] classifier_map_port_to_mem;     
logic   [72:0] classifier_map_profile_action_from_mem;
logic   [87:0] classifier_map_profile_action_to_mem;
logic   [88:0] classifier_map_profile_key0_from_mem;
logic  [109:0] classifier_map_profile_key0_to_mem;
logic   [88:0] classifier_map_profile_key1_from_mem;
logic  [109:0] classifier_map_profile_key1_to_mem;
logic   [88:0] classifier_map_profile_key_invert0_from_mem;
logic  [109:0] classifier_map_profile_key_invert0_to_mem;
logic   [88:0] classifier_map_profile_key_invert1_from_mem;
logic  [109:0] classifier_map_profile_key_invert1_to_mem;
logic   [72:0] classifier_map_prot_from_mem;   
logic   [85:0] classifier_map_prot_to_mem;     
logic   [72:0] classifier_map_rewrite_0_from_mem;
logic   [89:0] classifier_map_rewrite_0_to_mem;
logic   [72:0] classifier_map_rewrite_10_from_mem;
logic   [89:0] classifier_map_rewrite_10_to_mem;
logic   [72:0] classifier_map_rewrite_11_from_mem;
logic   [89:0] classifier_map_rewrite_11_to_mem;
logic   [72:0] classifier_map_rewrite_12_from_mem;
logic   [89:0] classifier_map_rewrite_12_to_mem;
logic   [72:0] classifier_map_rewrite_13_from_mem;
logic   [89:0] classifier_map_rewrite_13_to_mem;
logic   [72:0] classifier_map_rewrite_14_from_mem;
logic   [89:0] classifier_map_rewrite_14_to_mem;
logic   [72:0] classifier_map_rewrite_15_from_mem;
logic   [89:0] classifier_map_rewrite_15_to_mem;
logic   [72:0] classifier_map_rewrite_1_from_mem;
logic   [89:0] classifier_map_rewrite_1_to_mem;
logic   [72:0] classifier_map_rewrite_2_from_mem;
logic   [89:0] classifier_map_rewrite_2_to_mem;
logic   [72:0] classifier_map_rewrite_3_from_mem;
logic   [89:0] classifier_map_rewrite_3_to_mem;
logic   [72:0] classifier_map_rewrite_4_from_mem;
logic   [89:0] classifier_map_rewrite_4_to_mem;
logic   [72:0] classifier_map_rewrite_5_from_mem;
logic   [89:0] classifier_map_rewrite_5_to_mem;
logic   [72:0] classifier_map_rewrite_6_from_mem;
logic   [89:0] classifier_map_rewrite_6_to_mem;
logic   [72:0] classifier_map_rewrite_7_from_mem;
logic   [89:0] classifier_map_rewrite_7_to_mem;
logic   [72:0] classifier_map_rewrite_8_from_mem;
logic   [89:0] classifier_map_rewrite_8_to_mem;
logic   [72:0] classifier_map_rewrite_9_from_mem;
logic   [89:0] classifier_map_rewrite_9_to_mem;
logic   [72:0] classifier_map_type_from_mem;   
logic   [87:0] classifier_map_type_to_mem;     
logic   [72:0] classifier_map_vpri_from_mem;   
logic   [72:0] classifier_map_vpri_tc_from_mem;
logic   [89:0] classifier_map_vpri_tc_to_mem;  
logic   [89:0] classifier_map_vpri_to_mem;     
logic   [68:0] classifier_wcm_action_cfg_0_from_mem;
logic   [88:0] classifier_wcm_action_cfg_0_to_mem;
logic   [68:0] classifier_wcm_action_cfg_1_from_mem;
logic   [88:0] classifier_wcm_action_cfg_1_to_mem;
logic   [72:0] classifier_wcm_action_ram_0_from_mem;
logic   [90:0] classifier_wcm_action_ram_0_to_mem;
logic   [72:0] classifier_wcm_action_ram_10_from_mem;
logic   [90:0] classifier_wcm_action_ram_10_to_mem;
logic   [72:0] classifier_wcm_action_ram_11_from_mem;
logic   [90:0] classifier_wcm_action_ram_11_to_mem;
logic   [72:0] classifier_wcm_action_ram_12_from_mem;
logic   [90:0] classifier_wcm_action_ram_12_to_mem;
logic   [72:0] classifier_wcm_action_ram_13_from_mem;
logic   [90:0] classifier_wcm_action_ram_13_to_mem;
logic   [72:0] classifier_wcm_action_ram_14_from_mem;
logic   [90:0] classifier_wcm_action_ram_14_to_mem;
logic   [72:0] classifier_wcm_action_ram_15_from_mem;
logic   [90:0] classifier_wcm_action_ram_15_to_mem;
logic   [72:0] classifier_wcm_action_ram_16_from_mem;
logic   [90:0] classifier_wcm_action_ram_16_to_mem;
logic   [72:0] classifier_wcm_action_ram_17_from_mem;
logic   [90:0] classifier_wcm_action_ram_17_to_mem;
logic   [72:0] classifier_wcm_action_ram_18_from_mem;
logic   [90:0] classifier_wcm_action_ram_18_to_mem;
logic   [72:0] classifier_wcm_action_ram_19_from_mem;
logic   [90:0] classifier_wcm_action_ram_19_to_mem;
logic   [72:0] classifier_wcm_action_ram_1_from_mem;
logic   [90:0] classifier_wcm_action_ram_1_to_mem;
logic   [72:0] classifier_wcm_action_ram_20_from_mem;
logic   [90:0] classifier_wcm_action_ram_20_to_mem;
logic   [72:0] classifier_wcm_action_ram_21_from_mem;
logic   [90:0] classifier_wcm_action_ram_21_to_mem;
logic   [72:0] classifier_wcm_action_ram_22_from_mem;
logic   [90:0] classifier_wcm_action_ram_22_to_mem;
logic   [72:0] classifier_wcm_action_ram_23_from_mem;
logic   [90:0] classifier_wcm_action_ram_23_to_mem;
logic   [72:0] classifier_wcm_action_ram_2_from_mem;
logic   [90:0] classifier_wcm_action_ram_2_to_mem;
logic   [72:0] classifier_wcm_action_ram_3_from_mem;
logic   [90:0] classifier_wcm_action_ram_3_to_mem;
logic   [72:0] classifier_wcm_action_ram_4_from_mem;
logic   [90:0] classifier_wcm_action_ram_4_to_mem;
logic   [72:0] classifier_wcm_action_ram_5_from_mem;
logic   [90:0] classifier_wcm_action_ram_5_to_mem;
logic   [72:0] classifier_wcm_action_ram_6_from_mem;
logic   [90:0] classifier_wcm_action_ram_6_to_mem;
logic   [72:0] classifier_wcm_action_ram_7_from_mem;
logic   [90:0] classifier_wcm_action_ram_7_to_mem;
logic   [72:0] classifier_wcm_action_ram_8_from_mem;
logic   [90:0] classifier_wcm_action_ram_8_to_mem;
logic   [72:0] classifier_wcm_action_ram_9_from_mem;
logic   [90:0] classifier_wcm_action_ram_9_to_mem;
logic   [72:0] classifier_wcm_data_path_buffer0_from_mem;
logic   [85:0] classifier_wcm_data_path_buffer0_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_0_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_0_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_10_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_10_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_11_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_11_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_12_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_12_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_13_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_13_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_14_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_14_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_15_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_15_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_16_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_16_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_17_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_17_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_18_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_18_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_19_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_19_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_1_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_1_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_2_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_2_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_3_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_3_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_4_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_4_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_5_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_5_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_6_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_6_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_7_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_7_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_8_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_8_to_mem;
logic  [345:0] classifier_wcm_data_path_buffer1_9_from_mem;
logic  [362:0] classifier_wcm_data_path_buffer1_9_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_0_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_0_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_10_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_10_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_11_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_11_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_12_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_12_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_13_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_13_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_14_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_14_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_15_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_15_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_16_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_16_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_17_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_17_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_18_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_18_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_19_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_19_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_1_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_1_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_2_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_2_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_3_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_3_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_4_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_4_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_5_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_5_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_6_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_6_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_7_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_7_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_8_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_8_to_mem;
logic   [70:0] classifier_wcm_tcam_cfg_ram_9_from_mem;
logic   [88:0] classifier_wcm_tcam_cfg_ram_9_to_mem;
logic reset_n; 
assign reset_n = !reset;


// module classifier_shells_wrapper    from classifier_shells_wrapper using classifier_shells_wrapper.map 
classifier_shells_wrapper    classifier_shells_wrapper(
/* input  logic           */ .LPM_TREE_STATE_32_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_32_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_33_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_33_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_34_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_34_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_35_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_35_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_36_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_36_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_37_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_37_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_38_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_38_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_39_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_39_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_3_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_3_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_40_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_40_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_41_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_41_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_42_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_42_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_43_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_43_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_44_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_44_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_45_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_45_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_46_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_46_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_47_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_47_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_48_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_48_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_49_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_49_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_4_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_4_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_50_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_50_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_51_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_51_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_52_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_52_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_53_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_53_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_54_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_54_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_55_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_55_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_56_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_56_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_57_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_57_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_58_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_58_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_59_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_59_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_5_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_61_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_62_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_62_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_63_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_63_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_64_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_64_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_65_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_65_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_66_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_66_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_67_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_67_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_68_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_68_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_69_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_69_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_6_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_6_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_70_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_70_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_71_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_71_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_72_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_72_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_73_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_73_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_74_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_74_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_75_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_75_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_76_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_76_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_77_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_77_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_78_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_78_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_79_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_79_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_7_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_7_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_80_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_80_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_81_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_81_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_82_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_82_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_83_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_83_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_84_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_84_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_85_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_85_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_86_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_86_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_87_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_87_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_88_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_88_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_89_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_89_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_8_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_8_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_90_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_90_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_91_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_91_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_92_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_92_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_93_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_93_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_94_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_94_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_95_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_95_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_9_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_9_STATUS_reg_sel              (),                                           
/* input  logic           */ .MAP_DOMAIN_ACTION0_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_DOMAIN_ACTION0_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_DOMAIN_ACTION1_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_DOMAIN_ACTION1_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_DOMAIN_TCAM_CFG_reg_sel                  (),                                           
/* input  logic           */ .MAP_DOMAIN_TCAM_STATUS_reg_sel               (),                                           
/* input  logic           */ .MAP_DSCP_TC_CFG_reg_sel                      (),                                           
/* input  logic           */ .MAP_DSCP_TC_STATUS_reg_sel                   (),                                           
/* input  logic           */ .MAP_EXP_TC_CFG_reg_sel                       (),                                           
/* input  logic           */ .MAP_EXP_TC_STATUS_reg_sel                    (),                                           
/* input  logic           */ .MAP_EXTRACT_0_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_EXTRACT_0_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_EXTRACT_1_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_EXTRACT_1_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_EXTRACT_2_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_EXTRACT_2_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_IP_CFG_CFG_reg_sel                       (),                                           
/* input  logic           */ .MAP_IP_CFG_STATUS_reg_sel                    (),                                           
/* input  logic           */ .MAP_IP_HI_CFG_reg_sel                        (),                                           
/* input  logic           */ .MAP_IP_HI_STATUS_reg_sel                     (),                                           
/* input  logic           */ .MAP_IP_LO_CFG_reg_sel                        (),                                           
/* input  logic           */ .MAP_IP_LO_STATUS_reg_sel                     (),                                           
/* input  logic           */ .MAP_L4_DST_CFG_reg_sel                       (),                                           
/* input  logic           */ .MAP_L4_DST_STATUS_reg_sel                    (),                                           
/* input  logic           */ .MAP_L4_SRC_CFG_reg_sel                       (),                                           
/* input  logic           */ .MAP_L4_SRC_STATUS_reg_sel                    (),                                           
/* input  logic           */ .MAP_LEN_LIMIT_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_LEN_LIMIT_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_MAC_CFG_reg_sel                          (),                                           
/* input  logic           */ .MAP_MAC_STATUS_reg_sel                       (),                                           
/* input  logic           */ .MAP_PORT_CFG_CFG_reg_sel                     (),                                           
/* input  logic           */ .MAP_PORT_CFG_STATUS_reg_sel                  (),                                           
/* input  logic           */ .MAP_PORT_CFG_reg_sel                         (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_0_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_0_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_10_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_10_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_11_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_11_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_12_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_12_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_13_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_13_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_14_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_14_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_15_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_15_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_16_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_16_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_17_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_17_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_18_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_18_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_19_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_19_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_1_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_1_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_20_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_20_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_21_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_21_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_22_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_22_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_23_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_23_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_24_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_24_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_25_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_25_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_26_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_26_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_27_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_27_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_28_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_28_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_29_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_29_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_2_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_2_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_30_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_30_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_31_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_31_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_32_CFG_reg_sel              (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_32_STATUS_reg_sel           (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_3_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_3_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_4_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_6_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_7_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_7_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_8_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_8_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_9_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_9_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_STATUS_reg_sel                      (),                                           
/* input  logic           */ .MAP_PROFILE_ACTION_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PROFILE_ACTION_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PROFILE_KEY0_CFG_reg_sel                 (),                                           
/* input  logic           */ .MAP_PROFILE_KEY0_STATUS_reg_sel              (),                                           
/* input  logic           */ .MAP_PROFILE_KEY1_CFG_reg_sel                 (),                                           
/* input  logic           */ .MAP_PROFILE_KEY1_STATUS_reg_sel              (),                                           
/* input  logic           */ .MAP_PROFILE_KEY_INVERT0_CFG_reg_sel          (),                                           
/* input  logic           */ .MAP_PROFILE_KEY_INVERT0_STATUS_reg_sel       (),                                           
/* input  logic           */ .MAP_PROFILE_KEY_INVERT1_CFG_reg_sel          (),                                           
/* input  logic           */ .MAP_PROFILE_KEY_INVERT1_STATUS_reg_sel       (),                                           
/* input  logic           */ .MAP_PROT_CFG_reg_sel                         (),                                           
/* input  logic           */ .MAP_PROT_STATUS_reg_sel                      (),                                           
/* input  logic           */ .MAP_REWRITE_0_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_0_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_10_CFG_reg_sel                   (),                                           
/* input  logic           */ .MAP_REWRITE_10_STATUS_reg_sel                (),                                           
/* input  logic           */ .MAP_REWRITE_11_CFG_reg_sel                   (),                                           
/* input  logic           */ .MAP_REWRITE_11_STATUS_reg_sel                (),                                           
/* input  logic           */ .MAP_REWRITE_12_CFG_reg_sel                   (),                                           
/* input  logic           */ .MAP_REWRITE_12_STATUS_reg_sel                (),                                           
/* input  logic           */ .MAP_REWRITE_13_CFG_reg_sel                   (),                                           
/* input  logic           */ .MAP_REWRITE_13_STATUS_reg_sel                (),                                           
/* input  logic           */ .MAP_REWRITE_14_CFG_reg_sel                   (),                                           
/* input  logic           */ .MAP_REWRITE_14_STATUS_reg_sel                (),                                           
/* input  logic           */ .MAP_REWRITE_15_CFG_reg_sel                   (),                                           
/* input  logic           */ .MAP_REWRITE_15_STATUS_reg_sel                (),                                           
/* input  logic           */ .MAP_REWRITE_1_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_1_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_2_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_2_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_3_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_3_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_4_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_4_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_5_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_5_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_6_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_6_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_7_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_7_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_8_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_8_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_REWRITE_9_CFG_reg_sel                    (),                                           
/* input  logic           */ .MAP_REWRITE_9_STATUS_reg_sel                 (),                                           
/* input  logic           */ .MAP_TYPE_CFG_reg_sel                         (),                                           
/* input  logic           */ .MAP_TYPE_STATUS_reg_sel                      (),                                           
/* input  logic           */ .MAP_VPRI_CFG_reg_sel                         (),                                           
/* input  logic           */ .MAP_VPRI_STATUS_reg_sel                      (),                                           
/* input  logic           */ .MAP_VPRI_TC_CFG_reg_sel                      (),                                           
/* input  logic           */ .MAP_VPRI_TC_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_ACTION_CFG_0_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_CFG_0_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_CFG_1_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_CFG_1_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_0_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_0_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_10_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_10_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_11_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_11_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_12_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_12_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_13_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_13_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_14_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_14_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_15_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_15_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_16_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_16_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_17_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_17_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_18_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_1_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_20_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_20_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_21_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_21_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_22_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_22_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_23_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_23_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_2_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_2_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_3_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_3_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_4_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_4_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_5_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_5_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_6_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_6_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_7_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_7_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_8_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_8_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_ACTION_RAM_9_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_ACTION_RAM_9_STATUS_reg_sel              (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER0_CFG_reg_sel            (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER0_STATUS_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_0_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_0_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_10_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_10_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_11_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_11_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_12_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_12_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_13_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_13_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_14_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_14_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_15_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_15_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_16_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_16_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_17_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_17_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_18_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_18_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_19_CFG_reg_sel         (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_19_STATUS_reg_sel      (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_1_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_1_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_2_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_2_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_3_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_3_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_4_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_4_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_5_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_5_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_6_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_6_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_7_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_7_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_8_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_8_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_9_CFG_reg_sel          (),                                           
/* input  logic           */ .WCM_DATA_PATH_BUFFER1_9_STATUS_reg_sel       (),                                           
/* input  logic           */ .WCM_TCAM_0_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_0_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_10_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_10_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_11_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_11_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_12_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_12_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_13_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_13_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_14_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_14_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_15_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_17_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_18_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_18_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_19_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_19_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_1_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_1_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_2_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_2_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_3_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_3_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_4_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_4_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_5_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_5_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_6_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_6_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_7_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_7_STATUS_reg_sel                    (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_30_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_30_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_31_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_31_mem_ls_enter               (),                                           
/* input  logic           */ .WCM_TCAM_8_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_8_STATUS_reg_sel                    (),                                           
/* input  logic           */ .WCM_TCAM_9_CFG_reg_sel                       (),                                           
/* input  logic           */ .WCM_TCAM_9_STATUS_reg_sel                    (),                                           
/* input  logic           */ .lpm_tree_state_32_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_32_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_32_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_32_wr_en                      (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_0_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_0_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_10_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_10_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_11_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_11_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_12_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_12_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_13_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_13_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_14_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_14_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_15_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_15_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_16_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_16_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_17_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_17_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_18_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_18_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_19_CFG_reg_sel              (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_19_STATUS_reg_sel           (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_1_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_1_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_2_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_2_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_3_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_3_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_4_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_4_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_5_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_5_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_6_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_6_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_7_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_7_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_8_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_8_STATUS_reg_sel            (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_9_CFG_reg_sel               (),                                           
/* input  logic           */ .WCM_TCAM_CFG_RAM_9_STATUS_reg_sel            (),                                           
/* input  logic   [266:0] */ .classifier_em_a_delay_fifo_0_from_mem        (classifier_em_a_delay_fifo_0_from_mem),      
/* input  logic   [266:0] */ .classifier_em_a_delay_fifo_1_from_mem        (classifier_em_a_delay_fifo_1_from_mem),      
/* input  logic   [266:0] */ .classifier_em_a_delay_fifo_2_from_mem        (classifier_em_a_delay_fifo_2_from_mem),      
/* input  logic   [266:0] */ .classifier_em_a_delay_fifo_3_from_mem        (classifier_em_a_delay_fifo_3_from_mem),      
/* input  logic    [60:0] */ .classifier_em_a_hash_cfg_from_mem            (classifier_em_a_hash_cfg_from_mem),          
/* input  logic    [80:0] */ .classifier_em_a_hash_lookup_from_mem         (classifier_em_a_hash_lookup_from_mem),       
/* input  logic   [137:0] */ .classifier_em_a_hash_miss_from_mem           (classifier_em_a_hash_miss_from_mem),         
/* input  logic    [72:0] */ .classifier_em_a_key_mask_0_from_mem          (classifier_em_a_key_mask_0_from_mem),        
/* input  logic    [72:0] */ .classifier_em_a_key_mask_1_from_mem          (classifier_em_a_key_mask_1_from_mem),        
/* input  logic    [72:0] */ .classifier_em_a_key_mask_2_from_mem          (classifier_em_a_key_mask_2_from_mem),        
/* input  logic    [60:0] */ .classifier_em_b_hash_cfg_from_mem            (classifier_em_b_hash_cfg_from_mem),          
/* input  logic    [80:0] */ .classifier_em_b_hash_lookup_from_mem         (classifier_em_b_hash_lookup_from_mem),       
/* input  logic   [137:0] */ .classifier_em_b_hash_miss_from_mem           (classifier_em_b_hash_miss_from_mem),         
/* input  logic    [72:0] */ .classifier_em_b_key_mask_from_mem            (classifier_em_b_key_mask_from_mem),          
/* input  logic   [326:0] */ .classifier_lpm_key_cam_from_tcam             (classifier_lpm_key_cam_from_tcam),           
/* input  logic   [306:0] */ .classifier_lpm_tree_state_0_from_mem         (classifier_lpm_tree_state_0_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_10_from_mem        (classifier_lpm_tree_state_10_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_11_from_mem        (classifier_lpm_tree_state_11_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_12_from_mem        (classifier_lpm_tree_state_12_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_13_from_mem        (classifier_lpm_tree_state_13_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_14_from_mem        (classifier_lpm_tree_state_14_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_15_from_mem        (classifier_lpm_tree_state_15_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_16_from_mem        (classifier_lpm_tree_state_16_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_17_from_mem        (classifier_lpm_tree_state_17_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_18_from_mem        (classifier_lpm_tree_state_18_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_19_from_mem        (classifier_lpm_tree_state_19_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_1_from_mem         (classifier_lpm_tree_state_1_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_20_from_mem        (classifier_lpm_tree_state_20_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_21_from_mem        (classifier_lpm_tree_state_21_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_26_from_mem        (classifier_lpm_tree_state_26_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_27_from_mem        (classifier_lpm_tree_state_27_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_28_from_mem        (classifier_lpm_tree_state_28_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_29_from_mem        (classifier_lpm_tree_state_29_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_2_from_mem         (classifier_lpm_tree_state_2_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_30_from_mem        (classifier_lpm_tree_state_30_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_31_from_mem        (classifier_lpm_tree_state_31_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_32_from_mem        (classifier_lpm_tree_state_32_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_33_from_mem        (classifier_lpm_tree_state_33_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_34_from_mem        (classifier_lpm_tree_state_34_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_35_from_mem        (classifier_lpm_tree_state_35_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_36_from_mem        (classifier_lpm_tree_state_36_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_37_from_mem        (classifier_lpm_tree_state_37_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_38_from_mem        (classifier_lpm_tree_state_38_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_39_from_mem        (classifier_lpm_tree_state_39_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_3_from_mem         (classifier_lpm_tree_state_3_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_40_from_mem        (classifier_lpm_tree_state_40_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_41_from_mem        (classifier_lpm_tree_state_41_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_42_from_mem        (classifier_lpm_tree_state_42_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_43_from_mem        (classifier_lpm_tree_state_43_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_44_from_mem        (classifier_lpm_tree_state_44_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_45_from_mem        (classifier_lpm_tree_state_45_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_46_from_mem        (classifier_lpm_tree_state_46_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_47_from_mem        (classifier_lpm_tree_state_47_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_48_from_mem        (classifier_lpm_tree_state_48_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_49_from_mem        (classifier_lpm_tree_state_49_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_4_from_mem         (classifier_lpm_tree_state_4_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_50_from_mem        (classifier_lpm_tree_state_50_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_51_from_mem        (classifier_lpm_tree_state_51_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_52_from_mem        (classifier_lpm_tree_state_52_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_53_from_mem        (classifier_lpm_tree_state_53_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_54_from_mem        (classifier_lpm_tree_state_54_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_55_from_mem        (classifier_lpm_tree_state_55_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_56_from_mem        (classifier_lpm_tree_state_56_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_57_from_mem        (classifier_lpm_tree_state_57_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_58_from_mem        (classifier_lpm_tree_state_58_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_59_from_mem        (classifier_lpm_tree_state_59_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_5_from_mem         (classifier_lpm_tree_state_5_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_60_from_mem        (classifier_lpm_tree_state_60_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_61_from_mem        (classifier_lpm_tree_state_61_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_62_from_mem        (classifier_lpm_tree_state_62_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_63_from_mem        (classifier_lpm_tree_state_63_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_64_from_mem        (classifier_lpm_tree_state_64_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_65_from_mem        (classifier_lpm_tree_state_65_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_66_from_mem        (classifier_lpm_tree_state_66_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_67_from_mem        (classifier_lpm_tree_state_67_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_68_from_mem        (classifier_lpm_tree_state_68_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_69_from_mem        (classifier_lpm_tree_state_69_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_6_from_mem         (classifier_lpm_tree_state_6_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_70_from_mem        (classifier_lpm_tree_state_70_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_71_from_mem        (classifier_lpm_tree_state_71_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_72_from_mem        (classifier_lpm_tree_state_72_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_73_from_mem        (classifier_lpm_tree_state_73_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_74_from_mem        (classifier_lpm_tree_state_74_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_75_from_mem        (classifier_lpm_tree_state_75_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_76_from_mem        (classifier_lpm_tree_state_76_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_77_from_mem        (classifier_lpm_tree_state_77_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_78_from_mem        (classifier_lpm_tree_state_78_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_79_from_mem        (classifier_lpm_tree_state_79_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_7_from_mem         (classifier_lpm_tree_state_7_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_80_from_mem        (classifier_lpm_tree_state_80_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_81_from_mem        (classifier_lpm_tree_state_81_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_82_from_mem        (classifier_lpm_tree_state_82_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_83_from_mem        (classifier_lpm_tree_state_83_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_84_from_mem        (classifier_lpm_tree_state_84_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_85_from_mem        (classifier_lpm_tree_state_85_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_86_from_mem        (classifier_lpm_tree_state_86_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_87_from_mem        (classifier_lpm_tree_state_87_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_88_from_mem        (classifier_lpm_tree_state_88_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_89_from_mem        (classifier_lpm_tree_state_89_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_8_from_mem         (classifier_lpm_tree_state_8_from_mem),       
/* input  logic   [306:0] */ .classifier_lpm_tree_state_90_from_mem        (classifier_lpm_tree_state_90_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_91_from_mem        (classifier_lpm_tree_state_91_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_92_from_mem        (classifier_lpm_tree_state_92_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_93_from_mem        (classifier_lpm_tree_state_93_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_94_from_mem        (classifier_lpm_tree_state_94_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_95_from_mem        (classifier_lpm_tree_state_95_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_9_from_mem         (classifier_lpm_tree_state_9_from_mem),       
/* input  logic    [72:0] */ .classifier_map_domain_action0_from_mem       (classifier_map_domain_action0_from_mem),     
/* input  logic    [72:0] */ .classifier_map_domain_action1_from_mem       (classifier_map_domain_action1_from_mem),     
/* input  logic    [72:0] */ .classifier_map_domain_pol_cfg_from_mem       (classifier_map_domain_pol_cfg_from_mem),     
/* input  logic    [72:0] */ .classifier_map_domain_profile_from_mem       (classifier_map_domain_profile_from_mem),     
/* input  logic  [4181:0] */ .classifier_map_domain_tcam_from_tcam         (classifier_map_domain_tcam_from_tcam),       
/* input  logic    [72:0] */ .classifier_map_dscp_tc_from_mem              (classifier_map_dscp_tc_from_mem),            
/* input  logic    [72:0] */ .classifier_map_exp_tc_from_mem               (classifier_map_exp_tc_from_mem),             
/* input  logic    [72:0] */ .classifier_map_extract_0_from_mem            (classifier_map_extract_0_from_mem),          
/* input  logic    [72:0] */ .classifier_map_extract_1_from_mem            (classifier_map_extract_1_from_mem),          
/* input  logic    [72:0] */ .classifier_map_extract_2_from_mem            (classifier_map_extract_2_from_mem),          
/* input  logic    [72:0] */ .classifier_map_ip_cfg_from_mem               (classifier_map_ip_cfg_from_mem),             
/* input  logic    [72:0] */ .classifier_map_ip_hi_from_mem                (classifier_map_ip_hi_from_mem),              
/* input  logic    [72:0] */ .classifier_map_ip_lo_from_mem                (classifier_map_ip_lo_from_mem),              
/* input  logic    [72:0] */ .classifier_map_l4_dst_from_mem               (classifier_map_l4_dst_from_mem),             
/* input  logic    [72:0] */ .classifier_map_l4_src_from_mem               (classifier_map_l4_src_from_mem),             
/* input  logic    [72:0] */ .classifier_map_len_limit_from_mem            (classifier_map_len_limit_from_mem),          
/* input  logic   [137:0] */ .classifier_map_mac_from_mem                  (classifier_map_mac_from_mem),                
/* input  logic    [72:0] */ .classifier_map_port_cfg_from_mem             (classifier_map_port_cfg_from_mem),           
/* input  logic    [72:0] */ .classifier_map_port_default_0_from_mem       (classifier_map_port_default_0_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_10_from_mem      (classifier_map_port_default_10_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_11_from_mem      (classifier_map_port_default_11_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_12_from_mem      (classifier_map_port_default_12_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_13_from_mem      (classifier_map_port_default_13_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_14_from_mem      (classifier_map_port_default_14_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_15_from_mem      (classifier_map_port_default_15_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_16_from_mem      (classifier_map_port_default_16_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_17_from_mem      (classifier_map_port_default_17_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_18_from_mem      (classifier_map_port_default_18_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_19_from_mem      (classifier_map_port_default_19_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_1_from_mem       (classifier_map_port_default_1_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_20_from_mem      (classifier_map_port_default_20_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_21_from_mem      (classifier_map_port_default_21_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_22_from_mem      (classifier_map_port_default_22_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_23_from_mem      (classifier_map_port_default_23_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_24_from_mem      (classifier_map_port_default_24_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_25_from_mem      (classifier_map_port_default_25_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_26_from_mem      (classifier_map_port_default_26_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_27_from_mem      (classifier_map_port_default_27_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_28_from_mem      (classifier_map_port_default_28_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_29_from_mem      (classifier_map_port_default_29_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_2_from_mem       (classifier_map_port_default_2_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_4_from_mem       (classifier_map_port_default_4_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_5_from_mem       (classifier_map_port_default_5_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_6_from_mem       (classifier_map_port_default_6_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_7_from_mem       (classifier_map_port_default_7_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_8_from_mem       (classifier_map_port_default_8_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_default_9_from_mem       (classifier_map_port_default_9_from_mem),     
/* input  logic    [72:0] */ .classifier_map_port_from_mem                 (classifier_map_port_from_mem),               
/* input  logic    [72:0] */ .classifier_map_profile_action_from_mem       (classifier_map_profile_action_from_mem),     
/* input  logic    [88:0] */ .classifier_map_profile_key0_from_mem         (classifier_map_profile_key0_from_mem),       
/* input  logic    [88:0] */ .classifier_map_profile_key1_from_mem         (classifier_map_profile_key1_from_mem),       
/* input  logic    [88:0] */ .classifier_map_profile_key_invert0_from_mem  (classifier_map_profile_key_invert0_from_mem), 
/* input  logic    [88:0] */ .classifier_map_profile_key_invert1_from_mem  (classifier_map_profile_key_invert1_from_mem), 
/* input  logic    [72:0] */ .classifier_map_prot_from_mem                 (classifier_map_prot_from_mem),               
/* input  logic    [72:0] */ .classifier_map_rewrite_0_from_mem            (classifier_map_rewrite_0_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_10_from_mem           (classifier_map_rewrite_10_from_mem),         
/* input  logic    [72:0] */ .classifier_map_rewrite_11_from_mem           (classifier_map_rewrite_11_from_mem),         
/* input  logic    [72:0] */ .classifier_map_rewrite_12_from_mem           (classifier_map_rewrite_12_from_mem),         
/* input  logic    [72:0] */ .classifier_map_rewrite_13_from_mem           (classifier_map_rewrite_13_from_mem),         
/* input  logic    [72:0] */ .classifier_map_rewrite_14_from_mem           (classifier_map_rewrite_14_from_mem),         
/* input  logic    [72:0] */ .classifier_map_rewrite_15_from_mem           (classifier_map_rewrite_15_from_mem),         
/* input  logic    [72:0] */ .classifier_map_rewrite_1_from_mem            (classifier_map_rewrite_1_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_2_from_mem            (classifier_map_rewrite_2_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_3_from_mem            (classifier_map_rewrite_3_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_4_from_mem            (classifier_map_rewrite_4_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_5_from_mem            (classifier_map_rewrite_5_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_6_from_mem            (classifier_map_rewrite_6_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_7_from_mem            (classifier_map_rewrite_7_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_8_from_mem            (classifier_map_rewrite_8_from_mem),          
/* input  logic    [72:0] */ .classifier_map_rewrite_9_from_mem            (classifier_map_rewrite_9_from_mem),          
/* input  logic    [72:0] */ .classifier_map_type_from_mem                 (classifier_map_type_from_mem),               
/* input  logic    [72:0] */ .classifier_map_vpri_from_mem                 (classifier_map_vpri_from_mem),               
/* input  logic    [72:0] */ .classifier_map_vpri_tc_from_mem              (classifier_map_vpri_tc_from_mem),            
/* input  logic    [68:0] */ .classifier_wcm_action_cfg_0_from_mem         (classifier_wcm_action_cfg_0_from_mem),       
/* input  logic    [68:0] */ .classifier_wcm_action_cfg_1_from_mem         (classifier_wcm_action_cfg_1_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_0_from_mem         (classifier_wcm_action_ram_0_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_10_from_mem        (classifier_wcm_action_ram_10_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_11_from_mem        (classifier_wcm_action_ram_11_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_12_from_mem        (classifier_wcm_action_ram_12_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_13_from_mem        (classifier_wcm_action_ram_13_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_14_from_mem        (classifier_wcm_action_ram_14_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_15_from_mem        (classifier_wcm_action_ram_15_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_16_from_mem        (classifier_wcm_action_ram_16_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_17_from_mem        (classifier_wcm_action_ram_17_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_18_from_mem        (classifier_wcm_action_ram_18_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_19_from_mem        (classifier_wcm_action_ram_19_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_1_from_mem         (classifier_wcm_action_ram_1_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_20_from_mem        (classifier_wcm_action_ram_20_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_21_from_mem        (classifier_wcm_action_ram_21_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_22_from_mem        (classifier_wcm_action_ram_22_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_23_from_mem        (classifier_wcm_action_ram_23_from_mem),      
/* input  logic    [72:0] */ .classifier_wcm_action_ram_2_from_mem         (classifier_wcm_action_ram_2_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_3_from_mem         (classifier_wcm_action_ram_3_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_4_from_mem         (classifier_wcm_action_ram_4_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_5_from_mem         (classifier_wcm_action_ram_5_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_6_from_mem         (classifier_wcm_action_ram_6_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_7_from_mem         (classifier_wcm_action_ram_7_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_8_from_mem         (classifier_wcm_action_ram_8_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_action_ram_9_from_mem         (classifier_wcm_action_ram_9_from_mem),       
/* input  logic    [72:0] */ .classifier_wcm_data_path_buffer0_from_mem    (classifier_wcm_data_path_buffer0_from_mem),  
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_0_from_mem  (classifier_wcm_data_path_buffer1_0_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_10_from_mem (classifier_wcm_data_path_buffer1_10_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_11_from_mem (classifier_wcm_data_path_buffer1_11_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_12_from_mem (classifier_wcm_data_path_buffer1_12_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_13_from_mem (classifier_wcm_data_path_buffer1_13_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_14_from_mem (classifier_wcm_data_path_buffer1_14_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_15_from_mem (classifier_wcm_data_path_buffer1_15_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_16_from_mem (classifier_wcm_data_path_buffer1_16_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_17_from_mem (classifier_wcm_data_path_buffer1_17_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_18_from_mem (classifier_wcm_data_path_buffer1_18_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_19_from_mem (classifier_wcm_data_path_buffer1_19_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_1_from_mem  (classifier_wcm_data_path_buffer1_1_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_2_from_mem  (classifier_wcm_data_path_buffer1_2_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_3_from_mem  (classifier_wcm_data_path_buffer1_3_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_4_from_mem  (classifier_wcm_data_path_buffer1_4_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_5_from_mem  (classifier_wcm_data_path_buffer1_5_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_6_from_mem  (classifier_wcm_data_path_buffer1_6_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_7_from_mem  (classifier_wcm_data_path_buffer1_7_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_8_from_mem  (classifier_wcm_data_path_buffer1_8_from_mem), 
/* input  logic   [345:0] */ .classifier_wcm_data_path_buffer1_9_from_mem  (classifier_wcm_data_path_buffer1_9_from_mem), 
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_0_from_mem       (classifier_wcm_tcam_cfg_ram_0_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_10_from_mem      (classifier_wcm_tcam_cfg_ram_10_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_11_from_mem      (classifier_wcm_tcam_cfg_ram_11_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_12_from_mem      (classifier_wcm_tcam_cfg_ram_12_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_13_from_mem      (classifier_wcm_tcam_cfg_ram_13_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_14_from_mem      (classifier_wcm_tcam_cfg_ram_14_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_15_from_mem      (classifier_wcm_tcam_cfg_ram_15_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_16_from_mem      (classifier_wcm_tcam_cfg_ram_16_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_17_from_mem      (classifier_wcm_tcam_cfg_ram_17_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_18_from_mem      (classifier_wcm_tcam_cfg_ram_18_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_19_from_mem      (classifier_wcm_tcam_cfg_ram_19_from_mem),    
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_1_from_mem       (classifier_wcm_tcam_cfg_ram_1_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_2_from_mem       (classifier_wcm_tcam_cfg_ram_2_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_3_from_mem       (classifier_wcm_tcam_cfg_ram_3_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_4_from_mem       (classifier_wcm_tcam_cfg_ram_4_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_5_from_mem       (classifier_wcm_tcam_cfg_ram_5_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_6_from_mem       (classifier_wcm_tcam_cfg_ram_6_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_7_from_mem       (classifier_wcm_tcam_cfg_ram_7_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_8_from_mem       (classifier_wcm_tcam_cfg_ram_8_from_mem),     
/* input  logic    [70:0] */ .classifier_wcm_tcam_cfg_ram_9_from_mem       (classifier_wcm_tcam_cfg_ram_9_from_mem),     
/* input  logic  [1069:0] */ .classifier_wcm_tcam_from_tcam                (),                                           
/* input  logic           */ .clk                                          (cclk),                                       
/* input  logic           */ .em_a_delay_fifo_0_mem_ls_enter               (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_0_rd_adr                     (),                                           
/* input  logic           */ .em_a_delay_fifo_0_rd_en                      (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_0_wr_adr                     (),                                           
/* input  logic   [255:0] */ .em_a_delay_fifo_0_wr_data                    (),                                           
/* input  logic           */ .em_a_delay_fifo_0_wr_en                      (),                                           
/* input  logic           */ .em_a_delay_fifo_1_mem_ls_enter               (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_1_rd_adr                     (),                                           
/* input  logic           */ .em_a_delay_fifo_1_rd_en                      (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_1_wr_adr                     (),                                           
/* input  logic   [255:0] */ .em_a_delay_fifo_1_wr_data                    (),                                           
/* input  logic           */ .em_a_delay_fifo_1_wr_en                      (),                                           
/* input  logic           */ .em_a_delay_fifo_2_mem_ls_enter               (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_2_rd_adr                     (),                                           
/* input  logic           */ .em_a_delay_fifo_3_mem_ls_enter               (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_3_rd_adr                     (),                                           
/* input  logic           */ .em_a_delay_fifo_3_rd_en                      (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_3_wr_adr                     (),                                           
/* input  logic   [255:0] */ .em_a_delay_fifo_3_wr_data                    (),                                           
/* input  logic           */ .em_a_delay_fifo_3_wr_en                      (),                                           
/* input  logic           */ .em_a_hash_cfg_mem_ls_enter                   (),                                           
/* input  logic     [5:0] */ .em_a_hash_cfg_rd_adr                         (),                                           
/* input  logic           */ .em_a_hash_cfg_rd_en                          (),                                           
/* input  logic     [5:0] */ .em_a_hash_cfg_wr_adr                         (),                                           
/* input  logic    [52:0] */ .em_a_hash_cfg_wr_data                        (),                                           
/* input  logic           */ .em_a_hash_cfg_wr_en                          (),                                           
/* input  logic    [15:0] */ .em_a_hash_lookup_adr                         (),                                           
/* input  logic           */ .em_a_hash_lookup_mem_ls_enter                (),                                           
/* input  logic           */ .em_a_hash_lookup_rd_en                       (),                                           
/* input  logic    [71:0] */ .em_a_hash_lookup_wr_data                     (),                                           
/* input  logic           */ .em_a_hash_lookup_wr_en                       (),                                           
/* input  logic           */ .em_a_hash_miss_mem_ls_enter                  (),                                           
/* input  logic     [5:0] */ .em_a_hash_miss_rd_adr                        (),                                           
/* input  logic           */ .em_a_hash_miss_rd_en                         (),                                           
/* input  logic     [5:0] */ .em_a_hash_miss_wr_adr                        (),                                           
/* input  logic   [127:0] */ .em_a_hash_miss_wr_data                       (),                                           
/* input  logic           */ .em_a_hash_miss_wr_en                         (),                                           
/* input  logic           */ .em_a_key_mask_0_mem_ls_enter                 (),                                           
/* input  logic     [5:0] */ .em_a_key_mask_0_rd_adr                       (),                                           
/* input  logic           */ .em_a_key_mask_0_rd_en                        (),                                           
/* input  logic     [5:0] */ .em_a_key_mask_0_wr_adr                       (),                                           
/* input  logic    [63:0] */ .em_a_key_mask_0_wr_data                      (),                                           
/* input  logic           */ .em_a_key_mask_0_wr_en                        (),                                           
/* input  logic           */ .em_a_key_mask_1_mem_ls_enter                 (),                                           
/* input  logic     [5:0] */ .em_a_key_mask_1_rd_adr                       (),                                           
/* input  logic           */ .em_a_key_mask_1_rd_en                        (),                                           
/* input  logic     [5:0] */ .em_a_key_mask_1_wr_adr                       (),                                           
/* input  logic    [63:0] */ .em_a_key_mask_1_wr_data                      (),                                           
/* input  logic           */ .em_a_key_mask_1_wr_en                        (),                                           
/* input  logic           */ .em_a_key_mask_2_mem_ls_enter                 (),                                           
/* input  logic     [5:0] */ .em_a_key_mask_2_rd_adr                       (),                                           
/* input  logic           */ .em_a_key_mask_2_rd_en                        (),                                           
/* input  logic     [5:0] */ .em_a_key_mask_2_wr_adr                       (),                                           
/* input  logic    [63:0] */ .em_a_key_mask_2_wr_data                      (),                                           
/* input  logic           */ .em_a_key_mask_2_wr_en                        (),                                           
/* input  logic           */ .em_b_hash_cfg_mem_ls_enter                   (),                                           
/* input  logic     [5:0] */ .em_b_hash_cfg_rd_adr                         (),                                           
/* input  logic           */ .em_b_hash_cfg_rd_en                          (),                                           
/* input  logic     [5:0] */ .em_b_hash_cfg_wr_adr                         (),                                           
/* input  logic    [52:0] */ .em_b_hash_cfg_wr_data                        (),                                           
/* input  logic           */ .em_b_hash_cfg_wr_en                          (),                                           
/* input  logic    [12:0] */ .em_b_hash_lookup_adr                         (),                                           
/* input  logic           */ .em_b_hash_lookup_mem_ls_enter                (),                                           
/* input  logic           */ .em_b_hash_lookup_rd_en                       (),                                           
/* input  logic    [71:0] */ .em_b_hash_lookup_wr_data                     (),                                           
/* input  logic           */ .em_b_hash_lookup_wr_en                       (),                                           
/* input  logic           */ .em_b_hash_miss_mem_ls_enter                  (),                                           
/* input  logic     [5:0] */ .em_b_hash_miss_rd_adr                        (),                                           
/* input  logic           */ .em_b_hash_miss_rd_en                         (),                                           
/* input  logic     [5:0] */ .em_b_hash_miss_wr_adr                        (),                                           
/* input  logic   [127:0] */ .em_b_hash_miss_wr_data                       (),                                           
/* input  logic           */ .em_b_hash_miss_wr_en                         (),                                           
/* input  logic           */ .em_b_key_mask_mem_ls_enter                   (),                                           
/* input  logic     [5:0] */ .em_b_key_mask_rd_adr                         (),                                           
/* input  logic           */ .em_b_key_mask_rd_en                          (),                                           
/* input  logic     [5:0] */ .em_b_key_mask_wr_adr                         (),                                           
/* input  logic    [63:0] */ .em_b_key_mask_wr_data                        (),                                           
/* input  logic           */ .em_b_key_mask_wr_en                          (),                                           
/* input  logic     [8:0] */ .lpm_key_cam_adr                              (),                                           
/* input  logic           */ .lpm_key_cam_chk_en                           (),                                           
/* input  logic           */ .lpm_key_cam_chk_for_err_trig                 (),                                           
/* input  logic    [64:0] */ .lpm_key_cam_chk_key                          (),                                           
/* input  logic    [64:0] */ .lpm_key_cam_chk_mask                         (),                                           
/* input  logic   [255:0] */ .lpm_key_cam_raw_hit_in                       (),                                           
/* input  logic           */ .lpm_key_cam_rd_en                            (),                                           
/* input  logic     [3:0] */ .lpm_key_cam_slice_en                         (),                                           
/* input  logic    [64:0] */ .lpm_key_cam_wr_data                          (),                                           
/* input  logic           */ .lpm_key_cam_wr_en                            (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_0_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_0_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_0_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_0_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_0_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_10_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_10_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_11_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_11_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_11_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_11_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_12_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_12_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_12_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_12_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_12_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_13_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_13_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_13_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_13_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_13_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_14_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_14_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_14_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_14_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_14_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_15_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_15_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_15_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_15_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_15_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_16_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_16_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_16_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_16_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_16_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_17_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_17_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_17_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_17_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_17_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_18_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_18_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_18_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_18_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_18_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_19_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_19_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_19_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_19_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_19_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_1_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_1_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_1_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_1_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_1_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_20_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_20_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_20_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_20_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_20_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_21_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_21_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_21_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_21_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_21_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_22_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_22_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_22_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_22_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_22_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_23_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_23_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_23_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_23_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_23_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_24_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_24_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_24_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_24_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_24_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_25_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_25_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_25_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_25_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_25_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_26_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_26_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_26_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_26_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_26_wr_en                      (),                                           
/* input  logic           */ .lpm_tree_state_27_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_28_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_28_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_28_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_28_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_28_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_29_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_29_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_29_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_29_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_29_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_2_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_2_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_2_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_2_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_2_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_30_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_30_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_30_rd_en                      (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_1_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_1_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_1_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_1_wr_data              (),                                           
/* input  logic           */ .lpm_tree_state_31_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_31_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_31_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_32_adr                        (),                                           
/* input  logic           */ .wcm_data_path_buffer1_1_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_2_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_2_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_2_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_2_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_2_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_2_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_3_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_3_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_3_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_3_wr_adr               (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_33_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_33_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_33_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_33_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_33_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_34_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_34_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_34_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_34_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_34_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_35_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_35_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_35_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_35_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_35_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_36_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_36_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_36_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_36_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_36_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_37_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_37_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_37_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_37_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_37_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_38_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_38_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_38_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_38_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_38_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_39_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_39_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_39_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_39_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_39_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_3_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_3_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_3_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_3_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_3_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_40_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_40_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_40_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_40_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_40_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_41_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_41_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_41_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_41_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_41_wr_en                      (),                                           
/* input  logic           */ .lpm_tree_state_42_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_43_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_43_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_43_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_43_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_43_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_44_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_44_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_44_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_44_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_44_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_45_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_45_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_45_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_45_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_45_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_46_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_46_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_46_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_46_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_46_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_47_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_47_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_47_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_47_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_47_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_48_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_48_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_48_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_48_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_48_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_49_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_49_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_49_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_49_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_49_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_4_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_4_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_4_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_4_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_4_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_50_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_50_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_50_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_50_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_50_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_51_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_51_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_51_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_51_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_51_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_52_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_52_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_52_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_52_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_52_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_53_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_53_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_53_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_53_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_53_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_54_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_54_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_54_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_54_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_54_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_55_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_55_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_55_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_55_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_55_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_56_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_56_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_56_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_56_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_56_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_57_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_57_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_57_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_57_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_57_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_58_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_58_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_58_rd_en                      (),                                           
/* input  logic           */ .lpm_tree_state_59_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_59_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_59_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_5_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_5_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_5_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_5_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_5_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_60_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_60_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_60_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_60_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_60_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_61_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_61_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_61_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_61_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_61_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_62_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_62_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_62_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_62_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_62_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_63_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_63_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_63_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_63_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_63_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_64_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_64_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_64_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_64_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_64_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_65_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_65_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_65_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_65_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_65_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_66_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_66_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_66_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_66_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_66_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_67_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_67_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_67_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_67_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_67_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_68_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_68_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_68_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_68_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_68_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_69_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_69_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_69_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_69_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_69_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_6_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_6_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_6_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_6_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_6_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_70_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_70_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_70_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_70_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_70_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_71_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_71_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_71_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_71_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_71_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_72_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_72_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_72_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_72_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_72_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_73_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_73_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_73_rd_en                      (),                                           
/* input  logic           */ .lpm_tree_state_74_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_74_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_74_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_74_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_75_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_75_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_75_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_75_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_75_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_76_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_76_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_76_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_76_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_76_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_77_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_77_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_77_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_77_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_77_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_78_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_78_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_78_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_78_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_78_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_79_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_79_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_79_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_79_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_79_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_7_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_7_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_7_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_7_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_7_wr_en                       (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_80_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_80_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_80_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_80_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_80_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_81_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_81_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_81_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_81_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_81_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_82_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_82_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_82_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_82_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_82_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_83_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_83_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_83_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_83_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_83_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_84_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_84_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_84_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_84_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_84_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_85_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_85_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_85_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_85_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_85_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_86_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_86_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_86_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_86_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_86_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_87_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_87_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_87_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_87_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_87_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_88_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_88_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_88_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_88_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_88_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_89_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_89_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_89_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_89_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_89_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_8_adr                         (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_90_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_90_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_90_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_90_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_90_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_91_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_91_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_91_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_91_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_91_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_92_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_92_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_92_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_92_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_92_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_93_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_93_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_93_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_93_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_93_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_94_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_94_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_94_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_94_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_94_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_95_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_95_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_95_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_95_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_95_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_9_adr                         (),                                           
/* input  logic           */ .lpm_tree_state_9_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_9_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_9_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_9_wr_en                       (),                                           
/* input  logic    [11:0] */ .map_domain_action0_adr                       (),                                           
/* input  logic           */ .map_domain_action0_mem_ls_enter              (),                                           
/* input  logic           */ .map_domain_action0_rd_en                     (),                                           
/* input  logic    [63:0] */ .map_domain_action0_wr_data                   (),                                           
/* input  logic           */ .map_domain_action0_wr_en                     (),                                           
/* input  logic    [11:0] */ .map_domain_action1_adr                       (),                                           
/* input  logic           */ .map_domain_action1_mem_ls_enter              (),                                           
/* input  logic           */ .map_domain_action1_rd_en                     (),                                           
/* input  logic    [63:0] */ .map_domain_action1_wr_data                   (),                                           
/* input  logic           */ .map_domain_action1_wr_en                     (),                                           
/* input  logic           */ .map_domain_pol_cfg_mem_ls_enter              (),                                           
/* input  logic     [0:0] */ .map_domain_pol_cfg_rd_adr                    (),                                           
/* input  logic           */ .map_domain_pol_cfg_rd_en                     (),                                           
/* input  logic     [0:0] */ .map_domain_pol_cfg_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_domain_pol_cfg_wr_data                   (),                                           
/* input  logic           */ .map_domain_pol_cfg_wr_en                     (),                                           
/* input  logic     [8:0] */ .map_domain_profile_adr                       (),                                           
/* input  logic           */ .map_domain_profile_mem_ls_enter              (),                                           
/* input  logic           */ .map_domain_profile_rd_en                     (),                                           
/* input  logic    [63:0] */ .map_domain_profile_wr_data                   (),                                           
/* input  logic           */ .map_domain_profile_wr_en                     (),                                           
/* input  logic    [12:0] */ .map_domain_tcam_adr                          (),                                           
/* input  logic           */ .map_domain_tcam_chk_en                       (),                                           
/* input  logic           */ .map_domain_tcam_chk_for_err_trig             (),                                           
/* input  logic    [79:0] */ .map_domain_tcam_chk_key                      (),                                           
/* input  logic    [79:0] */ .map_domain_tcam_chk_mask                     (),                                           
/* input  logic  [4095:0] */ .map_domain_tcam_raw_hit_in                   (),                                           
/* input  logic           */ .map_domain_tcam_rd_en                        (),                                           
/* input  logic    [63:0] */ .map_domain_tcam_slice_en                     (),                                           
/* input  logic    [79:0] */ .map_domain_tcam_wr_data                      (),                                           
/* input  logic           */ .map_domain_tcam_wr_en                        (),                                           
/* input  logic    [10:0] */ .map_dscp_tc_adr                              (),                                           
/* input  logic           */ .map_dscp_tc_mem_ls_enter                     (),                                           
/* input  logic           */ .map_dscp_tc_rd_en                            (),                                           
/* input  logic    [63:0] */ .map_dscp_tc_wr_data                          (),                                           
/* input  logic           */ .map_dscp_tc_wr_en                            (),                                           
/* input  logic           */ .map_exp_tc_mem_ls_enter                      (),                                           
/* input  logic     [4:0] */ .map_exp_tc_rd_adr                            (),                                           
/* input  logic           */ .map_exp_tc_rd_en                             (),                                           
/* input  logic     [4:0] */ .map_exp_tc_wr_adr                            (),                                           
/* input  logic    [63:0] */ .map_exp_tc_wr_data                           (),                                           
/* input  logic           */ .map_exp_tc_wr_en                             (),                                           
/* input  logic           */ .map_extract_0_mem_ls_enter                   (),                                           
/* input  logic     [3:0] */ .map_extract_0_rd_adr                         (),                                           
/* input  logic           */ .map_extract_0_rd_en                          (),                                           
/* input  logic     [3:0] */ .map_extract_1_rd_adr                         (),                                           
/* input  logic           */ .map_extract_1_rd_en                          (),                                           
/* input  logic     [3:0] */ .map_extract_1_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_extract_1_wr_data                        (),                                           
/* input  logic           */ .map_extract_1_wr_en                          (),                                           
/* input  logic           */ .map_extract_2_mem_ls_enter                   (),                                           
/* input  logic     [3:0] */ .map_extract_2_rd_adr                         (),                                           
/* input  logic           */ .map_extract_2_rd_en                          (),                                           
/* input  logic     [3:0] */ .map_extract_2_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_extract_2_wr_data                        (),                                           
/* input  logic           */ .map_extract_2_wr_en                          (),                                           
/* input  logic           */ .map_ip_cfg_mem_ls_enter                      (),                                           
/* input  logic     [3:0] */ .map_ip_cfg_rd_adr                            (),                                           
/* input  logic           */ .map_ip_cfg_rd_en                             (),                                           
/* input  logic     [3:0] */ .map_ip_cfg_wr_adr                            (),                                           
/* input  logic    [63:0] */ .map_ip_cfg_wr_data                           (),                                           
/* input  logic           */ .map_ip_cfg_wr_en                             (),                                           
/* input  logic           */ .map_ip_hi_mem_ls_enter                       (),                                           
/* input  logic     [3:0] */ .map_ip_hi_rd_adr                             (),                                           
/* input  logic           */ .map_ip_hi_rd_en                              (),                                           
/* input  logic     [3:0] */ .map_ip_hi_wr_adr                             (),                                           
/* input  logic    [63:0] */ .map_ip_hi_wr_data                            (),                                           
/* input  logic           */ .map_ip_hi_wr_en                              (),                                           
/* input  logic           */ .map_ip_lo_mem_ls_enter                       (),                                           
/* input  logic     [3:0] */ .map_ip_lo_rd_adr                             (),                                           
/* input  logic           */ .map_ip_lo_rd_en                              (),                                           
/* input  logic     [3:0] */ .map_ip_lo_wr_adr                             (),                                           
/* input  logic    [63:0] */ .map_ip_lo_wr_data                            (),                                           
/* input  logic           */ .map_ip_lo_wr_en                              (),                                           
/* input  logic     [5:0] */ .map_l4_dst_adr                               (),                                           
/* input  logic           */ .map_l4_dst_mem_ls_enter                      (),                                           
/* input  logic           */ .map_l4_dst_rd_en                             (),                                           
/* input  logic    [63:0] */ .map_l4_dst_wr_data                           (),                                           
/* input  logic           */ .map_l4_dst_wr_en                             (),                                           
/* input  logic     [5:0] */ .map_l4_src_adr                               (),                                           
/* input  logic           */ .map_l4_src_mem_ls_enter                      (),                                           
/* input  logic           */ .map_l4_src_rd_en                             (),                                           
/* input  logic    [63:0] */ .map_l4_src_wr_data                           (),                                           
/* input  logic           */ .map_l4_src_wr_en                             (),                                           
/* input  logic           */ .map_len_limit_mem_ls_enter                   (),                                           
/* input  logic     [5:0] */ .map_len_limit_rd_adr                         (),                                           
/* input  logic           */ .map_len_limit_rd_en                          (),                                           
/* input  logic     [5:0] */ .map_len_limit_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_len_limit_wr_data                        (),                                           
/* input  logic           */ .map_len_limit_wr_en                          (),                                           
/* input  logic     [6:0] */ .map_mac_adr                                  (),                                           
/* input  logic           */ .map_mac_mem_ls_enter                         (),                                           
/* input  logic           */ .map_mac_rd_en                                (),                                           
/* input  logic   [127:0] */ .map_mac_wr_data                              (),                                           
/* input  logic           */ .map_mac_wr_en                                (),                                           
/* input  logic           */ .map_port_cfg_mem_ls_enter                    (),                                           
/* input  logic     [5:0] */ .map_port_cfg_rd_adr                          (),                                           
/* input  logic           */ .map_port_cfg_rd_en                           (),                                           
/* input  logic     [5:0] */ .map_port_cfg_wr_adr                          (),                                           
/* input  logic    [63:0] */ .map_port_cfg_wr_data                         (),                                           
/* input  logic           */ .map_port_cfg_wr_en                           (),                                           
/* input  logic           */ .map_port_default_0_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_0_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_0_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_0_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_0_wr_data                   (),                                           
/* input  logic           */ .map_port_default_0_wr_en                     (),                                           
/* input  logic           */ .map_port_default_10_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_10_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_10_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_10_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_10_wr_data                  (),                                           
/* input  logic           */ .map_port_default_10_wr_en                    (),                                           
/* input  logic           */ .map_port_default_11_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_11_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_11_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_11_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_11_wr_data                  (),                                           
/* input  logic           */ .map_port_default_11_wr_en                    (),                                           
/* input  logic           */ .map_port_default_12_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_12_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_12_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_12_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_12_wr_data                  (),                                           
/* input  logic           */ .map_port_default_12_wr_en                    (),                                           
/* input  logic           */ .map_port_default_13_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_13_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_13_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_13_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_13_wr_data                  (),                                           
/* input  logic     [2:0] */ .map_port_default_14_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_14_wr_data                  (),                                           
/* input  logic           */ .map_port_default_14_wr_en                    (),                                           
/* input  logic           */ .map_port_default_15_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_15_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_15_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_15_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_15_wr_data                  (),                                           
/* input  logic           */ .map_port_default_15_wr_en                    (),                                           
/* input  logic           */ .map_port_default_16_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_16_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_16_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_16_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_16_wr_data                  (),                                           
/* input  logic           */ .map_port_default_16_wr_en                    (),                                           
/* input  logic           */ .map_port_default_17_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_17_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_17_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_17_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_17_wr_data                  (),                                           
/* input  logic           */ .map_port_default_17_wr_en                    (),                                           
/* input  logic           */ .map_port_default_18_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_18_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_18_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_18_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_18_wr_data                  (),                                           
/* input  logic           */ .map_port_default_18_wr_en                    (),                                           
/* input  logic           */ .map_port_default_19_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_19_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_19_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_19_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_19_wr_data                  (),                                           
/* input  logic           */ .map_port_default_19_wr_en                    (),                                           
/* input  logic           */ .map_port_default_1_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_1_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_1_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_1_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_1_wr_data                   (),                                           
/* input  logic           */ .map_port_default_1_wr_en                     (),                                           
/* input  logic           */ .map_port_default_20_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_20_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_20_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_20_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_20_wr_data                  (),                                           
/* input  logic           */ .map_port_default_20_wr_en                    (),                                           
/* input  logic           */ .map_port_default_21_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_21_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_21_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_21_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_21_wr_data                  (),                                           
/* input  logic           */ .map_port_default_21_wr_en                    (),                                           
/* input  logic           */ .map_port_default_22_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_22_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_22_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_22_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_22_wr_data                  (),                                           
/* input  logic           */ .map_port_default_22_wr_en                    (),                                           
/* input  logic           */ .map_port_default_23_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_23_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_23_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_23_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_23_wr_data                  (),                                           
/* input  logic           */ .map_port_default_23_wr_en                    (),                                           
/* input  logic           */ .map_port_default_24_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_24_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_24_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_24_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_24_wr_data                  (),                                           
/* input  logic           */ .map_port_default_24_wr_en                    (),                                           
/* input  logic           */ .map_port_default_25_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_25_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_25_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_25_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_25_wr_data                  (),                                           
/* input  logic           */ .map_port_default_25_wr_en                    (),                                           
/* input  logic           */ .map_port_default_26_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_26_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_26_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_26_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_26_wr_data                  (),                                           
/* input  logic     [2:0] */ .map_port_default_27_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_27_wr_data                  (),                                           
/* input  logic           */ .map_port_default_27_wr_en                    (),                                           
/* input  logic           */ .map_port_default_28_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_28_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_28_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_28_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_28_wr_data                  (),                                           
/* input  logic           */ .map_port_default_28_wr_en                    (),                                           
/* input  logic           */ .map_port_default_29_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_29_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_29_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_29_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_29_wr_data                  (),                                           
/* input  logic           */ .map_port_default_29_wr_en                    (),                                           
/* input  logic           */ .map_port_default_2_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_2_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_2_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_2_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_2_wr_data                   (),                                           
/* input  logic           */ .map_port_default_2_wr_en                     (),                                           
/* input  logic           */ .map_port_default_30_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_30_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_30_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_30_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_30_wr_data                  (),                                           
/* input  logic           */ .map_port_default_30_wr_en                    (),                                           
/* input  logic           */ .map_port_default_31_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_31_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_31_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_31_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_31_wr_data                  (),                                           
/* input  logic           */ .map_port_default_31_wr_en                    (),                                           
/* input  logic           */ .map_port_default_32_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_32_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_32_rd_en                    (),                                           
/* input  logic     [2:0] */ .map_port_default_32_wr_adr                   (),                                           
/* input  logic    [63:0] */ .map_port_default_32_wr_data                  (),                                           
/* input  logic           */ .map_port_default_32_wr_en                    (),                                           
/* input  logic           */ .map_port_default_3_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_3_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_3_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_3_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_3_wr_data                   (),                                           
/* input  logic           */ .map_port_default_3_wr_en                     (),                                           
/* input  logic           */ .map_port_default_4_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_4_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_4_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_4_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_4_wr_data                   (),                                           
/* input  logic           */ .map_port_default_4_wr_en                     (),                                           
/* input  logic           */ .map_port_default_5_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_5_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_5_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_5_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_5_wr_data                   (),                                           
/* input  logic           */ .map_port_default_5_wr_en                     (),                                           
/* input  logic           */ .map_port_default_6_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_6_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_6_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_6_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_6_wr_data                   (),                                           
/* input  logic           */ .map_port_default_6_wr_en                     (),                                           
/* input  logic           */ .map_port_default_7_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_7_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_7_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_7_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_7_wr_data                   (),                                           
/* input  logic           */ .map_port_default_7_wr_en                     (),                                           
/* input  logic           */ .map_port_default_8_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_8_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_8_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_8_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_8_wr_data                   (),                                           
/* input  logic           */ .map_port_default_8_wr_en                     (),                                           
/* input  logic           */ .map_port_default_9_mem_ls_enter              (),                                           
/* input  logic     [2:0] */ .map_port_default_9_rd_adr                    (),                                           
/* input  logic           */ .map_port_default_9_rd_en                     (),                                           
/* input  logic     [2:0] */ .map_port_default_9_wr_adr                    (),                                           
/* input  logic    [63:0] */ .map_port_default_9_wr_data                   (),                                           
/* input  logic           */ .map_port_default_9_wr_en                     (),                                           
/* input  logic    [79:0] */ .map_profile_key0_wr_data                     (),                                           
/* input  logic           */ .map_profile_key0_wr_en                       (),                                           
/* input  logic           */ .map_profile_key1_mem_ls_enter                (),                                           
/* input  logic     [6:0] */ .map_profile_key1_rd_adr                      (),                                           
/* input  logic           */ .map_profile_key1_rd_en                       (),                                           
/* input  logic     [6:0] */ .map_profile_key1_wr_adr                      (),                                           
/* input  logic    [79:0] */ .map_profile_key1_wr_data                     (),                                           
/* input  logic           */ .map_profile_key1_wr_en                       (),                                           
/* input  logic           */ .map_profile_key_invert0_mem_ls_enter         (),                                           
/* input  logic     [6:0] */ .map_profile_key_invert0_rd_adr               (),                                           
/* input  logic           */ .map_profile_key_invert0_rd_en                (),                                           
/* input  logic     [6:0] */ .map_profile_key_invert0_wr_adr               (),                                           
/* input  logic    [79:0] */ .map_profile_key_invert0_wr_data              (),                                           
/* input  logic           */ .map_profile_key_invert0_wr_en                (),                                           
/* input  logic           */ .map_profile_key_invert1_mem_ls_enter         (),                                           
/* input  logic     [6:0] */ .map_profile_key_invert1_rd_adr               (),                                           
/* input  logic           */ .map_profile_key_invert1_rd_en                (),                                           
/* input  logic     [6:0] */ .map_profile_key_invert1_wr_adr               (),                                           
/* input  logic    [79:0] */ .map_profile_key_invert1_wr_data              (),                                           
/* input  logic           */ .map_profile_key_invert1_wr_en                (),                                           
/* input  logic           */ .map_prot_mem_ls_enter                        (),                                           
/* input  logic     [2:0] */ .map_prot_rd_adr                              (),                                           
/* input  logic           */ .map_prot_rd_en                               (),                                           
/* input  logic     [2:0] */ .map_prot_wr_adr                              (),                                           
/* input  logic    [63:0] */ .map_prot_wr_data                             (),                                           
/* input  logic           */ .map_prot_wr_en                               (),                                           
/* input  logic           */ .map_rewrite_0_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_0_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_0_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_0_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_0_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_0_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_10_mem_ls_enter                  (),                                           
/* input  logic     [4:0] */ .map_rewrite_10_rd_adr                        (),                                           
/* input  logic           */ .map_rewrite_10_rd_en                         (),                                           
/* input  logic     [4:0] */ .map_rewrite_10_wr_adr                        (),                                           
/* input  logic    [63:0] */ .map_rewrite_10_wr_data                       (),                                           
/* input  logic           */ .map_rewrite_10_wr_en                         (),                                           
/* input  logic           */ .map_rewrite_11_mem_ls_enter                  (),                                           
/* input  logic     [4:0] */ .map_rewrite_11_rd_adr                        (),                                           
/* input  logic           */ .map_rewrite_11_rd_en                         (),                                           
/* input  logic     [4:0] */ .map_rewrite_11_wr_adr                        (),                                           
/* input  logic    [63:0] */ .map_rewrite_11_wr_data                       (),                                           
/* input  logic           */ .map_rewrite_11_wr_en                         (),                                           
/* input  logic           */ .map_rewrite_12_mem_ls_enter                  (),                                           
/* input  logic     [4:0] */ .map_rewrite_12_rd_adr                        (),                                           
/* input  logic           */ .map_rewrite_12_rd_en                         (),                                           
/* input  logic     [4:0] */ .map_rewrite_12_wr_adr                        (),                                           
/* input  logic    [63:0] */ .map_rewrite_12_wr_data                       (),                                           
/* input  logic           */ .map_rewrite_12_wr_en                         (),                                           
/* input  logic           */ .map_rewrite_13_mem_ls_enter                  (),                                           
/* input  logic     [4:0] */ .map_rewrite_13_rd_adr                        (),                                           
/* input  logic           */ .map_rewrite_13_rd_en                         (),                                           
/* input  logic     [4:0] */ .map_rewrite_13_wr_adr                        (),                                           
/* input  logic    [63:0] */ .map_rewrite_13_wr_data                       (),                                           
/* input  logic           */ .map_rewrite_13_wr_en                         (),                                           
/* input  logic           */ .map_rewrite_14_mem_ls_enter                  (),                                           
/* input  logic     [4:0] */ .map_rewrite_14_rd_adr                        (),                                           
/* input  logic           */ .map_rewrite_14_rd_en                         (),                                           
/* input  logic     [4:0] */ .map_rewrite_14_wr_adr                        (),                                           
/* input  logic    [63:0] */ .map_rewrite_14_wr_data                       (),                                           
/* input  logic           */ .map_rewrite_14_wr_en                         (),                                           
/* input  logic           */ .map_rewrite_15_mem_ls_enter                  (),                                           
/* input  logic     [4:0] */ .map_rewrite_15_rd_adr                        (),                                           
/* input  logic           */ .map_rewrite_15_rd_en                         (),                                           
/* input  logic     [4:0] */ .map_rewrite_15_wr_adr                        (),                                           
/* input  logic    [63:0] */ .map_rewrite_15_wr_data                       (),                                           
/* input  logic           */ .map_rewrite_15_wr_en                         (),                                           
/* input  logic           */ .map_rewrite_1_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_1_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_1_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_1_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_1_wr_data                        (),                                           
/* input  logic     [4:0] */ .map_rewrite_2_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_2_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_2_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_3_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_3_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_3_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_3_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_3_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_3_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_4_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_4_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_4_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_4_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_4_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_4_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_5_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_5_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_5_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_5_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_5_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_5_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_6_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_6_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_6_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_6_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_6_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_6_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_7_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_7_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_7_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_7_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_7_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_7_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_8_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_8_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_8_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_8_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_8_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_8_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_9_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_9_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_9_rd_en                          (),                                           
/* input  logic     [4:0] */ .map_rewrite_9_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_rewrite_9_wr_data                        (),                                           
/* input  logic           */ .map_rewrite_9_wr_en                          (),                                           
/* input  logic           */ .map_type_mem_ls_enter                        (),                                           
/* input  logic     [3:0] */ .map_type_rd_adr                              (),                                           
/* input  logic           */ .map_type_rd_en                               (),                                           
/* input  logic     [3:0] */ .map_type_wr_adr                              (),                                           
/* input  logic    [63:0] */ .map_type_wr_data                             (),                                           
/* input  logic           */ .map_type_wr_en                               (),                                           
/* input  logic           */ .map_vpri_mem_ls_enter                        (),                                           
/* input  logic     [4:0] */ .map_vpri_rd_adr                              (),                                           
/* input  logic           */ .map_vpri_rd_en                               (),                                           
/* input  logic           */ .map_vpri_tc_mem_ls_enter                     (),                                           
/* input  logic     [4:0] */ .map_vpri_tc_rd_adr                           (),                                           
/* input  logic           */ .map_vpri_tc_rd_en                            (),                                           
/* input  logic     [4:0] */ .map_vpri_tc_wr_adr                           (),                                           
/* input  logic    [63:0] */ .map_vpri_tc_wr_data                          (),                                           
/* input  logic           */ .map_vpri_tc_wr_en                            (),                                           
/* input  logic     [4:0] */ .map_vpri_wr_adr                              (),                                           
/* input  logic    [63:0] */ .map_vpri_wr_data                             (),                                           
/* input  logic           */ .map_vpri_wr_en                               (),                                           
/* input  logic           */ .reset_n                                      (reset_n),                                    
/* input  logic           */ .unified_regs_rd                              (),                                           
/* input  logic    [31:0] */ .unified_regs_wr_data                         (),                                           
/* input  logic    [11:0] */ .wcm_action_cfg_0_adr                         (),                                           
/* input  logic           */ .wcm_action_cfg_0_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_cfg_0_rd_en                       (),                                           
/* input  logic    [59:0] */ .wcm_action_cfg_0_wr_data                     (),                                           
/* input  logic           */ .wcm_action_cfg_0_wr_en                       (),                                           
/* input  logic    [11:0] */ .wcm_action_cfg_1_adr                         (),                                           
/* input  logic           */ .wcm_action_cfg_1_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_cfg_1_rd_en                       (),                                           
/* input  logic    [59:0] */ .wcm_action_cfg_1_wr_data                     (),                                           
/* input  logic           */ .wcm_action_cfg_1_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_0_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_0_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_0_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_0_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_0_wr_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_10_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_10_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_11_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_11_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_11_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_11_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_11_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_12_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_12_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_12_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_12_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_12_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_13_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_13_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_13_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_13_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_13_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_14_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_14_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_14_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_14_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_14_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_15_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_15_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_15_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_15_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_15_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_16_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_16_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_16_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_16_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_16_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_17_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_17_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_17_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_17_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_17_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_18_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_18_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_18_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_18_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_18_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_19_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_19_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_19_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_19_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_19_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_1_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_1_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_1_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_1_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_1_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_20_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_20_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_20_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_20_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_20_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_21_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_21_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_21_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_21_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_21_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_22_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_22_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_22_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_22_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_22_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_23_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_23_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_23_rd_en                      (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_23_wr_data                    (),                                           
/* input  logic           */ .wcm_action_ram_23_wr_en                      (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_2_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_2_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_2_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_2_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_2_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_3_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_3_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_3_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_3_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_3_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_4_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_4_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_4_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_4_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_4_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_5_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_5_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_5_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_5_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_5_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_6_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_6_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_6_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_6_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_6_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_7_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_7_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_7_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_7_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_7_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_8_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_8_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_8_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_8_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_8_wr_en                       (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_9_adr                         (),                                           
/* input  logic           */ .wcm_action_ram_9_mem_ls_enter                (),                                           
/* input  logic           */ .wcm_action_ram_9_rd_en                       (),                                           
/* input  logic    [63:0] */ .wcm_action_ram_9_wr_data                     (),                                           
/* input  logic           */ .wcm_action_ram_9_wr_en                       (),                                           
/* input  logic           */ .wcm_data_path_buffer0_mem_ls_enter           (),                                           
/* input  logic     [2:0] */ .wcm_data_path_buffer0_rd_adr                 (),                                           
/* input  logic           */ .wcm_data_path_buffer0_rd_en                  (),                                           
/* input  logic     [2:0] */ .wcm_data_path_buffer0_wr_adr                 (),                                           
/* input  logic    [63:0] */ .wcm_data_path_buffer0_wr_data                (),                                           
/* input  logic           */ .wcm_data_path_buffer0_wr_en                  (),                                           
/* input  logic           */ .wcm_data_path_buffer1_0_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_0_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_0_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_0_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_0_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_0_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_10_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_10_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_10_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_10_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_10_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_10_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_11_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_11_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_11_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_11_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_11_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_11_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_12_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_12_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_12_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_12_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_12_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_12_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_13_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_13_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_13_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_13_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_13_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_13_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_14_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_14_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_14_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_14_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_14_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_14_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_15_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_15_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_15_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_15_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_15_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_15_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_16_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_16_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_16_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_16_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_16_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_16_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_17_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_17_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_17_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_18_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_18_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_18_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_18_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_18_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_19_mem_ls_enter        (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_19_rd_adr              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_19_rd_en               (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_19_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_19_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_19_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_1_mem_ls_enter         (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_3_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_3_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_4_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_4_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_4_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_4_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_4_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_4_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_5_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_5_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_5_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_5_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_5_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_5_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_6_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_6_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_6_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_6_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_6_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_6_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_7_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_7_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_7_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_7_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_7_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_7_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_8_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_8_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_8_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_8_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_8_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_8_wr_en                (),                                           
/* input  logic           */ .wcm_data_path_buffer1_9_mem_ls_enter         (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_9_rd_adr               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_9_rd_en                (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_9_wr_adr               (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_9_wr_data              (),                                           
/* input  logic           */ .wcm_data_path_buffer1_9_wr_en                (),                                           
/* input  logic    [10:0] */ .wcm_tcam_0_adr                               (),                                           
/* input  logic           */ .wcm_tcam_0_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_0_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_0_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_0_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_0_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_0_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_0_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_0_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_0_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_10_adr                              (),                                           
/* input  logic           */ .wcm_tcam_10_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_10_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_10_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_10_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_10_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_10_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_10_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_10_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_10_wr_en                            (),                                           
/* input  logic    [39:0] */ .wcm_tcam_11_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_11_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_11_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_11_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_11_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_11_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_12_adr                              (),                                           
/* input  logic           */ .wcm_tcam_12_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_12_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_12_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_12_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_12_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_12_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_12_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_12_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_12_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_13_adr                              (),                                           
/* input  logic           */ .wcm_tcam_13_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_13_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_13_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_13_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_13_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_13_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_13_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_13_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_13_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_14_adr                              (),                                           
/* input  logic           */ .wcm_tcam_14_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_14_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_14_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_14_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_14_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_14_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_14_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_14_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_14_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_15_adr                              (),                                           
/* input  logic           */ .wcm_tcam_15_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_15_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_15_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_15_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_15_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_15_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_15_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_15_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_15_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_16_adr                              (),                                           
/* input  logic           */ .wcm_tcam_16_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_16_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_16_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_16_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_16_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_16_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_16_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_16_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_16_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_17_adr                              (),                                           
/* input  logic           */ .wcm_tcam_17_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_17_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_17_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_17_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_17_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_17_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_17_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_17_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_17_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_18_adr                              (),                                           
/* input  logic           */ .wcm_tcam_18_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_18_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_18_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_18_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_18_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_18_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_18_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_18_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_18_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_19_adr                              (),                                           
/* input  logic           */ .wcm_tcam_19_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_19_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_19_chk_key                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_19_wr_data                          (),                                           
/* input  logic           */ .wcm_tcam_19_wr_en                            (),                                           
/* input  logic    [10:0] */ .wcm_tcam_1_adr                               (),                                           
/* input  logic           */ .wcm_tcam_1_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_1_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_1_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_1_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_1_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_1_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_1_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_1_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_1_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_2_adr                               (),                                           
/* input  logic           */ .wcm_tcam_2_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_2_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_2_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_2_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_2_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_2_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_2_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_2_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_2_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_3_adr                               (),                                           
/* input  logic           */ .wcm_tcam_3_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_3_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_3_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_3_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_3_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_3_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_3_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_3_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_3_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_4_adr                               (),                                           
/* input  logic           */ .wcm_tcam_4_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_4_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_4_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_4_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_4_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_4_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_4_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_4_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_4_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_5_adr                               (),                                           
/* input  logic           */ .wcm_tcam_5_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_5_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_5_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_5_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_5_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_5_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_5_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_5_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_5_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_6_adr                               (),                                           
/* input  logic           */ .wcm_tcam_6_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_6_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_6_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_6_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_6_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_6_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_6_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_6_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_6_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_7_adr                               (),                                           
/* input  logic           */ .wcm_tcam_7_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_7_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_7_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_7_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_7_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_7_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_7_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_7_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_7_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_8_adr                               (),                                           
/* input  logic           */ .wcm_tcam_8_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_8_chk_for_err_trig                  (),                                           
/* input  logic    [39:0] */ .wcm_tcam_8_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_8_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_8_raw_hit_in                        (),                                           
/* input  logic           */ .wcm_tcam_8_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_8_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_8_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_8_wr_en                             (),                                           
/* input  logic    [10:0] */ .wcm_tcam_9_adr                               (),                                           
/* input  logic           */ .wcm_tcam_9_chk_en                            (),                                           
/* input  logic           */ .wcm_tcam_9_chk_for_err_trig                  (),                                           
/* input  logic           */ .wcm_tcam_9_rd_en                             (),                                           
/* input  logic    [15:0] */ .wcm_tcam_9_slice_en                          (),                                           
/* input  logic    [39:0] */ .wcm_tcam_9_wr_data                           (),                                           
/* input  logic           */ .wcm_tcam_9_wr_en                             (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_0_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_0_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_0_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_0_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_0_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_10_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_10_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_10_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_10_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_10_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_11_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_11_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_11_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_11_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_11_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_12_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_12_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_12_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_12_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_12_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_13_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_13_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_13_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_13_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_13_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_14_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_14_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_14_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_14_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_14_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_15_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_15_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_15_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_15_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_15_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_16_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_16_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_16_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_16_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_16_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_17_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_17_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_17_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_17_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_17_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_18_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_18_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_18_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_18_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_18_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_19_adr                      (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_19_mem_ls_enter             (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_19_rd_en                    (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_19_wr_data                  (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_19_wr_en                    (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_1_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_1_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_1_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_1_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_1_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_2_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_2_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_2_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_2_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_2_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_3_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_3_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_3_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_3_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_3_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_4_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_4_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_4_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_4_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_4_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_5_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_5_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_6_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_6_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_6_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_6_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_7_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_7_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_7_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_7_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_7_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_8_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_8_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_8_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_8_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_8_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_9_adr                       (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_9_mem_ls_enter              (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_9_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_9_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_9_wr_en                     (),                                           
/* input  logic    [63:0] */ .map_port_wr_data                             (),                                           
/* input  logic           */ .map_port_wr_en                               (),                                           
/* input  logic     [6:0] */ .map_profile_action_adr                       (),                                           
/* input  logic           */ .map_profile_action_mem_ls_enter              (),                                           
/* input  logic           */ .map_profile_action_rd_en                     (),                                           
/* input  logic    [63:0] */ .map_profile_action_wr_data                   (),                                           
/* input  logic           */ .map_profile_action_wr_en                     (),                                           
/* input  logic           */ .map_profile_key0_mem_ls_enter                (),                                           
/* input  logic     [6:0] */ .map_profile_key0_rd_adr                      (),                                           
/* input  logic           */ .map_profile_key0_rd_en                       (),                                           
/* input  logic     [6:0] */ .map_profile_key0_wr_adr                      (),                                           
/* input  logic           */ .CLASSIFIER_ECC_COR_ERR_reg_sel               (),                                           
/* input  logic           */ .CLASSIFIER_ECC_UNCOR_ERR_reg_sel             (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_0_CFG_reg_sel                (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_0_STATUS_reg_sel             (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_1_CFG_reg_sel                (),                                           
/* input  logic     [3:0] */ .map_extract_0_wr_adr                         (),                                           
/* input  logic    [63:0] */ .map_extract_0_wr_data                        (),                                           
/* input  logic           */ .map_extract_0_wr_en                          (),                                           
/* input  logic           */ .map_extract_1_mem_ls_enter                   (),                                           
/* input  logic           */ .map_port_default_13_wr_en                    (),                                           
/* input  logic           */ .map_port_default_14_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_14_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_14_rd_en                    (),                                           
/* input  logic   [306:0] */ .classifier_lpm_tree_state_22_from_mem        (classifier_lpm_tree_state_22_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_23_from_mem        (classifier_lpm_tree_state_23_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_24_from_mem        (classifier_lpm_tree_state_24_from_mem),      
/* input  logic   [306:0] */ .classifier_lpm_tree_state_25_from_mem        (classifier_lpm_tree_state_25_from_mem),      
/* input  logic           */ .lpm_tree_state_10_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_10_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_10_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_11_adr                        (),                                           
/* input  logic           */ .MAP_DOMAIN_POL_CFG_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_DOMAIN_POL_CFG_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_DOMAIN_PROFILE_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_DOMAIN_PROFILE_STATUS_reg_sel            (),                                           
/* input  logic     [9:0] */ .wcm_action_ram_10_adr                        (),                                           
/* input  logic           */ .wcm_action_ram_10_mem_ls_enter               (),                                           
/* input  logic           */ .wcm_action_ram_10_rd_en                      (),                                           
/* input  logic     [4:0] */ .wcm_data_path_buffer1_17_wr_adr              (),                                           
/* input  logic   [334:0] */ .wcm_data_path_buffer1_17_wr_data             (),                                           
/* input  logic           */ .wcm_data_path_buffer1_17_wr_en               (),                                           
/* input  logic           */ .wcm_data_path_buffer1_18_mem_ls_enter        (),                                           
/* input  logic    [10:0] */ .wcm_tcam_11_adr                              (),                                           
/* input  logic           */ .wcm_tcam_11_chk_en                           (),                                           
/* input  logic           */ .wcm_tcam_11_chk_for_err_trig                 (),                                           
/* input  logic    [39:0] */ .wcm_tcam_11_chk_key                          (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_5_rd_en                     (),                                           
/* input  logic    [61:0] */ .wcm_tcam_cfg_ram_5_wr_data                   (),                                           
/* input  logic           */ .wcm_tcam_cfg_ram_5_wr_en                     (),                                           
/* input  logic     [9:0] */ .wcm_tcam_cfg_ram_6_adr                       (),                                           
/* input  logic    [72:0] */ .classifier_map_port_default_30_from_mem      (classifier_map_port_default_30_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_31_from_mem      (classifier_map_port_default_31_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_32_from_mem      (classifier_map_port_default_32_from_mem),    
/* input  logic    [72:0] */ .classifier_map_port_default_3_from_mem       (classifier_map_port_default_3_from_mem),     
/* input  logic           */ .em_a_delay_fifo_2_rd_en                      (),                                           
/* input  logic     [5:0] */ .em_a_delay_fifo_2_wr_adr                     (),                                           
/* input  logic   [255:0] */ .em_a_delay_fifo_2_wr_data                    (),                                           
/* input  logic           */ .em_a_delay_fifo_2_wr_en                      (),                                           
/* input  logic           */ .LPM_TREE_STATE_5_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_60_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_60_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_61_CFG_reg_sel                (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_4_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_5_CFG_reg_sel               (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_5_STATUS_reg_sel            (),                                           
/* input  logic           */ .MAP_PORT_DEFAULT_6_CFG_reg_sel               (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_27_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_27_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_27_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_27_wr_data                    (),                                           
/* input  logic           */ .WCM_ACTION_RAM_18_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_19_CFG_reg_sel                (),                                           
/* input  logic           */ .WCM_ACTION_RAM_19_STATUS_reg_sel             (),                                           
/* input  logic           */ .WCM_ACTION_RAM_1_CFG_reg_sel                 (),                                           
/* input  logic           */ .WCM_TCAM_15_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_16_CFG_reg_sel                      (),                                           
/* input  logic           */ .WCM_TCAM_16_STATUS_reg_sel                   (),                                           
/* input  logic           */ .WCM_TCAM_17_CFG_reg_sel                      (),                                           
/* input  logic           */ .LPM_TREE_STATE_21_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_22_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_22_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_23_CFG_reg_sel                (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_42_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_42_mem_ls_enter               (),                                           
/* input  logic           */ .lpm_tree_state_42_rd_en                      (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_42_wr_data                    (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_58_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_58_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_59_adr                        (),                                           
/* input  logic           */ .lpm_tree_state_59_mem_ls_enter               (),                                           
/* input  logic           */ .map_port_mem_ls_enter                        (),                                           
/* input  logic     [5:0] */ .map_port_rd_adr                              (),                                           
/* input  logic           */ .map_port_rd_en                               (),                                           
/* input  logic     [5:0] */ .map_port_wr_adr                              (),                                           
/* input  logic           */ .map_rewrite_1_wr_en                          (),                                           
/* input  logic           */ .map_rewrite_2_mem_ls_enter                   (),                                           
/* input  logic     [4:0] */ .map_rewrite_2_rd_adr                         (),                                           
/* input  logic           */ .map_rewrite_2_rd_en                          (),                                           
/* input  logic           */ .lpm_tree_state_8_mem_ls_enter                (),                                           
/* input  logic           */ .lpm_tree_state_8_rd_en                       (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_8_wr_data                     (),                                           
/* input  logic           */ .lpm_tree_state_8_wr_en                       (),                                           
/* input  logic           */ .map_port_default_26_wr_en                    (),                                           
/* input  logic           */ .map_port_default_27_mem_ls_enter             (),                                           
/* input  logic     [2:0] */ .map_port_default_27_rd_adr                   (),                                           
/* input  logic           */ .map_port_default_27_rd_en                    (),                                           
/* input  logic   [295:0] */ .lpm_tree_state_73_wr_data                    (),                                           
/* input  logic           */ .lpm_tree_state_73_wr_en                      (),                                           
/* input  logic     [8:0] */ .lpm_tree_state_74_adr                        (),                                           
/* input  logic    [39:0] */ .wcm_tcam_19_chk_mask                         (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_19_raw_hit_in                       (),                                           
/* input  logic           */ .wcm_tcam_19_rd_en                            (),                                           
/* input  logic    [15:0] */ .wcm_tcam_19_slice_en                         (),                                           
/* input  logic    [39:0] */ .wcm_tcam_9_chk_key                           (),                                           
/* input  logic    [39:0] */ .wcm_tcam_9_chk_mask                          (),                                           
/* input  logic  [1023:0] */ .wcm_tcam_9_raw_hit_in                        (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_1_STATUS_reg_sel             (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_2_CFG_reg_sel                (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_2_STATUS_reg_sel             (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_3_CFG_reg_sel                (),                                           
/* input  logic           */ .EM_A_DELAY_FIFO_3_STATUS_reg_sel             (),                                           
/* input  logic           */ .EM_A_HASH_CFG_CFG_reg_sel                    (),                                           
/* input  logic           */ .EM_A_HASH_CFG_STATUS_reg_sel                 (),                                           
/* input  logic           */ .EM_A_HASH_LOOKUP_CFG_reg_sel                 (),                                           
/* input  logic           */ .EM_A_HASH_LOOKUP_STATUS_reg_sel              (),                                           
/* input  logic           */ .EM_A_HASH_MISS_CFG_reg_sel                   (),                                           
/* input  logic           */ .EM_A_HASH_MISS_STATUS_reg_sel                (),                                           
/* input  logic           */ .EM_A_KEY_MASK_0_CFG_reg_sel                  (),                                           
/* input  logic           */ .EM_A_KEY_MASK_0_STATUS_reg_sel               (),                                           
/* input  logic           */ .EM_A_KEY_MASK_1_CFG_reg_sel                  (),                                           
/* input  logic           */ .EM_A_KEY_MASK_1_STATUS_reg_sel               (),                                           
/* input  logic           */ .EM_A_KEY_MASK_2_CFG_reg_sel                  (),                                           
/* input  logic           */ .EM_A_KEY_MASK_2_STATUS_reg_sel               (),                                           
/* input  logic           */ .EM_B_HASH_CFG_CFG_reg_sel                    (),                                           
/* input  logic           */ .EM_B_HASH_CFG_STATUS_reg_sel                 (),                                           
/* input  logic           */ .EM_B_HASH_LOOKUP_CFG_reg_sel                 (),                                           
/* input  logic           */ .EM_B_HASH_LOOKUP_STATUS_reg_sel              (),                                           
/* input  logic           */ .EM_B_HASH_MISS_CFG_reg_sel                   (),                                           
/* input  logic           */ .EM_B_HASH_MISS_STATUS_reg_sel                (),                                           
/* input  logic           */ .EM_B_KEY_MASK_CFG_reg_sel                    (),                                           
/* input  logic           */ .EM_B_KEY_MASK_STATUS_reg_sel                 (),                                           
/* input  logic           */ .LPM_KEY_CAM_CFG_reg_sel                      (),                                           
/* input  logic           */ .LPM_KEY_CAM_STATUS_reg_sel                   (),                                           
/* input  logic           */ .LPM_TREE_STATE_0_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_0_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_10_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_10_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_11_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_11_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_12_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_12_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_13_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_13_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_14_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_14_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_15_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_15_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_16_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_16_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_17_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_17_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_18_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_18_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_19_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_19_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_1_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_1_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_20_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_20_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_21_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_23_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_24_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_24_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_25_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_25_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_26_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_26_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_27_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_27_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_28_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_28_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_29_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_29_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_2_CFG_reg_sel                 (),                                           
/* input  logic           */ .LPM_TREE_STATE_2_STATUS_reg_sel              (),                                           
/* input  logic           */ .LPM_TREE_STATE_30_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_30_STATUS_reg_sel             (),                                           
/* input  logic           */ .LPM_TREE_STATE_31_CFG_reg_sel                (),                                           
/* input  logic           */ .LPM_TREE_STATE_31_STATUS_reg_sel             (),                                           
/* output logic           */ .classifier_ecc_int                           (),                                           
/* output logic   [285:0] */ .classifier_em_a_delay_fifo_0_to_mem          (classifier_em_a_delay_fifo_0_to_mem),        
/* output logic   [285:0] */ .classifier_em_a_delay_fifo_1_to_mem          (classifier_em_a_delay_fifo_1_to_mem),        
/* output logic   [285:0] */ .classifier_em_a_delay_fifo_2_to_mem          (classifier_em_a_delay_fifo_2_to_mem),        
/* output logic   [285:0] */ .classifier_em_a_delay_fifo_3_to_mem          (classifier_em_a_delay_fifo_3_to_mem),        
/* output logic    [79:0] */ .classifier_em_a_hash_cfg_to_mem              (classifier_em_a_hash_cfg_to_mem),            
/* output logic   [104:0] */ .classifier_em_a_hash_lookup_to_mem           (classifier_em_a_hash_lookup_to_mem),         
/* output logic   [156:0] */ .classifier_em_a_hash_miss_to_mem             (classifier_em_a_hash_miss_to_mem),           
/* output logic    [91:0] */ .classifier_em_a_key_mask_0_to_mem            (classifier_em_a_key_mask_0_to_mem),          
/* output logic    [91:0] */ .classifier_em_a_key_mask_1_to_mem            (classifier_em_a_key_mask_1_to_mem),          
/* output logic    [91:0] */ .classifier_em_a_key_mask_2_to_mem            (classifier_em_a_key_mask_2_to_mem),          
/* output logic    [79:0] */ .classifier_em_b_hash_cfg_to_mem              (classifier_em_b_hash_cfg_to_mem),            
/* output logic   [101:0] */ .classifier_em_b_hash_lookup_to_mem           (classifier_em_b_hash_lookup_to_mem),         
/* output logic   [156:0] */ .classifier_em_b_hash_miss_to_mem             (classifier_em_b_hash_miss_to_mem),           
/* output logic    [91:0] */ .classifier_em_b_key_mask_to_mem              (classifier_em_b_key_mask_to_mem),            
/* output logic           */ .classifier_init_done                         (),                                           
/* output logic   [485:0] */ .classifier_lpm_key_cam_to_tcam               (classifier_lpm_key_cam_to_tcam),             
/* output logic   [323:0] */ .classifier_lpm_tree_state_0_to_mem           (classifier_lpm_tree_state_0_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_10_to_mem          (classifier_lpm_tree_state_10_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_11_to_mem          (classifier_lpm_tree_state_11_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_12_to_mem          (classifier_lpm_tree_state_12_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_13_to_mem          (classifier_lpm_tree_state_13_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_14_to_mem          (classifier_lpm_tree_state_14_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_15_to_mem          (classifier_lpm_tree_state_15_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_16_to_mem          (classifier_lpm_tree_state_16_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_17_to_mem          (classifier_lpm_tree_state_17_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_18_to_mem          (classifier_lpm_tree_state_18_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_19_to_mem          (classifier_lpm_tree_state_19_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_1_to_mem           (classifier_lpm_tree_state_1_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_20_to_mem          (classifier_lpm_tree_state_20_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_21_to_mem          (classifier_lpm_tree_state_21_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_22_to_mem          (classifier_lpm_tree_state_22_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_23_to_mem          (classifier_lpm_tree_state_23_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_24_to_mem          (classifier_lpm_tree_state_24_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_25_to_mem          (classifier_lpm_tree_state_25_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_26_to_mem          (classifier_lpm_tree_state_26_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_27_to_mem          (classifier_lpm_tree_state_27_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_28_to_mem          (classifier_lpm_tree_state_28_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_29_to_mem          (classifier_lpm_tree_state_29_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_2_to_mem           (classifier_lpm_tree_state_2_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_30_to_mem          (classifier_lpm_tree_state_30_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_31_to_mem          (classifier_lpm_tree_state_31_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_32_to_mem          (classifier_lpm_tree_state_32_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_33_to_mem          (classifier_lpm_tree_state_33_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_34_to_mem          (classifier_lpm_tree_state_34_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_35_to_mem          (classifier_lpm_tree_state_35_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_36_to_mem          (classifier_lpm_tree_state_36_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_37_to_mem          (classifier_lpm_tree_state_37_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_38_to_mem          (classifier_lpm_tree_state_38_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_39_to_mem          (classifier_lpm_tree_state_39_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_3_to_mem           (classifier_lpm_tree_state_3_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_40_to_mem          (classifier_lpm_tree_state_40_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_41_to_mem          (classifier_lpm_tree_state_41_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_42_to_mem          (classifier_lpm_tree_state_42_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_43_to_mem          (classifier_lpm_tree_state_43_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_44_to_mem          (classifier_lpm_tree_state_44_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_45_to_mem          (classifier_lpm_tree_state_45_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_46_to_mem          (classifier_lpm_tree_state_46_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_47_to_mem          (classifier_lpm_tree_state_47_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_48_to_mem          (classifier_lpm_tree_state_48_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_49_to_mem          (classifier_lpm_tree_state_49_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_4_to_mem           (classifier_lpm_tree_state_4_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_50_to_mem          (classifier_lpm_tree_state_50_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_51_to_mem          (classifier_lpm_tree_state_51_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_52_to_mem          (classifier_lpm_tree_state_52_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_53_to_mem          (classifier_lpm_tree_state_53_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_54_to_mem          (classifier_lpm_tree_state_54_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_55_to_mem          (classifier_lpm_tree_state_55_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_56_to_mem          (classifier_lpm_tree_state_56_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_57_to_mem          (classifier_lpm_tree_state_57_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_58_to_mem          (classifier_lpm_tree_state_58_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_59_to_mem          (classifier_lpm_tree_state_59_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_5_to_mem           (classifier_lpm_tree_state_5_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_60_to_mem          (classifier_lpm_tree_state_60_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_61_to_mem          (classifier_lpm_tree_state_61_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_62_to_mem          (classifier_lpm_tree_state_62_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_63_to_mem          (classifier_lpm_tree_state_63_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_64_to_mem          (classifier_lpm_tree_state_64_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_65_to_mem          (classifier_lpm_tree_state_65_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_66_to_mem          (classifier_lpm_tree_state_66_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_67_to_mem          (classifier_lpm_tree_state_67_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_68_to_mem          (classifier_lpm_tree_state_68_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_69_to_mem          (classifier_lpm_tree_state_69_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_6_to_mem           (classifier_lpm_tree_state_6_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_70_to_mem          (classifier_lpm_tree_state_70_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_74_to_mem          (classifier_lpm_tree_state_74_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_75_to_mem          (classifier_lpm_tree_state_75_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_76_to_mem          (classifier_lpm_tree_state_76_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_77_to_mem          (classifier_lpm_tree_state_77_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_78_to_mem          (classifier_lpm_tree_state_78_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_79_to_mem          (classifier_lpm_tree_state_79_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_7_to_mem           (classifier_lpm_tree_state_7_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_80_to_mem          (classifier_lpm_tree_state_80_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_81_to_mem          (classifier_lpm_tree_state_81_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_82_to_mem          (classifier_lpm_tree_state_82_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_83_to_mem          (classifier_lpm_tree_state_83_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_84_to_mem          (classifier_lpm_tree_state_84_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_85_to_mem          (classifier_lpm_tree_state_85_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_86_to_mem          (classifier_lpm_tree_state_86_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_87_to_mem          (classifier_lpm_tree_state_87_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_88_to_mem          (classifier_lpm_tree_state_88_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_89_to_mem          (classifier_lpm_tree_state_89_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_8_to_mem           (classifier_lpm_tree_state_8_to_mem),         
/* output logic   [323:0] */ .classifier_lpm_tree_state_90_to_mem          (classifier_lpm_tree_state_90_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_91_to_mem          (classifier_lpm_tree_state_91_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_92_to_mem          (classifier_lpm_tree_state_92_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_93_to_mem          (classifier_lpm_tree_state_93_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_94_to_mem          (classifier_lpm_tree_state_94_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_95_to_mem          (classifier_lpm_tree_state_95_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_9_to_mem           (classifier_lpm_tree_state_9_to_mem),         
/* output logic    [92:0] */ .classifier_map_domain_action0_to_mem         (classifier_map_domain_action0_to_mem),       
/* output logic    [92:0] */ .classifier_map_domain_action1_to_mem         (classifier_map_domain_action1_to_mem),       
/* output logic    [81:0] */ .classifier_map_domain_pol_cfg_to_mem         (classifier_map_domain_pol_cfg_to_mem),       
/* output logic    [89:0] */ .classifier_map_domain_profile_to_mem         (classifier_map_domain_profile_to_mem),       
/* output logic  [4434:0] */ .classifier_map_domain_tcam_to_tcam           (classifier_map_domain_tcam_to_tcam),         
/* output logic    [91:0] */ .classifier_map_dscp_tc_to_mem                (classifier_map_dscp_tc_to_mem),              
/* output logic    [89:0] */ .classifier_map_exp_tc_to_mem                 (classifier_map_exp_tc_to_mem),               
/* output logic    [87:0] */ .classifier_map_extract_0_to_mem              (classifier_map_extract_0_to_mem),            
/* output logic    [87:0] */ .classifier_map_extract_1_to_mem              (classifier_map_extract_1_to_mem),            
/* output logic    [87:0] */ .classifier_map_extract_2_to_mem              (classifier_map_extract_2_to_mem),            
/* output logic    [87:0] */ .classifier_map_ip_cfg_to_mem                 (classifier_map_ip_cfg_to_mem),               
/* output logic    [87:0] */ .classifier_map_ip_hi_to_mem                  (classifier_map_ip_hi_to_mem),                
/* output logic    [87:0] */ .classifier_map_ip_lo_to_mem                  (classifier_map_ip_lo_to_mem),                
/* output logic    [86:0] */ .classifier_map_l4_dst_to_mem                 (classifier_map_l4_dst_to_mem),               
/* output logic    [86:0] */ .classifier_map_l4_src_to_mem                 (classifier_map_l4_src_to_mem),               
/* output logic    [91:0] */ .classifier_map_len_limit_to_mem              (classifier_map_len_limit_to_mem),            
/* output logic   [152:0] */ .classifier_map_mac_to_mem                    (classifier_map_mac_to_mem),                  
/* output logic    [91:0] */ .classifier_map_port_cfg_to_mem               (classifier_map_port_cfg_to_mem),             
/* output logic    [85:0] */ .classifier_map_port_default_0_to_mem         (classifier_map_port_default_0_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_10_to_mem        (classifier_map_port_default_10_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_11_to_mem        (classifier_map_port_default_11_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_12_to_mem        (classifier_map_port_default_12_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_13_to_mem        (classifier_map_port_default_13_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_14_to_mem        (classifier_map_port_default_14_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_15_to_mem        (classifier_map_port_default_15_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_16_to_mem        (classifier_map_port_default_16_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_17_to_mem        (classifier_map_port_default_17_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_18_to_mem        (classifier_map_port_default_18_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_19_to_mem        (classifier_map_port_default_19_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_1_to_mem         (classifier_map_port_default_1_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_20_to_mem        (classifier_map_port_default_20_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_21_to_mem        (classifier_map_port_default_21_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_22_to_mem        (classifier_map_port_default_22_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_23_to_mem        (classifier_map_port_default_23_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_24_to_mem        (classifier_map_port_default_24_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_25_to_mem        (classifier_map_port_default_25_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_26_to_mem        (classifier_map_port_default_26_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_27_to_mem        (classifier_map_port_default_27_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_28_to_mem        (classifier_map_port_default_28_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_29_to_mem        (classifier_map_port_default_29_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_2_to_mem         (classifier_map_port_default_2_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_30_to_mem        (classifier_map_port_default_30_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_31_to_mem        (classifier_map_port_default_31_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_32_to_mem        (classifier_map_port_default_32_to_mem),      
/* output logic    [85:0] */ .classifier_map_port_default_3_to_mem         (classifier_map_port_default_3_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_4_to_mem         (classifier_map_port_default_4_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_5_to_mem         (classifier_map_port_default_5_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_6_to_mem         (classifier_map_port_default_6_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_7_to_mem         (classifier_map_port_default_7_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_8_to_mem         (classifier_map_port_default_8_to_mem),       
/* output logic    [85:0] */ .classifier_map_port_default_9_to_mem         (classifier_map_port_default_9_to_mem),       
/* output logic    [91:0] */ .classifier_map_port_to_mem                   (classifier_map_port_to_mem),                 
/* output logic    [87:0] */ .classifier_map_profile_action_to_mem         (classifier_map_profile_action_to_mem),       
/* output logic   [109:0] */ .classifier_map_profile_key0_to_mem           (classifier_map_profile_key0_to_mem),         
/* output logic   [109:0] */ .classifier_map_profile_key1_to_mem           (classifier_map_profile_key1_to_mem),         
/* output logic   [109:0] */ .classifier_map_profile_key_invert0_to_mem    (classifier_map_profile_key_invert0_to_mem),  
/* output logic   [109:0] */ .classifier_map_profile_key_invert1_to_mem    (classifier_map_profile_key_invert1_to_mem),  
/* output logic    [85:0] */ .classifier_map_prot_to_mem                   (classifier_map_prot_to_mem),                 
/* output logic    [89:0] */ .classifier_map_rewrite_0_to_mem              (classifier_map_rewrite_0_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_10_to_mem             (classifier_map_rewrite_10_to_mem),           
/* output logic    [89:0] */ .classifier_map_rewrite_11_to_mem             (classifier_map_rewrite_11_to_mem),           
/* output logic    [89:0] */ .classifier_map_rewrite_12_to_mem             (classifier_map_rewrite_12_to_mem),           
/* output logic    [89:0] */ .classifier_map_rewrite_13_to_mem             (classifier_map_rewrite_13_to_mem),           
/* output logic    [89:0] */ .classifier_map_rewrite_14_to_mem             (classifier_map_rewrite_14_to_mem),           
/* output logic    [89:0] */ .classifier_map_rewrite_15_to_mem             (classifier_map_rewrite_15_to_mem),           
/* output logic    [89:0] */ .classifier_map_rewrite_1_to_mem              (classifier_map_rewrite_1_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_2_to_mem              (classifier_map_rewrite_2_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_3_to_mem              (classifier_map_rewrite_3_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_4_to_mem              (classifier_map_rewrite_4_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_5_to_mem              (classifier_map_rewrite_5_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_6_to_mem              (classifier_map_rewrite_6_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_7_to_mem              (classifier_map_rewrite_7_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_8_to_mem              (classifier_map_rewrite_8_to_mem),            
/* output logic    [89:0] */ .classifier_map_rewrite_9_to_mem              (classifier_map_rewrite_9_to_mem),            
/* output logic    [87:0] */ .classifier_map_type_to_mem                   (classifier_map_type_to_mem),                 
/* output logic    [89:0] */ .classifier_map_vpri_tc_to_mem                (classifier_map_vpri_tc_to_mem),              
/* output logic    [89:0] */ .classifier_map_vpri_to_mem                   (classifier_map_vpri_to_mem),                 
/* output logic    [88:0] */ .classifier_wcm_action_cfg_0_to_mem           (classifier_wcm_action_cfg_0_to_mem),         
/* output logic    [88:0] */ .classifier_wcm_action_cfg_1_to_mem           (classifier_wcm_action_cfg_1_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_0_to_mem           (classifier_wcm_action_ram_0_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_10_to_mem          (classifier_wcm_action_ram_10_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_11_to_mem          (classifier_wcm_action_ram_11_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_12_to_mem          (classifier_wcm_action_ram_12_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_13_to_mem          (classifier_wcm_action_ram_13_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_14_to_mem          (classifier_wcm_action_ram_14_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_15_to_mem          (classifier_wcm_action_ram_15_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_16_to_mem          (classifier_wcm_action_ram_16_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_17_to_mem          (classifier_wcm_action_ram_17_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_18_to_mem          (classifier_wcm_action_ram_18_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_19_to_mem          (classifier_wcm_action_ram_19_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_1_to_mem           (classifier_wcm_action_ram_1_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_2_to_mem           (classifier_wcm_action_ram_2_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_3_to_mem           (classifier_wcm_action_ram_3_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_4_to_mem           (classifier_wcm_action_ram_4_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_5_to_mem           (classifier_wcm_action_ram_5_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_6_to_mem           (classifier_wcm_action_ram_6_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_7_to_mem           (classifier_wcm_action_ram_7_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_8_to_mem           (classifier_wcm_action_ram_8_to_mem),         
/* output logic    [90:0] */ .classifier_wcm_action_ram_9_to_mem           (classifier_wcm_action_ram_9_to_mem),         
/* output logic    [85:0] */ .classifier_wcm_data_path_buffer0_to_mem      (classifier_wcm_data_path_buffer0_to_mem),    
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_0_to_mem    (classifier_wcm_data_path_buffer1_0_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_10_to_mem   (classifier_wcm_data_path_buffer1_10_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_11_to_mem   (classifier_wcm_data_path_buffer1_11_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_12_to_mem   (classifier_wcm_data_path_buffer1_12_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_13_to_mem   (classifier_wcm_data_path_buffer1_13_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_14_to_mem   (classifier_wcm_data_path_buffer1_14_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_15_to_mem   (classifier_wcm_data_path_buffer1_15_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_16_to_mem   (classifier_wcm_data_path_buffer1_16_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_17_to_mem   (classifier_wcm_data_path_buffer1_17_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_18_to_mem   (classifier_wcm_data_path_buffer1_18_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_19_to_mem   (classifier_wcm_data_path_buffer1_19_to_mem), 
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_1_to_mem    (classifier_wcm_data_path_buffer1_1_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_2_to_mem    (classifier_wcm_data_path_buffer1_2_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_3_to_mem    (classifier_wcm_data_path_buffer1_3_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_4_to_mem    (classifier_wcm_data_path_buffer1_4_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_5_to_mem    (classifier_wcm_data_path_buffer1_5_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_6_to_mem    (classifier_wcm_data_path_buffer1_6_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_7_to_mem    (classifier_wcm_data_path_buffer1_7_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_8_to_mem    (classifier_wcm_data_path_buffer1_8_to_mem),  
/* output logic   [362:0] */ .classifier_wcm_data_path_buffer1_9_to_mem    (classifier_wcm_data_path_buffer1_9_to_mem),  
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_0_to_mem         (classifier_wcm_tcam_cfg_ram_0_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_10_to_mem        (classifier_wcm_tcam_cfg_ram_10_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_11_to_mem        (classifier_wcm_tcam_cfg_ram_11_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_12_to_mem        (classifier_wcm_tcam_cfg_ram_12_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_13_to_mem        (classifier_wcm_tcam_cfg_ram_13_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_14_to_mem        (classifier_wcm_tcam_cfg_ram_14_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_15_to_mem        (classifier_wcm_tcam_cfg_ram_15_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_16_to_mem        (classifier_wcm_tcam_cfg_ram_16_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_17_to_mem        (classifier_wcm_tcam_cfg_ram_17_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_18_to_mem        (classifier_wcm_tcam_cfg_ram_18_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_19_to_mem        (classifier_wcm_tcam_cfg_ram_19_to_mem),      
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_1_to_mem         (classifier_wcm_tcam_cfg_ram_1_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_2_to_mem         (classifier_wcm_tcam_cfg_ram_2_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_3_to_mem         (classifier_wcm_tcam_cfg_ram_3_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_4_to_mem         (classifier_wcm_tcam_cfg_ram_4_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_5_to_mem         (classifier_wcm_tcam_cfg_ram_5_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_6_to_mem         (classifier_wcm_tcam_cfg_ram_6_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_7_to_mem         (classifier_wcm_tcam_cfg_ram_7_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_8_to_mem         (classifier_wcm_tcam_cfg_ram_8_to_mem),       
/* output logic    [88:0] */ .classifier_wcm_tcam_cfg_ram_9_to_mem         (classifier_wcm_tcam_cfg_ram_9_to_mem),       
/* output logic  [1192:0] */ .classifier_wcm_tcam_to_tcam                  (),                                           
/* output logic           */ .em_a_delay_fifo_0_ecc_uncor_err              (),                                           
/* output logic           */ .em_a_delay_fifo_0_init_done                  (),                                           
/* output logic   [255:0] */ .em_a_delay_fifo_0_rd_data                    (),                                           
/* output logic           */ .em_a_delay_fifo_0_rd_valid                   (),                                           
/* output logic           */ .em_a_delay_fifo_1_ecc_uncor_err              (),                                           
/* output logic           */ .em_a_delay_fifo_1_init_done                  (),                                           
/* output logic   [255:0] */ .em_a_delay_fifo_1_rd_data                    (),                                           
/* output logic           */ .em_a_delay_fifo_1_rd_valid                   (),                                           
/* output logic           */ .em_a_delay_fifo_2_ecc_uncor_err              (),                                           
/* output logic           */ .em_a_delay_fifo_2_init_done                  (),                                           
/* output logic   [255:0] */ .em_a_delay_fifo_2_rd_data                    (),                                           
/* output logic           */ .em_a_delay_fifo_2_rd_valid                   (),                                           
/* output logic           */ .em_a_delay_fifo_3_ecc_uncor_err              (),                                           
/* output logic           */ .em_a_delay_fifo_3_init_done                  (),                                           
/* output logic   [255:0] */ .em_a_delay_fifo_3_rd_data                    (),                                           
/* output logic           */ .em_a_delay_fifo_3_rd_valid                   (),                                           
/* output logic           */ .em_a_hash_cfg_ecc_uncor_err                  (),                                           
/* output logic           */ .em_a_hash_cfg_init_done                      (),                                           
/* output logic    [52:0] */ .em_a_hash_cfg_rd_data                        (),                                           
/* output logic           */ .em_a_hash_cfg_rd_valid                       (),                                           
/* output logic           */ .em_a_hash_lookup_ecc_uncor_err               (),                                           
/* output logic           */ .em_a_hash_lookup_init_done                   (),                                           
/* output logic    [71:0] */ .em_a_hash_lookup_rd_data                     (),                                           
/* output logic           */ .em_a_hash_lookup_rd_valid                    (),                                           
/* output logic           */ .em_a_hash_miss_ecc_uncor_err                 (),                                           
/* output logic           */ .em_a_hash_miss_init_done                     (),                                           
/* output logic   [127:0] */ .em_a_hash_miss_rd_data                       (),                                           
/* output logic           */ .em_a_hash_miss_rd_valid                      (),                                           
/* output logic           */ .em_a_key_mask_0_ecc_uncor_err                (),                                           
/* output logic           */ .em_a_key_mask_0_init_done                    (),                                           
/* output logic    [63:0] */ .em_a_key_mask_0_rd_data                      (),                                           
/* output logic           */ .em_a_key_mask_0_rd_valid                     (),                                           
/* output logic           */ .em_a_key_mask_1_ecc_uncor_err                (),                                           
/* output logic           */ .em_a_key_mask_1_init_done                    (),                                           
/* output logic    [63:0] */ .em_a_key_mask_1_rd_data                      (),                                           
/* output logic           */ .em_a_key_mask_1_rd_valid                     (),                                           
/* output logic           */ .em_a_key_mask_2_ecc_uncor_err                (),                                           
/* output logic           */ .em_a_key_mask_2_init_done                    (),                                           
/* output logic    [63:0] */ .em_a_key_mask_2_rd_data                      (),                                           
/* output logic           */ .em_a_key_mask_2_rd_valid                     (),                                           
/* output logic           */ .em_b_hash_cfg_ecc_uncor_err                  (),                                           
/* output logic           */ .em_b_hash_cfg_init_done                      (),                                           
/* output logic    [52:0] */ .em_b_hash_cfg_rd_data                        (),                                           
/* output logic           */ .em_b_hash_cfg_rd_valid                       (),                                           
/* output logic           */ .em_b_hash_lookup_ecc_uncor_err               (),                                           
/* output logic           */ .em_b_hash_lookup_init_done                   (),                                           
/* output logic           */ .em_b_hash_miss_init_done                     (),                                           
/* output logic   [127:0] */ .em_b_hash_miss_rd_data                       (),                                           
/* output logic           */ .em_b_hash_miss_rd_valid                      (),                                           
/* output logic           */ .em_b_key_mask_ecc_uncor_err                  (),                                           
/* output logic           */ .em_b_key_mask_init_done                      (),                                           
/* output logic    [63:0] */ .em_b_key_mask_rd_data                        (),                                           
/* output logic           */ .em_b_key_mask_rd_valid                       (),                                           
/* output logic           */ .lpm_key_cam_ecc_uncor_err                    (),                                           
/* output logic           */ .lpm_key_cam_init_done                        (),                                           
/* output logic   [255:0] */ .lpm_key_cam_raw_hit_out                      (),                                           
/* output logic    [64:0] */ .lpm_key_cam_rd_data                          (),                                           
/* output logic     [7:0] */ .lpm_key_cam_rule_hit_num                     (),                                           
/* output logic           */ .lpm_key_cam_rule_hit_num_vld                 (),                                           
/* output logic           */ .lpm_key_cam_tcam_chk_rdy                     (),                                           
/* output logic           */ .lpm_key_cam_tcam_chk_valid                   (),                                           
/* output logic           */ .lpm_key_cam_tcam_rd_valid                    (),                                           
/* output logic           */ .lpm_key_cam_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .lpm_tree_state_0_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_0_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_0_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_0_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_10_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_10_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_10_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_10_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_11_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_11_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_11_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_11_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_12_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_12_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_12_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_12_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_13_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_13_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_13_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_13_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_14_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_14_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_14_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_14_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_15_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_15_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_15_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_15_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_16_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_16_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_16_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_16_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_17_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_17_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_17_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_17_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_18_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_18_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_18_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_18_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_19_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_19_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_19_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_19_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_1_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_1_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_1_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_1_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_20_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_20_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_20_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_20_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_21_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_21_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_21_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_21_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_22_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_22_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_22_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_22_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_23_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_23_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_23_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_23_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_24_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_24_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_24_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_24_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_26_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_26_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_26_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_26_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_27_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_27_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_27_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_27_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_28_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_28_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_28_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_28_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_29_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_29_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_29_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_29_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_2_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_2_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_2_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_2_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_30_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_30_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_30_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_30_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_31_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_31_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_31_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_31_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_32_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_32_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_32_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_32_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_33_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_33_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_33_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_33_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_34_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_34_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_34_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_34_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_35_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_35_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_35_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_35_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_36_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_36_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_36_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_36_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_37_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_37_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_37_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_37_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_38_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_38_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_38_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_38_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_39_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_39_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_39_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_39_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_3_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_3_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_3_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_3_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_40_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_40_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_40_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_40_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_41_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_41_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_41_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_41_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_42_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_42_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_42_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_42_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_43_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_43_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_43_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_43_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_45_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_45_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_45_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_45_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_46_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_46_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_46_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_46_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_47_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_47_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_47_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_47_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_48_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_48_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_48_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_48_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_49_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_49_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_49_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_49_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_4_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_4_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_4_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_4_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_50_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_50_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_50_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_50_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_51_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_51_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_51_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_51_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_52_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_52_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_52_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_52_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_53_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_53_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_53_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_53_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_54_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_54_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_54_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_54_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_55_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_55_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_55_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_55_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_56_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_56_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_56_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_56_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_57_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_57_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_57_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_57_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_58_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_58_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_58_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_58_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_59_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_59_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_59_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_59_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_5_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_5_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_5_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_5_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_60_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_60_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_60_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_60_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_61_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_61_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_61_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_61_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_62_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_62_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_62_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_62_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_63_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_63_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_63_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_63_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_64_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_65_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_65_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_65_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_66_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_66_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_66_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_66_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_67_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_67_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_67_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_67_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_68_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_68_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_68_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_68_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_69_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_69_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_69_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_69_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_6_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_6_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_6_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_6_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_70_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_70_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_70_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_70_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_71_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_71_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_71_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_71_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_72_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_72_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_72_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_72_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_73_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_73_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_73_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_73_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_74_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_74_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_74_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_74_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_75_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_75_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_75_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_75_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_76_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_76_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_76_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_76_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_77_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_77_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_77_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_77_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_78_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_78_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_78_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_78_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_79_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_79_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_79_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_79_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_7_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_7_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_7_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_7_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_80_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_80_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_80_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_80_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_81_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_81_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_81_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_81_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_82_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_82_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_82_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_82_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_83_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_84_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_84_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_84_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_85_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_85_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_85_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_85_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_86_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_86_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_86_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_86_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_87_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_87_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_87_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_87_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_88_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_88_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_88_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_88_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_89_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_89_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_89_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_89_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_8_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_8_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_8_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_8_rd_valid                    (),                                           
/* output logic           */ .lpm_tree_state_90_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_90_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_90_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_90_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_91_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_91_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_91_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_91_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_92_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_92_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_92_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_92_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_93_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_93_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_93_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_93_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_94_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_94_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_94_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_94_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_95_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_95_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_95_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_95_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_9_ecc_uncor_err               (),                                           
/* output logic           */ .lpm_tree_state_9_init_done                   (),                                           
/* output logic   [295:0] */ .lpm_tree_state_9_rd_data                     (),                                           
/* output logic           */ .lpm_tree_state_9_rd_valid                    (),                                           
/* output logic           */ .map_domain_action0_ecc_uncor_err             (),                                           
/* output logic           */ .map_domain_action0_init_done                 (),                                           
/* output logic    [63:0] */ .map_domain_action0_rd_data                   (),                                           
/* output logic           */ .map_domain_action0_rd_valid                  (),                                           
/* output logic           */ .map_domain_action1_ecc_uncor_err             (),                                           
/* output logic           */ .map_domain_action1_init_done                 (),                                           
/* output logic    [63:0] */ .map_domain_action1_rd_data                   (),                                           
/* output logic           */ .map_domain_action1_rd_valid                  (),                                           
/* output logic           */ .map_domain_pol_cfg_ecc_uncor_err             (),                                           
/* output logic           */ .map_domain_pol_cfg_init_done                 (),                                           
/* output logic    [63:0] */ .map_domain_pol_cfg_rd_data                   (),                                           
/* output logic           */ .map_domain_pol_cfg_rd_valid                  (),                                           
/* output logic           */ .map_domain_profile_ecc_uncor_err             (),                                           
/* output logic           */ .map_domain_profile_init_done                 (),                                           
/* output logic    [63:0] */ .map_domain_profile_rd_data                   (),                                           
/* output logic           */ .map_domain_profile_rd_valid                  (),                                           
/* output logic           */ .map_domain_tcam_ecc_uncor_err                (),                                           
/* output logic           */ .map_domain_tcam_init_done                    (),                                           
/* output logic  [4095:0] */ .map_domain_tcam_raw_hit_out                  (),                                           
/* output logic    [79:0] */ .map_domain_tcam_rd_data                      (),                                           
/* output logic    [11:0] */ .map_domain_tcam_rule_hit_num                 (),                                           
/* output logic           */ .map_domain_tcam_rule_hit_num_vld             (),                                           
/* output logic           */ .map_domain_tcam_tcam_chk_rdy                 (),                                           
/* output logic           */ .map_domain_tcam_tcam_chk_valid               (),                                           
/* output logic           */ .map_domain_tcam_tcam_rd_valid                (),                                           
/* output logic           */ .map_domain_tcam_tcam_rdwr_rdy                (),                                           
/* output logic           */ .map_dscp_tc_ecc_uncor_err                    (),                                           
/* output logic           */ .map_dscp_tc_init_done                        (),                                           
/* output logic    [63:0] */ .map_dscp_tc_rd_data                          (),                                           
/* output logic           */ .map_dscp_tc_rd_valid                         (),                                           
/* output logic           */ .map_exp_tc_rd_valid                          (),                                           
/* output logic           */ .map_extract_0_ecc_uncor_err                  (),                                           
/* output logic           */ .map_extract_0_init_done                      (),                                           
/* output logic    [63:0] */ .map_extract_0_rd_data                        (),                                           
/* output logic           */ .map_extract_0_rd_valid                       (),                                           
/* output logic           */ .map_extract_1_ecc_uncor_err                  (),                                           
/* output logic           */ .map_extract_1_init_done                      (),                                           
/* output logic    [63:0] */ .map_extract_1_rd_data                        (),                                           
/* output logic           */ .map_extract_1_rd_valid                       (),                                           
/* output logic           */ .map_extract_2_ecc_uncor_err                  (),                                           
/* output logic           */ .map_extract_2_init_done                      (),                                           
/* output logic    [63:0] */ .map_extract_2_rd_data                        (),                                           
/* output logic           */ .map_extract_2_rd_valid                       (),                                           
/* output logic           */ .map_ip_cfg_ecc_uncor_err                     (),                                           
/* output logic           */ .map_ip_cfg_init_done                         (),                                           
/* output logic    [63:0] */ .map_ip_cfg_rd_data                           (),                                           
/* output logic           */ .map_ip_cfg_rd_valid                          (),                                           
/* output logic           */ .map_ip_hi_ecc_uncor_err                      (),                                           
/* output logic           */ .map_ip_hi_init_done                          (),                                           
/* output logic    [63:0] */ .map_ip_hi_rd_data                            (),                                           
/* output logic           */ .map_ip_hi_rd_valid                           (),                                           
/* output logic           */ .map_ip_lo_ecc_uncor_err                      (),                                           
/* output logic           */ .map_ip_lo_init_done                          (),                                           
/* output logic    [63:0] */ .map_ip_lo_rd_data                            (),                                           
/* output logic           */ .map_ip_lo_rd_valid                           (),                                           
/* output logic           */ .map_l4_dst_ecc_uncor_err                     (),                                           
/* output logic           */ .map_l4_dst_init_done                         (),                                           
/* output logic    [63:0] */ .map_l4_dst_rd_data                           (),                                           
/* output logic           */ .map_l4_dst_rd_valid                          (),                                           
/* output logic           */ .map_l4_src_ecc_uncor_err                     (),                                           
/* output logic           */ .map_l4_src_init_done                         (),                                           
/* output logic    [63:0] */ .map_l4_src_rd_data                           (),                                           
/* output logic           */ .map_l4_src_rd_valid                          (),                                           
/* output logic           */ .map_len_limit_ecc_uncor_err                  (),                                           
/* output logic           */ .map_len_limit_init_done                      (),                                           
/* output logic    [63:0] */ .map_len_limit_rd_data                        (),                                           
/* output logic           */ .map_len_limit_rd_valid                       (),                                           
/* output logic           */ .map_mac_ecc_uncor_err                        (),                                           
/* output logic           */ .map_mac_init_done                            (),                                           
/* output logic   [127:0] */ .map_mac_rd_data                              (),                                           
/* output logic           */ .map_mac_rd_valid                             (),                                           
/* output logic           */ .map_port_cfg_ecc_uncor_err                   (),                                           
/* output logic           */ .map_port_cfg_init_done                       (),                                           
/* output logic    [63:0] */ .map_port_cfg_rd_data                         (),                                           
/* output logic           */ .map_port_cfg_rd_valid                        (),                                           
/* output logic           */ .map_port_default_0_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_0_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_0_rd_data                   (),                                           
/* output logic           */ .map_port_default_0_rd_valid                  (),                                           
/* output logic           */ .map_port_default_10_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_10_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_10_rd_data                  (),                                           
/* output logic           */ .map_port_default_10_rd_valid                 (),                                           
/* output logic           */ .map_port_default_11_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_11_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_11_rd_data                  (),                                           
/* output logic           */ .map_port_default_11_rd_valid                 (),                                           
/* output logic           */ .map_port_default_12_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_12_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_12_rd_data                  (),                                           
/* output logic           */ .map_port_default_12_rd_valid                 (),                                           
/* output logic           */ .map_port_default_13_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_13_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_13_rd_data                  (),                                           
/* output logic           */ .map_port_default_13_rd_valid                 (),                                           
/* output logic           */ .map_port_default_14_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_14_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_14_rd_data                  (),                                           
/* output logic           */ .map_port_default_14_rd_valid                 (),                                           
/* output logic           */ .map_port_default_15_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_15_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_15_rd_data                  (),                                           
/* output logic           */ .map_port_default_15_rd_valid                 (),                                           
/* output logic           */ .map_port_default_16_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_16_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_16_rd_data                  (),                                           
/* output logic           */ .map_port_default_16_rd_valid                 (),                                           
/* output logic           */ .map_port_default_17_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_17_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_17_rd_data                  (),                                           
/* output logic           */ .map_port_default_17_rd_valid                 (),                                           
/* output logic           */ .map_port_default_19_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_19_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_19_rd_data                  (),                                           
/* output logic           */ .map_port_default_19_rd_valid                 (),                                           
/* output logic           */ .map_port_default_1_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_1_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_1_rd_data                   (),                                           
/* output logic           */ .map_port_default_1_rd_valid                  (),                                           
/* output logic           */ .map_port_default_20_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_20_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_20_rd_data                  (),                                           
/* output logic           */ .map_port_default_20_rd_valid                 (),                                           
/* output logic           */ .map_port_default_21_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_21_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_21_rd_data                  (),                                           
/* output logic           */ .map_port_default_21_rd_valid                 (),                                           
/* output logic           */ .map_port_default_22_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_22_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_22_rd_data                  (),                                           
/* output logic           */ .map_port_default_22_rd_valid                 (),                                           
/* output logic           */ .map_port_default_23_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_23_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_23_rd_data                  (),                                           
/* output logic           */ .map_port_default_23_rd_valid                 (),                                           
/* output logic           */ .map_port_default_24_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_24_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_24_rd_data                  (),                                           
/* output logic           */ .map_port_default_24_rd_valid                 (),                                           
/* output logic           */ .map_port_default_25_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_25_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_25_rd_data                  (),                                           
/* output logic           */ .map_port_default_25_rd_valid                 (),                                           
/* output logic           */ .map_port_default_26_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_26_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_26_rd_data                  (),                                           
/* output logic           */ .map_port_default_26_rd_valid                 (),                                           
/* output logic           */ .map_port_default_27_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_27_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_27_rd_data                  (),                                           
/* output logic           */ .map_port_default_27_rd_valid                 (),                                           
/* output logic           */ .map_port_default_28_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_28_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_28_rd_data                  (),                                           
/* output logic           */ .map_port_default_28_rd_valid                 (),                                           
/* output logic           */ .map_port_default_29_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_29_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_29_rd_data                  (),                                           
/* output logic           */ .map_port_default_29_rd_valid                 (),                                           
/* output logic           */ .map_port_default_2_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_2_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_2_rd_data                   (),                                           
/* output logic           */ .map_port_default_2_rd_valid                  (),                                           
/* output logic           */ .map_port_default_30_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_30_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_30_rd_data                  (),                                           
/* output logic           */ .map_port_default_30_rd_valid                 (),                                           
/* output logic           */ .map_port_default_31_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_31_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_31_rd_data                  (),                                           
/* output logic           */ .map_port_default_31_rd_valid                 (),                                           
/* output logic           */ .map_port_default_32_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_32_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_32_rd_data                  (),                                           
/* output logic           */ .map_port_default_32_rd_valid                 (),                                           
/* output logic           */ .map_port_default_3_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_3_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_3_rd_data                   (),                                           
/* output logic           */ .map_port_default_3_rd_valid                  (),                                           
/* output logic           */ .map_port_default_4_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_4_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_4_rd_data                   (),                                           
/* output logic           */ .map_port_default_4_rd_valid                  (),                                           
/* output logic           */ .map_port_default_5_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_5_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_5_rd_data                   (),                                           
/* output logic           */ .map_port_default_5_rd_valid                  (),                                           
/* output logic           */ .map_port_default_6_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_6_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_6_rd_data                   (),                                           
/* output logic           */ .map_port_default_6_rd_valid                  (),                                           
/* output logic           */ .map_port_default_7_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_7_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_7_rd_data                   (),                                           
/* output logic           */ .map_port_default_7_rd_valid                  (),                                           
/* output logic           */ .map_port_default_9_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_9_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_9_rd_data                   (),                                           
/* output logic           */ .map_port_default_9_rd_valid                  (),                                           
/* output logic           */ .map_port_ecc_uncor_err                       (),                                           
/* output logic           */ .map_port_init_done                           (),                                           
/* output logic    [63:0] */ .map_port_rd_data                             (),                                           
/* output logic           */ .map_port_rd_valid                            (),                                           
/* output logic           */ .map_profile_action_ecc_uncor_err             (),                                           
/* output logic           */ .map_profile_action_init_done                 (),                                           
/* output logic    [63:0] */ .map_profile_action_rd_data                   (),                                           
/* output logic           */ .map_profile_action_rd_valid                  (),                                           
/* output logic           */ .map_profile_key0_ecc_uncor_err               (),                                           
/* output logic           */ .map_profile_key0_init_done                   (),                                           
/* output logic    [79:0] */ .map_profile_key0_rd_data                     (),                                           
/* output logic           */ .map_profile_key0_rd_valid                    (),                                           
/* output logic           */ .map_profile_key1_ecc_uncor_err               (),                                           
/* output logic           */ .map_profile_key1_init_done                   (),                                           
/* output logic    [79:0] */ .map_profile_key1_rd_data                     (),                                           
/* output logic           */ .map_profile_key1_rd_valid                    (),                                           
/* output logic           */ .map_profile_key_invert0_ecc_uncor_err        (),                                           
/* output logic           */ .map_profile_key_invert0_init_done            (),                                           
/* output logic    [79:0] */ .map_profile_key_invert0_rd_data              (),                                           
/* output logic           */ .map_profile_key_invert0_rd_valid             (),                                           
/* output logic           */ .map_profile_key_invert1_ecc_uncor_err        (),                                           
/* output logic           */ .map_profile_key_invert1_init_done            (),                                           
/* output logic    [79:0] */ .map_profile_key_invert1_rd_data              (),                                           
/* output logic           */ .map_profile_key_invert1_rd_valid             (),                                           
/* output logic           */ .map_prot_ecc_uncor_err                       (),                                           
/* output logic           */ .map_prot_init_done                           (),                                           
/* output logic    [63:0] */ .map_prot_rd_data                             (),                                           
/* output logic           */ .map_prot_rd_valid                            (),                                           
/* output logic           */ .map_rewrite_0_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_0_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_0_rd_data                        (),                                           
/* output logic           */ .map_rewrite_0_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_10_ecc_uncor_err                 (),                                           
/* output logic           */ .map_rewrite_10_init_done                     (),                                           
/* output logic    [63:0] */ .map_rewrite_10_rd_data                       (),                                           
/* output logic           */ .map_rewrite_10_rd_valid                      (),                                           
/* output logic           */ .map_rewrite_11_ecc_uncor_err                 (),                                           
/* output logic           */ .map_rewrite_11_init_done                     (),                                           
/* output logic    [63:0] */ .map_rewrite_11_rd_data                       (),                                           
/* output logic           */ .map_rewrite_11_rd_valid                      (),                                           
/* output logic           */ .map_rewrite_12_ecc_uncor_err                 (),                                           
/* output logic           */ .map_rewrite_12_init_done                     (),                                           
/* output logic    [63:0] */ .map_rewrite_12_rd_data                       (),                                           
/* output logic           */ .map_rewrite_12_rd_valid                      (),                                           
/* output logic           */ .map_rewrite_13_ecc_uncor_err                 (),                                           
/* output logic           */ .map_rewrite_13_init_done                     (),                                           
/* output logic    [63:0] */ .map_rewrite_13_rd_data                       (),                                           
/* output logic           */ .map_rewrite_13_rd_valid                      (),                                           
/* output logic           */ .map_rewrite_14_ecc_uncor_err                 (),                                           
/* output logic           */ .map_rewrite_14_init_done                     (),                                           
/* output logic    [63:0] */ .map_rewrite_14_rd_data                       (),                                           
/* output logic           */ .map_rewrite_14_rd_valid                      (),                                           
/* output logic           */ .map_rewrite_15_ecc_uncor_err                 (),                                           
/* output logic           */ .map_rewrite_15_init_done                     (),                                           
/* output logic    [63:0] */ .map_rewrite_15_rd_data                       (),                                           
/* output logic           */ .map_rewrite_15_rd_valid                      (),                                           
/* output logic           */ .map_rewrite_1_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_1_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_1_rd_data                        (),                                           
/* output logic           */ .map_rewrite_1_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_2_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_2_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_2_rd_data                        (),                                           
/* output logic           */ .map_rewrite_2_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_3_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_3_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_3_rd_data                        (),                                           
/* output logic           */ .map_rewrite_3_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_4_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_4_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_4_rd_data                        (),                                           
/* output logic           */ .map_rewrite_4_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_5_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_5_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_5_rd_data                        (),                                           
/* output logic           */ .map_rewrite_5_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_6_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_7_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_7_rd_data                        (),                                           
/* output logic           */ .map_rewrite_7_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_8_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_8_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_8_rd_data                        (),                                           
/* output logic           */ .map_rewrite_8_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_9_ecc_uncor_err                  (),                                           
/* output logic           */ .map_rewrite_9_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_9_rd_data                        (),                                           
/* output logic           */ .map_rewrite_9_rd_valid                       (),                                           
/* output logic           */ .map_type_ecc_uncor_err                       (),                                           
/* output logic           */ .map_type_init_done                           (),                                           
/* output logic    [63:0] */ .map_type_rd_data                             (),                                           
/* output logic           */ .map_type_rd_valid                            (),                                           
/* output logic           */ .map_vpri_ecc_uncor_err                       (),                                           
/* output logic           */ .map_vpri_init_done                           (),                                           
/* output logic    [63:0] */ .map_vpri_rd_data                             (),                                           
/* output logic           */ .map_vpri_rd_valid                            (),                                           
/* output logic           */ .map_vpri_tc_ecc_uncor_err                    (),                                           
/* output logic           */ .map_vpri_tc_init_done                        (),                                           
/* output logic    [63:0] */ .map_vpri_tc_rd_data                          (),                                           
/* output logic           */ .map_vpri_tc_rd_valid                         (),                                           
/* output logic           */ .unified_regs_ack                             (),                                           
/* output logic    [31:0] */ .unified_regs_rd_data                         (),                                           
/* output logic           */ .wcm_action_cfg_0_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_cfg_0_init_done                   (),                                           
/* output logic    [59:0] */ .wcm_action_cfg_0_rd_data                     (),                                           
/* output logic           */ .wcm_action_cfg_0_rd_valid                    (),                                           
/* output logic           */ .wcm_action_cfg_1_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_cfg_1_init_done                   (),                                           
/* output logic    [59:0] */ .wcm_action_cfg_1_rd_data                     (),                                           
/* output logic           */ .wcm_action_cfg_1_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_0_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_0_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_0_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_0_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_10_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_10_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_10_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_10_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_11_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_11_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_11_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_11_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_12_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_12_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_12_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_12_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_13_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_13_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_13_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_13_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_14_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_14_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_14_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_14_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_15_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_15_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_15_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_15_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_16_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_16_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_16_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_16_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_17_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_17_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_17_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_17_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_18_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_18_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_18_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_18_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_19_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_19_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_19_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_19_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_1_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_1_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_1_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_20_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_21_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_21_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_21_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_21_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_22_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_22_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_22_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_22_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_23_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_23_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_23_rd_data                    (),                                           
/* output logic           */ .wcm_action_ram_23_rd_valid                   (),                                           
/* output logic           */ .wcm_action_ram_2_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_2_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_2_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_2_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_3_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_3_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_3_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_3_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_4_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_4_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_4_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_4_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_5_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_5_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_5_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_5_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_6_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_6_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_6_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_6_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_7_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_7_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_7_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_7_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_8_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_8_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_8_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_8_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_9_ecc_uncor_err               (),                                           
/* output logic           */ .wcm_action_ram_9_init_done                   (),                                           
/* output logic    [63:0] */ .wcm_action_ram_9_rd_data                     (),                                           
/* output logic           */ .wcm_action_ram_9_rd_valid                    (),                                           
/* output logic           */ .wcm_data_path_buffer0_ecc_uncor_err          (),                                           
/* output logic           */ .wcm_data_path_buffer0_init_done              (),                                           
/* output logic    [63:0] */ .wcm_data_path_buffer0_rd_data                (),                                           
/* output logic           */ .wcm_data_path_buffer0_rd_valid               (),                                           
/* output logic           */ .wcm_data_path_buffer1_0_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_0_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_0_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_0_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_10_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_10_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_10_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_10_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_11_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_11_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_11_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_11_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_12_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_12_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_12_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_12_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_13_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_13_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_13_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_13_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_14_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_14_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_14_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_14_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_15_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_15_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_15_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_15_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_16_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_16_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_16_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_16_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_17_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_17_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_17_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_17_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_19_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_19_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_19_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_19_rd_valid            (),                                           
/* output logic           */ .wcm_data_path_buffer1_1_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_1_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_1_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_1_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_2_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_2_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_2_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_2_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_3_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_3_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_3_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_3_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_4_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_4_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_4_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_4_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_5_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_5_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_5_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_5_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_6_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_6_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_6_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_6_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_7_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_7_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_7_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_7_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_8_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_8_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_8_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_8_rd_valid             (),                                           
/* output logic           */ .wcm_data_path_buffer1_9_ecc_uncor_err        (),                                           
/* output logic           */ .wcm_data_path_buffer1_9_init_done            (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_9_rd_data              (),                                           
/* output logic           */ .wcm_data_path_buffer1_9_rd_valid             (),                                           
/* output logic           */ .wcm_tcam_0_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_0_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_0_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_0_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_0_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_0_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_0_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_0_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_0_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_0_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_10_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_10_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_10_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_10_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_10_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_10_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_10_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_10_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_10_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_10_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_11_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_11_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_11_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_11_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_11_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_11_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_11_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_11_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_11_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_11_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_12_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_12_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_12_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_12_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_12_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_12_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_12_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_12_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_12_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_12_tcam_rdwr_rdy                    (),                                           
/* output logic     [9:0] */ .wcm_tcam_13_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_13_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_13_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_13_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_13_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_13_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_14_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_14_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_14_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_14_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_14_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_14_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_14_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_14_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_14_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_14_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_15_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_15_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_15_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_15_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_15_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_15_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_15_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_15_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_15_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_15_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_16_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_16_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_16_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_16_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_16_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_16_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_16_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_16_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_16_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_16_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_17_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_17_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_17_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_17_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_17_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_17_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_17_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_17_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_17_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_17_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_18_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_18_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_18_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_18_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_18_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_18_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_18_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_18_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_18_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_18_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_19_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_19_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_19_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_19_rd_data                          (),                                           
/* output logic     [9:0] */ .wcm_tcam_19_rule_hit_num                     (),                                           
/* output logic           */ .wcm_tcam_19_rule_hit_num_vld                 (),                                           
/* output logic           */ .wcm_tcam_19_tcam_chk_rdy                     (),                                           
/* output logic           */ .wcm_tcam_19_tcam_chk_valid                   (),                                           
/* output logic           */ .wcm_tcam_19_tcam_rd_valid                    (),                                           
/* output logic           */ .wcm_tcam_19_tcam_rdwr_rdy                    (),                                           
/* output logic           */ .wcm_tcam_1_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_1_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_1_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_1_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_1_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_1_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_1_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_1_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_1_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_1_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_2_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_2_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_2_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_2_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_2_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_2_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_2_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_2_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_2_tcam_rd_valid                     (),                                           
/* output logic  [1023:0] */ .wcm_tcam_3_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_3_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_3_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_3_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_3_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_3_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_3_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_3_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_4_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_4_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_4_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_4_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_4_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_4_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_4_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_4_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_4_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_4_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_5_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_5_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_5_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_5_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_5_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_5_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_5_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_5_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_5_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_5_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_6_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_6_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_6_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_6_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_6_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_6_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_6_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_6_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_6_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_6_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_7_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_7_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_7_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_7_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_7_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_7_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_7_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_7_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_7_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_7_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_8_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_8_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_8_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_8_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_8_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_8_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_8_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_8_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_8_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_8_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_9_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_9_init_done                         (),                                           
/* output logic  [1023:0] */ .wcm_tcam_9_raw_hit_out                       (),                                           
/* output logic    [39:0] */ .wcm_tcam_9_rd_data                           (),                                           
/* output logic     [9:0] */ .wcm_tcam_9_rule_hit_num                      (),                                           
/* output logic           */ .wcm_tcam_9_rule_hit_num_vld                  (),                                           
/* output logic           */ .wcm_tcam_9_tcam_chk_rdy                      (),                                           
/* output logic           */ .wcm_tcam_9_tcam_chk_valid                    (),                                           
/* output logic           */ .wcm_tcam_9_tcam_rd_valid                     (),                                           
/* output logic           */ .wcm_tcam_9_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_0_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_0_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_0_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_0_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_10_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_10_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_10_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_10_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_11_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_11_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_11_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_11_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_12_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_13_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_13_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_13_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_14_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_14_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_14_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_14_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_15_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_15_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_15_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_15_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_16_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_16_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_16_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_16_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_17_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_17_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_17_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_17_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_18_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_18_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_18_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_18_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_19_ecc_uncor_err            (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_19_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_19_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_19_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_1_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_1_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_1_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_1_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_2_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_2_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_2_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_2_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_3_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_3_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_3_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_3_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_4_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_4_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_4_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_4_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_5_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_5_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_5_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_5_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_6_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_6_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_6_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_6_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_7_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_7_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_7_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_7_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_8_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_8_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_8_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_8_rd_valid                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_9_ecc_uncor_err             (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_9_init_done                 (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_9_rd_data                   (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_9_rd_valid                  (),                                           
/* output logic   [323:0] */ .classifier_lpm_tree_state_71_to_mem          (classifier_lpm_tree_state_71_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_72_to_mem          (classifier_lpm_tree_state_72_to_mem),        
/* output logic   [323:0] */ .classifier_lpm_tree_state_73_to_mem          (classifier_lpm_tree_state_73_to_mem),        
/* output logic           */ .lpm_tree_state_64_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_64_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_64_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_65_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_25_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_25_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_25_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_25_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_44_ecc_uncor_err              (),                                           
/* output logic           */ .lpm_tree_state_44_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_44_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_44_rd_valid                   (),                                           
/* output logic    [90:0] */ .classifier_wcm_action_ram_20_to_mem          (classifier_wcm_action_ram_20_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_21_to_mem          (classifier_wcm_action_ram_21_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_22_to_mem          (classifier_wcm_action_ram_22_to_mem),        
/* output logic    [90:0] */ .classifier_wcm_action_ram_23_to_mem          (classifier_wcm_action_ram_23_to_mem),        
/* output logic           */ .wcm_tcam_2_tcam_rdwr_rdy                     (),                                           
/* output logic           */ .wcm_tcam_3_ecc_uncor_err                     (),                                           
/* output logic           */ .wcm_tcam_3_init_done                         (),                                           
/* output logic           */ .wcm_data_path_buffer1_18_ecc_uncor_err       (),                                           
/* output logic           */ .wcm_data_path_buffer1_18_init_done           (),                                           
/* output logic   [334:0] */ .wcm_data_path_buffer1_18_rd_data             (),                                           
/* output logic           */ .wcm_data_path_buffer1_18_rd_valid            (),                                           
/* output logic           */ .wcm_tcam_13_ecc_uncor_err                    (),                                           
/* output logic           */ .wcm_tcam_13_init_done                        (),                                           
/* output logic  [1023:0] */ .wcm_tcam_13_raw_hit_out                      (),                                           
/* output logic    [39:0] */ .wcm_tcam_13_rd_data                          (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_12_init_done                (),                                           
/* output logic    [61:0] */ .wcm_tcam_cfg_ram_12_rd_data                  (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_12_rd_valid                 (),                                           
/* output logic           */ .wcm_tcam_cfg_ram_13_ecc_uncor_err            (),                                           
/* output logic           */ .lpm_tree_state_83_init_done                  (),                                           
/* output logic   [295:0] */ .lpm_tree_state_83_rd_data                    (),                                           
/* output logic           */ .lpm_tree_state_83_rd_valid                   (),                                           
/* output logic           */ .lpm_tree_state_84_ecc_uncor_err              (),                                           
/* output logic           */ .map_exp_tc_ecc_uncor_err                     (),                                           
/* output logic           */ .map_exp_tc_init_done                         (),                                           
/* output logic    [63:0] */ .map_exp_tc_rd_data                           (),                                           
/* output logic    [71:0] */ .em_b_hash_lookup_rd_data                     (),                                           
/* output logic           */ .em_b_hash_lookup_rd_valid                    (),                                           
/* output logic           */ .em_b_hash_miss_ecc_uncor_err                 (),                                           
/* output logic           */ .map_rewrite_6_init_done                      (),                                           
/* output logic    [63:0] */ .map_rewrite_6_rd_data                        (),                                           
/* output logic           */ .map_rewrite_6_rd_valid                       (),                                           
/* output logic           */ .map_rewrite_7_ecc_uncor_err                  (),                                           
/* output logic           */ .wcm_action_ram_1_rd_valid                    (),                                           
/* output logic           */ .wcm_action_ram_20_ecc_uncor_err              (),                                           
/* output logic           */ .wcm_action_ram_20_init_done                  (),                                           
/* output logic    [63:0] */ .wcm_action_ram_20_rd_data                    (),                                           
/* output logic           */ .map_port_default_18_ecc_uncor_err            (),                                           
/* output logic           */ .map_port_default_18_init_done                (),                                           
/* output logic    [63:0] */ .map_port_default_18_rd_data                  (),                                           
/* output logic           */ .map_port_default_18_rd_valid                 (),                                           
/* output logic           */ .map_port_default_8_ecc_uncor_err             (),                                           
/* output logic           */ .map_port_default_8_init_done                 (),                                           
/* output logic    [63:0] */ .map_port_default_8_rd_data                   (),                                           
/* output logic           */ .map_port_default_8_rd_valid                  ());                                           
// End of module classifier_shells_wrapper from classifier_shells_wrapper


// module classifier_ff_mems    from classifier_ff_mems using classifier_ff_mems.map 
classifier_ff_mems    classifier_ff_mems(
/* input  logic         */ .car_raw_lan_power_good_with_byprst           (),                                           
/* input  logic         */ .cclk                                         (cclk),                                       
/* input  logic  [79:0] */ .classifier_em_a_hash_cfg_to_mem              (classifier_em_a_hash_cfg_to_mem),            
/* input  logic  [79:0] */ .classifier_em_b_hash_cfg_to_mem              (classifier_em_b_hash_cfg_to_mem),            
/* input  logic  [81:0] */ .classifier_map_domain_pol_cfg_to_mem         (classifier_map_domain_pol_cfg_to_mem),       
/* input  logic  [89:0] */ .classifier_map_exp_tc_to_mem                 (classifier_map_exp_tc_to_mem),               
/* input  logic  [87:0] */ .classifier_map_extract_0_to_mem              (classifier_map_extract_0_to_mem),            
/* input  logic  [87:0] */ .classifier_map_extract_1_to_mem              (classifier_map_extract_1_to_mem),            
/* input  logic  [87:0] */ .classifier_map_extract_2_to_mem              (classifier_map_extract_2_to_mem),            
/* input  logic  [91:0] */ .classifier_map_port_cfg_to_mem               (classifier_map_port_cfg_to_mem),             
/* input  logic  [85:0] */ .classifier_map_port_default_0_to_mem         (classifier_map_port_default_0_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_10_to_mem        (classifier_map_port_default_10_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_11_to_mem        (classifier_map_port_default_11_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_12_to_mem        (classifier_map_port_default_12_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_13_to_mem        (classifier_map_port_default_13_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_14_to_mem        (classifier_map_port_default_14_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_15_to_mem        (classifier_map_port_default_15_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_16_to_mem        (classifier_map_port_default_16_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_17_to_mem        (classifier_map_port_default_17_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_18_to_mem        (classifier_map_port_default_18_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_19_to_mem        (classifier_map_port_default_19_to_mem),      
/* input  logic  [87:0] */ .classifier_map_ip_cfg_to_mem                 (classifier_map_ip_cfg_to_mem),               
/* input  logic  [87:0] */ .classifier_map_ip_hi_to_mem                  (classifier_map_ip_hi_to_mem),                
/* input  logic  [87:0] */ .classifier_map_ip_lo_to_mem                  (classifier_map_ip_lo_to_mem),                
/* input  logic  [91:0] */ .classifier_map_len_limit_to_mem              (classifier_map_len_limit_to_mem),            
/* input  logic  [85:0] */ .classifier_map_port_default_1_to_mem         (classifier_map_port_default_1_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_20_to_mem        (classifier_map_port_default_20_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_21_to_mem        (classifier_map_port_default_21_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_22_to_mem        (classifier_map_port_default_22_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_23_to_mem        (classifier_map_port_default_23_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_24_to_mem        (classifier_map_port_default_24_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_25_to_mem        (classifier_map_port_default_25_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_26_to_mem        (classifier_map_port_default_26_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_27_to_mem        (classifier_map_port_default_27_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_28_to_mem        (classifier_map_port_default_28_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_29_to_mem        (classifier_map_port_default_29_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_2_to_mem         (classifier_map_port_default_2_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_30_to_mem        (classifier_map_port_default_30_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_31_to_mem        (classifier_map_port_default_31_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_32_to_mem        (classifier_map_port_default_32_to_mem),      
/* input  logic  [85:0] */ .classifier_map_port_default_3_to_mem         (classifier_map_port_default_3_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_4_to_mem         (classifier_map_port_default_4_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_5_to_mem         (classifier_map_port_default_5_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_6_to_mem         (classifier_map_port_default_6_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_7_to_mem         (classifier_map_port_default_7_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_8_to_mem         (classifier_map_port_default_8_to_mem),       
/* input  logic  [85:0] */ .classifier_map_port_default_9_to_mem         (classifier_map_port_default_9_to_mem),       
/* input  logic  [91:0] */ .classifier_map_port_to_mem                   (classifier_map_port_to_mem),                 
/* input  logic  [85:0] */ .classifier_map_prot_to_mem                   (classifier_map_prot_to_mem),                 
/* input  logic  [89:0] */ .classifier_map_rewrite_0_to_mem              (classifier_map_rewrite_0_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_10_to_mem             (classifier_map_rewrite_10_to_mem),           
/* input  logic  [89:0] */ .classifier_map_rewrite_11_to_mem             (classifier_map_rewrite_11_to_mem),           
/* input  logic  [89:0] */ .classifier_map_rewrite_12_to_mem             (classifier_map_rewrite_12_to_mem),           
/* input  logic  [89:0] */ .classifier_map_rewrite_13_to_mem             (classifier_map_rewrite_13_to_mem),           
/* input  logic  [89:0] */ .classifier_map_rewrite_14_to_mem             (classifier_map_rewrite_14_to_mem),           
/* input  logic  [89:0] */ .classifier_map_rewrite_15_to_mem             (classifier_map_rewrite_15_to_mem),           
/* input  logic  [89:0] */ .classifier_map_rewrite_1_to_mem              (classifier_map_rewrite_1_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_2_to_mem              (classifier_map_rewrite_2_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_3_to_mem              (classifier_map_rewrite_3_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_4_to_mem              (classifier_map_rewrite_4_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_5_to_mem              (classifier_map_rewrite_5_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_6_to_mem              (classifier_map_rewrite_6_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_7_to_mem              (classifier_map_rewrite_7_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_8_to_mem              (classifier_map_rewrite_8_to_mem),            
/* input  logic  [89:0] */ .classifier_map_rewrite_9_to_mem              (classifier_map_rewrite_9_to_mem),            
/* input  logic  [87:0] */ .classifier_map_type_to_mem                   (classifier_map_type_to_mem),                 
/* input  logic  [89:0] */ .classifier_map_vpri_tc_to_mem                (classifier_map_vpri_tc_to_mem),              
/* input  logic  [89:0] */ .classifier_map_vpri_to_mem                   (classifier_map_vpri_to_mem),                 
/* input  logic  [85:0] */ .classifier_wcm_data_path_buffer0_to_mem      (classifier_wcm_data_path_buffer0_to_mem),    
/* output logic  [72:0] */ .classifier_map_len_limit_from_mem            (classifier_map_len_limit_from_mem),          
/* output logic  [72:0] */ .classifier_map_port_cfg_from_mem             (classifier_map_port_cfg_from_mem),           
/* output logic  [72:0] */ .classifier_map_port_default_0_from_mem       (classifier_map_port_default_0_from_mem),     
/* output logic  [60:0] */ .classifier_em_a_hash_cfg_from_mem            (classifier_em_a_hash_cfg_from_mem),          
/* output logic  [60:0] */ .classifier_em_b_hash_cfg_from_mem            (classifier_em_b_hash_cfg_from_mem),          
/* output logic  [72:0] */ .classifier_map_domain_pol_cfg_from_mem       (classifier_map_domain_pol_cfg_from_mem),     
/* output logic  [72:0] */ .classifier_map_exp_tc_from_mem               (classifier_map_exp_tc_from_mem),             
/* output logic  [72:0] */ .classifier_map_extract_0_from_mem            (classifier_map_extract_0_from_mem),          
/* output logic  [72:0] */ .classifier_map_extract_1_from_mem            (classifier_map_extract_1_from_mem),          
/* output logic  [72:0] */ .classifier_map_extract_2_from_mem            (classifier_map_extract_2_from_mem),          
/* output logic  [72:0] */ .classifier_map_ip_cfg_from_mem               (classifier_map_ip_cfg_from_mem),             
/* output logic  [72:0] */ .classifier_map_ip_hi_from_mem                (classifier_map_ip_hi_from_mem),              
/* output logic  [72:0] */ .classifier_map_ip_lo_from_mem                (classifier_map_ip_lo_from_mem),              
/* output logic  [72:0] */ .classifier_map_port_default_10_from_mem      (classifier_map_port_default_10_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_11_from_mem      (classifier_map_port_default_11_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_12_from_mem      (classifier_map_port_default_12_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_13_from_mem      (classifier_map_port_default_13_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_14_from_mem      (classifier_map_port_default_14_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_15_from_mem      (classifier_map_port_default_15_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_16_from_mem      (classifier_map_port_default_16_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_17_from_mem      (classifier_map_port_default_17_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_18_from_mem      (classifier_map_port_default_18_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_19_from_mem      (classifier_map_port_default_19_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_1_from_mem       (classifier_map_port_default_1_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_20_from_mem      (classifier_map_port_default_20_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_21_from_mem      (classifier_map_port_default_21_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_22_from_mem      (classifier_map_port_default_22_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_23_from_mem      (classifier_map_port_default_23_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_24_from_mem      (classifier_map_port_default_24_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_25_from_mem      (classifier_map_port_default_25_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_26_from_mem      (classifier_map_port_default_26_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_27_from_mem      (classifier_map_port_default_27_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_28_from_mem      (classifier_map_port_default_28_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_29_from_mem      (classifier_map_port_default_29_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_2_from_mem       (classifier_map_port_default_2_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_30_from_mem      (classifier_map_port_default_30_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_31_from_mem      (classifier_map_port_default_31_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_32_from_mem      (classifier_map_port_default_32_from_mem),    
/* output logic  [72:0] */ .classifier_map_port_default_3_from_mem       (classifier_map_port_default_3_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_4_from_mem       (classifier_map_port_default_4_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_5_from_mem       (classifier_map_port_default_5_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_6_from_mem       (classifier_map_port_default_6_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_7_from_mem       (classifier_map_port_default_7_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_8_from_mem       (classifier_map_port_default_8_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_default_9_from_mem       (classifier_map_port_default_9_from_mem),     
/* output logic  [72:0] */ .classifier_map_port_from_mem                 (classifier_map_port_from_mem),               
/* output logic  [72:0] */ .classifier_map_prot_from_mem                 (classifier_map_prot_from_mem),               
/* output logic  [72:0] */ .classifier_map_rewrite_0_from_mem            (classifier_map_rewrite_0_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_10_from_mem           (classifier_map_rewrite_10_from_mem),         
/* output logic  [72:0] */ .classifier_map_rewrite_11_from_mem           (classifier_map_rewrite_11_from_mem),         
/* output logic  [72:0] */ .classifier_map_rewrite_12_from_mem           (classifier_map_rewrite_12_from_mem),         
/* output logic  [72:0] */ .classifier_map_rewrite_13_from_mem           (classifier_map_rewrite_13_from_mem),         
/* output logic  [72:0] */ .classifier_map_rewrite_14_from_mem           (classifier_map_rewrite_14_from_mem),         
/* output logic  [72:0] */ .classifier_map_rewrite_15_from_mem           (classifier_map_rewrite_15_from_mem),         
/* output logic  [72:0] */ .classifier_map_rewrite_1_from_mem            (classifier_map_rewrite_1_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_2_from_mem            (classifier_map_rewrite_2_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_3_from_mem            (classifier_map_rewrite_3_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_4_from_mem            (classifier_map_rewrite_4_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_5_from_mem            (classifier_map_rewrite_5_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_6_from_mem            (classifier_map_rewrite_6_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_7_from_mem            (classifier_map_rewrite_7_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_8_from_mem            (classifier_map_rewrite_8_from_mem),          
/* output logic  [72:0] */ .classifier_map_rewrite_9_from_mem            (classifier_map_rewrite_9_from_mem),          
/* output logic  [72:0] */ .classifier_map_type_from_mem                 (classifier_map_type_from_mem),               
/* output logic  [72:0] */ .classifier_map_vpri_from_mem                 (classifier_map_vpri_from_mem),               
/* output logic  [72:0] */ .classifier_map_vpri_tc_from_mem              (classifier_map_vpri_tc_from_mem),            
/* output logic  [72:0] */ .classifier_wcm_data_path_buffer0_from_mem    (classifier_wcm_data_path_buffer0_from_mem));  
// End of module classifier_ff_mems from classifier_ff_mems


// module classifier_rf_mems    from classifier_rf_mems using classifier_rf_mems.map 
classifier_rf_mems    classifier_rf_mems(
/* input  logic          */ .car_raw_lan_power_good_with_byprst           (),                                           
/* input  logic          */ .cclk                                         (cclk),                                       
/* input  logic  [285:0] */ .classifier_em_a_delay_fifo_0_to_mem          (classifier_em_a_delay_fifo_0_to_mem),        
/* input  logic  [285:0] */ .classifier_em_a_delay_fifo_1_to_mem          (classifier_em_a_delay_fifo_1_to_mem),        
/* input  logic  [285:0] */ .classifier_em_a_delay_fifo_2_to_mem          (classifier_em_a_delay_fifo_2_to_mem),        
/* input  logic  [285:0] */ .classifier_em_a_delay_fifo_3_to_mem          (classifier_em_a_delay_fifo_3_to_mem),        
/* input  logic  [156:0] */ .classifier_em_a_hash_miss_to_mem             (classifier_em_a_hash_miss_to_mem),           
/* input  logic   [91:0] */ .classifier_em_a_key_mask_0_to_mem            (classifier_em_a_key_mask_0_to_mem),          
/* input  logic   [91:0] */ .classifier_em_a_key_mask_1_to_mem            (classifier_em_a_key_mask_1_to_mem),          
/* input  logic   [91:0] */ .classifier_em_a_key_mask_2_to_mem            (classifier_em_a_key_mask_2_to_mem),          
/* input  logic  [156:0] */ .classifier_em_b_hash_miss_to_mem             (classifier_em_b_hash_miss_to_mem),           
/* input  logic   [91:0] */ .classifier_em_b_key_mask_to_mem              (classifier_em_b_key_mask_to_mem),            
/* input  logic   [86:0] */ .classifier_map_l4_dst_to_mem                 (classifier_map_l4_dst_to_mem),               
/* input  logic   [86:0] */ .classifier_map_l4_src_to_mem                 (classifier_map_l4_src_to_mem),               
/* input  logic  [152:0] */ .classifier_map_mac_to_mem                    (classifier_map_mac_to_mem),                  
/* input  logic   [87:0] */ .classifier_map_profile_action_to_mem         (classifier_map_profile_action_to_mem),       
/* input  logic  [109:0] */ .classifier_map_profile_key0_to_mem           (classifier_map_profile_key0_to_mem),         
/* input  logic  [109:0] */ .classifier_map_profile_key1_to_mem           (classifier_map_profile_key1_to_mem),         
/* input  logic  [109:0] */ .classifier_map_profile_key_invert0_to_mem    (classifier_map_profile_key_invert0_to_mem),  
/* input  logic  [109:0] */ .classifier_map_profile_key_invert1_to_mem    (classifier_map_profile_key_invert1_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_0_to_mem    (classifier_wcm_data_path_buffer1_0_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_10_to_mem   (classifier_wcm_data_path_buffer1_10_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_11_to_mem   (classifier_wcm_data_path_buffer1_11_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_12_to_mem   (classifier_wcm_data_path_buffer1_12_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_13_to_mem   (classifier_wcm_data_path_buffer1_13_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_14_to_mem   (classifier_wcm_data_path_buffer1_14_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_15_to_mem   (classifier_wcm_data_path_buffer1_15_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_16_to_mem   (classifier_wcm_data_path_buffer1_16_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_17_to_mem   (classifier_wcm_data_path_buffer1_17_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_18_to_mem   (classifier_wcm_data_path_buffer1_18_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_19_to_mem   (classifier_wcm_data_path_buffer1_19_to_mem), 
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_1_to_mem    (classifier_wcm_data_path_buffer1_1_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_2_to_mem    (classifier_wcm_data_path_buffer1_2_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_3_to_mem    (classifier_wcm_data_path_buffer1_3_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_4_to_mem    (classifier_wcm_data_path_buffer1_4_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_5_to_mem    (classifier_wcm_data_path_buffer1_5_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_6_to_mem    (classifier_wcm_data_path_buffer1_6_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_7_to_mem    (classifier_wcm_data_path_buffer1_7_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_8_to_mem    (classifier_wcm_data_path_buffer1_8_to_mem),  
/* input  logic  [362:0] */ .classifier_wcm_data_path_buffer1_9_to_mem    (classifier_wcm_data_path_buffer1_9_to_mem),  
/* input  logic    [5:0] */ .fary_ffuse_data_misc_rf                      (),                                           
/* input  logic          */ .fary_pwren_b_rf                              (),                                           
/* input  logic          */ .fdfx_lbist_test_mode                         (),                                           
/* input  logic          */ .fscan_byprst_b                               (),                                           
/* input  logic   [37:0] */ .fscan_ram_awt_mode                           (),                                           
/* input  logic   [37:0] */ .fscan_ram_awt_ren                            (),                                           
/* input  logic   [37:0] */ .fscan_ram_awt_wen                            (),                                           
/* input  logic   [37:0] */ .fscan_ram_bypsel                             (),                                           
/* input  logic          */ .fscan_ram_init_en                            (),                                           
/* input  logic          */ .fscan_ram_init_val                           (),                                           
/* input  logic   [37:0] */ .fscan_ram_odis_b                             (),                                           
/* input  logic          */ .fscan_ram_rddis_b                            (),                                           
/* input  logic          */ .fscan_ram_wrdis_b                            (),                                           
/* input  logic          */ .fscan_rstbypen                               (),                                           
/* output logic   [88:0] */ .classifier_map_profile_key_invert0_from_mem  (classifier_map_profile_key_invert0_from_mem), 
/* output logic   [88:0] */ .classifier_map_profile_key_invert1_from_mem  (classifier_map_profile_key_invert1_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_0_from_mem  (classifier_wcm_data_path_buffer1_0_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_10_from_mem (classifier_wcm_data_path_buffer1_10_from_mem), 
/* output logic          */ .aary_pwren_b_rf                              (),                                           
/* output logic  [266:0] */ .classifier_em_a_delay_fifo_0_from_mem        (classifier_em_a_delay_fifo_0_from_mem),      
/* output logic  [266:0] */ .classifier_em_a_delay_fifo_1_from_mem        (classifier_em_a_delay_fifo_1_from_mem),      
/* output logic  [266:0] */ .classifier_em_a_delay_fifo_2_from_mem        (classifier_em_a_delay_fifo_2_from_mem),      
/* output logic  [266:0] */ .classifier_em_a_delay_fifo_3_from_mem        (classifier_em_a_delay_fifo_3_from_mem),      
/* output logic  [137:0] */ .classifier_em_a_hash_miss_from_mem           (classifier_em_a_hash_miss_from_mem),         
/* output logic   [72:0] */ .classifier_em_a_key_mask_0_from_mem          (classifier_em_a_key_mask_0_from_mem),        
/* output logic   [72:0] */ .classifier_em_a_key_mask_1_from_mem          (classifier_em_a_key_mask_1_from_mem),        
/* output logic   [72:0] */ .classifier_em_a_key_mask_2_from_mem          (classifier_em_a_key_mask_2_from_mem),        
/* output logic  [137:0] */ .classifier_em_b_hash_miss_from_mem           (classifier_em_b_hash_miss_from_mem),         
/* output logic   [72:0] */ .classifier_em_b_key_mask_from_mem            (classifier_em_b_key_mask_from_mem),          
/* output logic   [72:0] */ .classifier_map_l4_dst_from_mem               (classifier_map_l4_dst_from_mem),             
/* output logic   [72:0] */ .classifier_map_l4_src_from_mem               (classifier_map_l4_src_from_mem),             
/* output logic  [137:0] */ .classifier_map_mac_from_mem                  (classifier_map_mac_from_mem),                
/* output logic   [72:0] */ .classifier_map_profile_action_from_mem       (classifier_map_profile_action_from_mem),     
/* output logic   [88:0] */ .classifier_map_profile_key0_from_mem         (classifier_map_profile_key0_from_mem),       
/* output logic   [88:0] */ .classifier_map_profile_key1_from_mem         (classifier_map_profile_key1_from_mem),       
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_11_from_mem (classifier_wcm_data_path_buffer1_11_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_12_from_mem (classifier_wcm_data_path_buffer1_12_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_13_from_mem (classifier_wcm_data_path_buffer1_13_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_14_from_mem (classifier_wcm_data_path_buffer1_14_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_15_from_mem (classifier_wcm_data_path_buffer1_15_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_16_from_mem (classifier_wcm_data_path_buffer1_16_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_17_from_mem (classifier_wcm_data_path_buffer1_17_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_18_from_mem (classifier_wcm_data_path_buffer1_18_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_19_from_mem (classifier_wcm_data_path_buffer1_19_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_1_from_mem  (classifier_wcm_data_path_buffer1_1_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_2_from_mem  (classifier_wcm_data_path_buffer1_2_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_3_from_mem  (classifier_wcm_data_path_buffer1_3_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_4_from_mem  (classifier_wcm_data_path_buffer1_4_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_5_from_mem  (classifier_wcm_data_path_buffer1_5_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_6_from_mem  (classifier_wcm_data_path_buffer1_6_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_7_from_mem  (classifier_wcm_data_path_buffer1_7_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_8_from_mem  (classifier_wcm_data_path_buffer1_8_from_mem), 
/* output logic  [345:0] */ .classifier_wcm_data_path_buffer1_9_from_mem  (classifier_wcm_data_path_buffer1_9_from_mem)); 
// End of module classifier_rf_mems from classifier_rf_mems


// module classifier_sram_mems    from classifier_sram_mems using classifier_sram_mems.map 
classifier_sram_mems    classifier_sram_mems(
/* input  logic          */ .car_raw_lan_power_good_with_byprst           (),                                           
/* input  logic          */ .cclk                                         (cclk),                                       
/* input  logic  [104:0] */ .classifier_em_a_hash_lookup_to_mem           (classifier_em_a_hash_lookup_to_mem),         
/* input  logic  [101:0] */ .classifier_em_b_hash_lookup_to_mem           (classifier_em_b_hash_lookup_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_0_to_mem           (classifier_lpm_tree_state_0_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_10_to_mem          (classifier_lpm_tree_state_10_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_11_to_mem          (classifier_lpm_tree_state_11_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_12_to_mem          (classifier_lpm_tree_state_12_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_13_to_mem          (classifier_lpm_tree_state_13_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_14_to_mem          (classifier_lpm_tree_state_14_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_15_to_mem          (classifier_lpm_tree_state_15_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_16_to_mem          (classifier_lpm_tree_state_16_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_17_to_mem          (classifier_lpm_tree_state_17_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_78_to_mem          (classifier_lpm_tree_state_78_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_79_to_mem          (classifier_lpm_tree_state_79_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_7_to_mem           (classifier_lpm_tree_state_7_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_18_to_mem          (classifier_lpm_tree_state_18_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_19_to_mem          (classifier_lpm_tree_state_19_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_1_to_mem           (classifier_lpm_tree_state_1_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_20_to_mem          (classifier_lpm_tree_state_20_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_21_to_mem          (classifier_lpm_tree_state_21_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_22_to_mem          (classifier_lpm_tree_state_22_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_23_to_mem          (classifier_lpm_tree_state_23_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_24_to_mem          (classifier_lpm_tree_state_24_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_25_to_mem          (classifier_lpm_tree_state_25_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_26_to_mem          (classifier_lpm_tree_state_26_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_27_to_mem          (classifier_lpm_tree_state_27_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_28_to_mem          (classifier_lpm_tree_state_28_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_29_to_mem          (classifier_lpm_tree_state_29_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_2_to_mem           (classifier_lpm_tree_state_2_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_30_to_mem          (classifier_lpm_tree_state_30_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_31_to_mem          (classifier_lpm_tree_state_31_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_32_to_mem          (classifier_lpm_tree_state_32_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_33_to_mem          (classifier_lpm_tree_state_33_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_34_to_mem          (classifier_lpm_tree_state_34_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_35_to_mem          (classifier_lpm_tree_state_35_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_36_to_mem          (classifier_lpm_tree_state_36_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_37_to_mem          (classifier_lpm_tree_state_37_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_38_to_mem          (classifier_lpm_tree_state_38_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_39_to_mem          (classifier_lpm_tree_state_39_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_3_to_mem           (classifier_lpm_tree_state_3_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_40_to_mem          (classifier_lpm_tree_state_40_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_41_to_mem          (classifier_lpm_tree_state_41_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_42_to_mem          (classifier_lpm_tree_state_42_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_43_to_mem          (classifier_lpm_tree_state_43_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_44_to_mem          (classifier_lpm_tree_state_44_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_45_to_mem          (classifier_lpm_tree_state_45_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_46_to_mem          (classifier_lpm_tree_state_46_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_47_to_mem          (classifier_lpm_tree_state_47_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_48_to_mem          (classifier_lpm_tree_state_48_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_49_to_mem          (classifier_lpm_tree_state_49_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_4_to_mem           (classifier_lpm_tree_state_4_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_50_to_mem          (classifier_lpm_tree_state_50_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_51_to_mem          (classifier_lpm_tree_state_51_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_52_to_mem          (classifier_lpm_tree_state_52_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_53_to_mem          (classifier_lpm_tree_state_53_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_54_to_mem          (classifier_lpm_tree_state_54_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_55_to_mem          (classifier_lpm_tree_state_55_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_56_to_mem          (classifier_lpm_tree_state_56_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_57_to_mem          (classifier_lpm_tree_state_57_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_58_to_mem          (classifier_lpm_tree_state_58_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_59_to_mem          (classifier_lpm_tree_state_59_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_5_to_mem           (classifier_lpm_tree_state_5_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_60_to_mem          (classifier_lpm_tree_state_60_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_61_to_mem          (classifier_lpm_tree_state_61_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_62_to_mem          (classifier_lpm_tree_state_62_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_63_to_mem          (classifier_lpm_tree_state_63_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_64_to_mem          (classifier_lpm_tree_state_64_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_65_to_mem          (classifier_lpm_tree_state_65_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_66_to_mem          (classifier_lpm_tree_state_66_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_67_to_mem          (classifier_lpm_tree_state_67_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_68_to_mem          (classifier_lpm_tree_state_68_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_69_to_mem          (classifier_lpm_tree_state_69_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_6_to_mem           (classifier_lpm_tree_state_6_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_70_to_mem          (classifier_lpm_tree_state_70_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_71_to_mem          (classifier_lpm_tree_state_71_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_72_to_mem          (classifier_lpm_tree_state_72_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_73_to_mem          (classifier_lpm_tree_state_73_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_74_to_mem          (classifier_lpm_tree_state_74_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_75_to_mem          (classifier_lpm_tree_state_75_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_76_to_mem          (classifier_lpm_tree_state_76_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_77_to_mem          (classifier_lpm_tree_state_77_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_80_to_mem          (classifier_lpm_tree_state_80_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_81_to_mem          (classifier_lpm_tree_state_81_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_82_to_mem          (classifier_lpm_tree_state_82_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_83_to_mem          (classifier_lpm_tree_state_83_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_84_to_mem          (classifier_lpm_tree_state_84_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_85_to_mem          (classifier_lpm_tree_state_85_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_86_to_mem          (classifier_lpm_tree_state_86_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_87_to_mem          (classifier_lpm_tree_state_87_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_88_to_mem          (classifier_lpm_tree_state_88_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_89_to_mem          (classifier_lpm_tree_state_89_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_8_to_mem           (classifier_lpm_tree_state_8_to_mem),         
/* input  logic  [323:0] */ .classifier_lpm_tree_state_90_to_mem          (classifier_lpm_tree_state_90_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_91_to_mem          (classifier_lpm_tree_state_91_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_92_to_mem          (classifier_lpm_tree_state_92_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_93_to_mem          (classifier_lpm_tree_state_93_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_94_to_mem          (classifier_lpm_tree_state_94_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_95_to_mem          (classifier_lpm_tree_state_95_to_mem),        
/* input  logic  [323:0] */ .classifier_lpm_tree_state_9_to_mem           (classifier_lpm_tree_state_9_to_mem),         
/* input  logic   [92:0] */ .classifier_map_domain_action0_to_mem         (classifier_map_domain_action0_to_mem),       
/* input  logic   [92:0] */ .classifier_map_domain_action1_to_mem         (classifier_map_domain_action1_to_mem),       
/* input  logic   [89:0] */ .classifier_map_domain_profile_to_mem         (classifier_map_domain_profile_to_mem),       
/* input  logic   [91:0] */ .classifier_map_dscp_tc_to_mem                (classifier_map_dscp_tc_to_mem),              
/* input  logic   [88:0] */ .classifier_wcm_action_cfg_0_to_mem           (classifier_wcm_action_cfg_0_to_mem),         
/* input  logic   [88:0] */ .classifier_wcm_action_cfg_1_to_mem           (classifier_wcm_action_cfg_1_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_0_to_mem           (classifier_wcm_action_ram_0_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_10_to_mem          (classifier_wcm_action_ram_10_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_11_to_mem          (classifier_wcm_action_ram_11_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_12_to_mem          (classifier_wcm_action_ram_12_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_13_to_mem          (classifier_wcm_action_ram_13_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_14_to_mem          (classifier_wcm_action_ram_14_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_15_to_mem          (classifier_wcm_action_ram_15_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_16_to_mem          (classifier_wcm_action_ram_16_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_17_to_mem          (classifier_wcm_action_ram_17_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_18_to_mem          (classifier_wcm_action_ram_18_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_19_to_mem          (classifier_wcm_action_ram_19_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_1_to_mem           (classifier_wcm_action_ram_1_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_20_to_mem          (classifier_wcm_action_ram_20_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_21_to_mem          (classifier_wcm_action_ram_21_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_22_to_mem          (classifier_wcm_action_ram_22_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_23_to_mem          (classifier_wcm_action_ram_23_to_mem),        
/* input  logic   [90:0] */ .classifier_wcm_action_ram_2_to_mem           (classifier_wcm_action_ram_2_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_3_to_mem           (classifier_wcm_action_ram_3_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_4_to_mem           (classifier_wcm_action_ram_4_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_5_to_mem           (classifier_wcm_action_ram_5_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_6_to_mem           (classifier_wcm_action_ram_6_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_7_to_mem           (classifier_wcm_action_ram_7_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_8_to_mem           (classifier_wcm_action_ram_8_to_mem),         
/* input  logic   [90:0] */ .classifier_wcm_action_ram_9_to_mem           (classifier_wcm_action_ram_9_to_mem),         
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_0_to_mem         (classifier_wcm_tcam_cfg_ram_0_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_10_to_mem        (classifier_wcm_tcam_cfg_ram_10_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_11_to_mem        (classifier_wcm_tcam_cfg_ram_11_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_12_to_mem        (classifier_wcm_tcam_cfg_ram_12_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_13_to_mem        (classifier_wcm_tcam_cfg_ram_13_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_14_to_mem        (classifier_wcm_tcam_cfg_ram_14_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_15_to_mem        (classifier_wcm_tcam_cfg_ram_15_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_16_to_mem        (classifier_wcm_tcam_cfg_ram_16_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_17_to_mem        (classifier_wcm_tcam_cfg_ram_17_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_18_to_mem        (classifier_wcm_tcam_cfg_ram_18_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_19_to_mem        (classifier_wcm_tcam_cfg_ram_19_to_mem),      
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_1_to_mem         (classifier_wcm_tcam_cfg_ram_1_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_2_to_mem         (classifier_wcm_tcam_cfg_ram_2_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_3_to_mem         (classifier_wcm_tcam_cfg_ram_3_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_4_to_mem         (classifier_wcm_tcam_cfg_ram_4_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_5_to_mem         (classifier_wcm_tcam_cfg_ram_5_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_6_to_mem         (classifier_wcm_tcam_cfg_ram_6_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_7_to_mem         (classifier_wcm_tcam_cfg_ram_7_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_8_to_mem         (classifier_wcm_tcam_cfg_ram_8_to_mem),       
/* input  logic   [88:0] */ .classifier_wcm_tcam_cfg_ram_9_to_mem         (classifier_wcm_tcam_cfg_ram_9_to_mem),       
/* input  logic          */ .fary_enblfloat_sram                          (),                                           
/* input  logic          */ .fary_ensleep_sram                            (),                                           
/* input  logic   [19:0] */ .fary_ffuse_data_misc_sram                    (),                                           
/* input  logic    [1:0] */ .fary_fwen_sram                               (),                                           
/* input  logic          */ .fary_pwren_b_sram                            (),                                           
/* input  logic          */ .fary_stm_enable                              (),                                           
/* input  logic          */ .fary_stm_hilo                                (),                                           
/* input  logic          */ .fary_wakeup_sram                             (),                                           
/* input  logic          */ .fdfx_lbist_test_mode                         (),                                           
/* input  logic          */ .fscan_byprst_b                               (),                                           
/* input  logic          */ .fscan_mode                                   (),                                           
/* input  logic  [147:0] */ .fscan_ram_awt_mode                           (),                                           
/* input  logic  [147:0] */ .fscan_ram_awt_ren                            (),                                           
/* input  logic  [147:0] */ .fscan_ram_awt_wen                            (),                                           
/* input  logic  [147:0] */ .fscan_ram_bypsel                             (),                                           
/* input  logic          */ .fscan_ram_init_en                            (),                                           
/* input  logic          */ .fscan_ram_init_val                           (),                                           
/* input  logic  [147:0] */ .fscan_ram_odis_b                             (),                                           
/* input  logic          */ .fscan_ram_rddis_b                            (),                                           
/* input  logic          */ .fscan_ram_wrdis_b                            (),                                           
/* input  logic          */ .fscan_rstbypen                               (),                                           
/* output logic  [306:0] */ .classifier_lpm_tree_state_10_from_mem        (classifier_lpm_tree_state_10_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_11_from_mem        (classifier_lpm_tree_state_11_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_12_from_mem        (classifier_lpm_tree_state_12_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_13_from_mem        (classifier_lpm_tree_state_13_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_14_from_mem        (classifier_lpm_tree_state_14_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_15_from_mem        (classifier_lpm_tree_state_15_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_16_from_mem        (classifier_lpm_tree_state_16_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_17_from_mem        (classifier_lpm_tree_state_17_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_18_from_mem        (classifier_lpm_tree_state_18_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_19_from_mem        (classifier_lpm_tree_state_19_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_1_from_mem         (classifier_lpm_tree_state_1_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_20_from_mem        (classifier_lpm_tree_state_20_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_21_from_mem        (classifier_lpm_tree_state_21_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_22_from_mem        (classifier_lpm_tree_state_22_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_23_from_mem        (classifier_lpm_tree_state_23_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_28_from_mem        (classifier_lpm_tree_state_28_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_29_from_mem        (classifier_lpm_tree_state_29_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_2_from_mem         (classifier_lpm_tree_state_2_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_30_from_mem        (classifier_lpm_tree_state_30_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_31_from_mem        (classifier_lpm_tree_state_31_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_32_from_mem        (classifier_lpm_tree_state_32_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_33_from_mem        (classifier_lpm_tree_state_33_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_34_from_mem        (classifier_lpm_tree_state_34_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_35_from_mem        (classifier_lpm_tree_state_35_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_36_from_mem        (classifier_lpm_tree_state_36_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_37_from_mem        (classifier_lpm_tree_state_37_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_38_from_mem        (classifier_lpm_tree_state_38_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_39_from_mem        (classifier_lpm_tree_state_39_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_3_from_mem         (classifier_lpm_tree_state_3_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_40_from_mem        (classifier_lpm_tree_state_40_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_41_from_mem        (classifier_lpm_tree_state_41_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_42_from_mem        (classifier_lpm_tree_state_42_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_43_from_mem        (classifier_lpm_tree_state_43_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_44_from_mem        (classifier_lpm_tree_state_44_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_45_from_mem        (classifier_lpm_tree_state_45_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_46_from_mem        (classifier_lpm_tree_state_46_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_47_from_mem        (classifier_lpm_tree_state_47_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_48_from_mem        (classifier_lpm_tree_state_48_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_49_from_mem        (classifier_lpm_tree_state_49_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_4_from_mem         (classifier_lpm_tree_state_4_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_50_from_mem        (classifier_lpm_tree_state_50_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_51_from_mem        (classifier_lpm_tree_state_51_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_52_from_mem        (classifier_lpm_tree_state_52_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_53_from_mem        (classifier_lpm_tree_state_53_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_54_from_mem        (classifier_lpm_tree_state_54_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_55_from_mem        (classifier_lpm_tree_state_55_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_56_from_mem        (classifier_lpm_tree_state_56_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_57_from_mem        (classifier_lpm_tree_state_57_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_58_from_mem        (classifier_lpm_tree_state_58_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_59_from_mem        (classifier_lpm_tree_state_59_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_5_from_mem         (classifier_lpm_tree_state_5_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_60_from_mem        (classifier_lpm_tree_state_60_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_61_from_mem        (classifier_lpm_tree_state_61_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_62_from_mem        (classifier_lpm_tree_state_62_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_63_from_mem        (classifier_lpm_tree_state_63_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_64_from_mem        (classifier_lpm_tree_state_64_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_65_from_mem        (classifier_lpm_tree_state_65_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_66_from_mem        (classifier_lpm_tree_state_66_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_67_from_mem        (classifier_lpm_tree_state_67_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_68_from_mem        (classifier_lpm_tree_state_68_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_69_from_mem        (classifier_lpm_tree_state_69_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_6_from_mem         (classifier_lpm_tree_state_6_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_70_from_mem        (classifier_lpm_tree_state_70_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_71_from_mem        (classifier_lpm_tree_state_71_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_72_from_mem        (classifier_lpm_tree_state_72_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_73_from_mem        (classifier_lpm_tree_state_73_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_74_from_mem        (classifier_lpm_tree_state_74_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_75_from_mem        (classifier_lpm_tree_state_75_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_76_from_mem        (classifier_lpm_tree_state_76_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_77_from_mem        (classifier_lpm_tree_state_77_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_78_from_mem        (classifier_lpm_tree_state_78_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_79_from_mem        (classifier_lpm_tree_state_79_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_7_from_mem         (classifier_lpm_tree_state_7_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_80_from_mem        (classifier_lpm_tree_state_80_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_81_from_mem        (classifier_lpm_tree_state_81_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_82_from_mem        (classifier_lpm_tree_state_82_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_83_from_mem        (classifier_lpm_tree_state_83_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_84_from_mem        (classifier_lpm_tree_state_84_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_85_from_mem        (classifier_lpm_tree_state_85_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_86_from_mem        (classifier_lpm_tree_state_86_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_87_from_mem        (classifier_lpm_tree_state_87_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_88_from_mem        (classifier_lpm_tree_state_88_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_89_from_mem        (classifier_lpm_tree_state_89_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_8_from_mem         (classifier_lpm_tree_state_8_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_90_from_mem        (classifier_lpm_tree_state_90_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_91_from_mem        (classifier_lpm_tree_state_91_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_92_from_mem        (classifier_lpm_tree_state_92_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_93_from_mem        (classifier_lpm_tree_state_93_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_94_from_mem        (classifier_lpm_tree_state_94_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_95_from_mem        (classifier_lpm_tree_state_95_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_9_from_mem         (classifier_lpm_tree_state_9_from_mem),       
/* output logic   [72:0] */ .classifier_map_domain_action0_from_mem       (classifier_map_domain_action0_from_mem),     
/* output logic   [72:0] */ .classifier_map_domain_action1_from_mem       (classifier_map_domain_action1_from_mem),     
/* output logic   [72:0] */ .classifier_map_domain_profile_from_mem       (classifier_map_domain_profile_from_mem),     
/* output logic   [72:0] */ .classifier_map_dscp_tc_from_mem              (classifier_map_dscp_tc_from_mem),            
/* output logic   [68:0] */ .classifier_wcm_action_cfg_0_from_mem         (classifier_wcm_action_cfg_0_from_mem),       
/* output logic   [68:0] */ .classifier_wcm_action_cfg_1_from_mem         (classifier_wcm_action_cfg_1_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_0_from_mem         (classifier_wcm_action_ram_0_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_10_from_mem        (classifier_wcm_action_ram_10_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_11_from_mem        (classifier_wcm_action_ram_11_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_12_from_mem        (classifier_wcm_action_ram_12_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_13_from_mem        (classifier_wcm_action_ram_13_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_14_from_mem        (classifier_wcm_action_ram_14_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_15_from_mem        (classifier_wcm_action_ram_15_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_16_from_mem        (classifier_wcm_action_ram_16_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_17_from_mem        (classifier_wcm_action_ram_17_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_18_from_mem        (classifier_wcm_action_ram_18_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_19_from_mem        (classifier_wcm_action_ram_19_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_1_from_mem         (classifier_wcm_action_ram_1_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_20_from_mem        (classifier_wcm_action_ram_20_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_21_from_mem        (classifier_wcm_action_ram_21_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_22_from_mem        (classifier_wcm_action_ram_22_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_23_from_mem        (classifier_wcm_action_ram_23_from_mem),      
/* output logic   [72:0] */ .classifier_wcm_action_ram_2_from_mem         (classifier_wcm_action_ram_2_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_3_from_mem         (classifier_wcm_action_ram_3_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_4_from_mem         (classifier_wcm_action_ram_4_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_5_from_mem         (classifier_wcm_action_ram_5_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_6_from_mem         (classifier_wcm_action_ram_6_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_7_from_mem         (classifier_wcm_action_ram_7_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_8_from_mem         (classifier_wcm_action_ram_8_from_mem),       
/* output logic   [72:0] */ .classifier_wcm_action_ram_9_from_mem         (classifier_wcm_action_ram_9_from_mem),       
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_0_from_mem       (classifier_wcm_tcam_cfg_ram_0_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_10_from_mem      (classifier_wcm_tcam_cfg_ram_10_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_11_from_mem      (classifier_wcm_tcam_cfg_ram_11_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_12_from_mem      (classifier_wcm_tcam_cfg_ram_12_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_13_from_mem      (classifier_wcm_tcam_cfg_ram_13_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_14_from_mem      (classifier_wcm_tcam_cfg_ram_14_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_15_from_mem      (classifier_wcm_tcam_cfg_ram_15_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_16_from_mem      (classifier_wcm_tcam_cfg_ram_16_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_17_from_mem      (classifier_wcm_tcam_cfg_ram_17_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_18_from_mem      (classifier_wcm_tcam_cfg_ram_18_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_19_from_mem      (classifier_wcm_tcam_cfg_ram_19_from_mem),    
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_1_from_mem       (classifier_wcm_tcam_cfg_ram_1_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_2_from_mem       (classifier_wcm_tcam_cfg_ram_2_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_3_from_mem       (classifier_wcm_tcam_cfg_ram_3_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_4_from_mem       (classifier_wcm_tcam_cfg_ram_4_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_5_from_mem       (classifier_wcm_tcam_cfg_ram_5_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_6_from_mem       (classifier_wcm_tcam_cfg_ram_6_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_7_from_mem       (classifier_wcm_tcam_cfg_ram_7_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_8_from_mem       (classifier_wcm_tcam_cfg_ram_8_from_mem),     
/* output logic   [70:0] */ .classifier_wcm_tcam_cfg_ram_9_from_mem       (classifier_wcm_tcam_cfg_ram_9_from_mem),     
/* output logic  [306:0] */ .classifier_lpm_tree_state_24_from_mem        (classifier_lpm_tree_state_24_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_25_from_mem        (classifier_lpm_tree_state_25_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_26_from_mem        (classifier_lpm_tree_state_26_from_mem),      
/* output logic  [306:0] */ .classifier_lpm_tree_state_27_from_mem        (classifier_lpm_tree_state_27_from_mem),      
/* output logic          */ .aary_pwren_b_sram                            (),                                           
/* output logic   [80:0] */ .classifier_em_a_hash_lookup_from_mem         (classifier_em_a_hash_lookup_from_mem),       
/* output logic   [80:0] */ .classifier_em_b_hash_lookup_from_mem         (classifier_em_b_hash_lookup_from_mem),       
/* output logic  [306:0] */ .classifier_lpm_tree_state_0_from_mem         (classifier_lpm_tree_state_0_from_mem));       
// End of module classifier_sram_mems from classifier_sram_mems


// module classifier_tcam_mems    from classifier_tcam_mems using classifier_tcam_mems.map 
classifier_tcam_mems    classifier_tcam_mems(
/* input  logic           */ .cclk                                         (cclk),                                       
/* input  logic   [485:0] */ .classifier_lpm_key_cam_to_tcam               (classifier_lpm_key_cam_to_tcam),             
/* input  logic  [4434:0] */ .classifier_map_domain_tcam_to_tcam           (classifier_map_domain_tcam_to_tcam),         
/* input  logic  [1192:0] */ .classifier_wcm_tcam_0_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_10_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_11_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_12_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_13_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_14_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_15_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_16_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_17_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_18_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_19_to_tcam               (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_1_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_2_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_3_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_4_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_5_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_6_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_7_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_8_to_tcam                (),                                           
/* input  logic  [1192:0] */ .classifier_wcm_tcam_9_to_tcam                (),                                           
/* input  logic    [11:0] */ .fary_ffuse_tune_tcam                         (),                                           
/* input  logic           */ .fary_pwren_b_tcam                            (),                                           
/* input  logic           */ .fary_stm_enable                              (),                                           
/* input  logic           */ .fary_stm_hilo                                (),                                           
/* input  logic           */ .fdfx_lbist_test_mode                         (),                                           
/* input  logic           */ .fscan_clkungate                              (),                                           
/* input  logic           */ .fscan_mode                                   (),                                           
/* input  logic           */ .fscan_shiften                                (),                                           
/* output logic           */ .aary_pwren_b_tcam                            (),                                           
/* output logic   [326:0] */ .classifier_lpm_key_cam_from_tcam             (classifier_lpm_key_cam_from_tcam),           
/* output logic  [4181:0] */ .classifier_map_domain_tcam_from_tcam         (classifier_map_domain_tcam_from_tcam),       
/* output logic  [1069:0] */ .classifier_wcm_tcam_0_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_10_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_11_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_12_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_13_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_14_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_15_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_16_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_17_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_18_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_19_from_tcam             (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_1_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_2_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_3_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_4_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_5_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_6_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_7_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_8_from_tcam              (),                                           
/* output logic  [1069:0] */ .classifier_wcm_tcam_9_from_tcam              ());                                           
// End of module classifier_tcam_mems from classifier_tcam_mems

endmodule // classifier_top
