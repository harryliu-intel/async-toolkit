magic
tech scmos
timestamp 965070614
<< ndiffusion >>
rect -9 85 -1 86
rect -9 77 -1 82
rect -9 69 -1 74
rect -9 61 -1 66
rect -9 53 -1 58
rect -9 45 -1 50
rect -9 41 -1 42
<< pdiffusion >>
rect 22 100 30 101
rect 22 96 30 97
rect 22 87 30 88
rect 22 83 30 84
rect 22 74 30 75
rect 22 70 30 71
rect 22 61 30 62
rect 22 57 30 58
rect 22 48 30 49
rect 22 44 30 45
rect 22 35 30 36
rect 22 31 30 32
<< ntransistor >>
rect -9 82 -1 85
rect -9 74 -1 77
rect -9 66 -1 69
rect -9 58 -1 61
rect -9 50 -1 53
rect -9 42 -1 45
<< ptransistor >>
rect 22 97 30 100
rect 22 84 30 87
rect 22 71 30 74
rect 22 58 30 61
rect 22 45 30 48
rect 22 32 30 35
<< polysilicon >>
rect 1 97 22 100
rect 30 97 34 100
rect 1 85 4 97
rect -13 82 -9 85
rect -1 82 4 85
rect 9 84 22 87
rect 30 84 34 87
rect 9 77 12 84
rect -13 74 -9 77
rect -1 74 12 77
rect 17 71 22 74
rect 30 71 34 74
rect 17 69 20 71
rect -13 66 -9 69
rect -1 66 20 69
rect -13 58 -9 61
rect -1 58 22 61
rect 30 58 34 61
rect -13 50 -9 53
rect -1 50 20 53
rect 17 48 20 50
rect 17 45 22 48
rect 30 45 34 48
rect -13 42 -9 45
rect -1 42 11 45
rect 8 35 11 42
rect 8 32 22 35
rect 30 32 34 35
<< ndcontact >>
rect -9 86 -1 94
rect -9 33 -1 41
<< pdcontact >>
rect 22 101 30 109
rect 22 88 30 96
rect 22 75 30 83
rect 22 62 30 70
rect 22 49 30 57
rect 22 36 30 44
rect 22 23 30 31
<< metal1 >>
rect 22 101 30 109
rect 11 94 30 96
rect -9 88 30 94
rect -9 86 18 88
rect 10 70 18 86
rect 22 75 30 83
rect 10 62 30 70
rect 10 44 18 62
rect 22 49 30 57
rect -9 33 -1 41
rect 10 36 30 44
rect 22 23 30 31
<< labels >>
rlabel metal1 26 40 26 40 1 x
rlabel metal1 26 53 26 53 5 Vdd!
rlabel metal1 26 27 26 27 1 Vdd!
rlabel polysilicon 31 46 31 46 1 b
rlabel polysilicon 31 33 31 33 1 a
rlabel metal1 26 66 26 66 5 x
rlabel polysilicon 31 59 31 59 1 c
rlabel metal1 26 79 26 79 1 Vdd!
rlabel polysilicon 31 72 31 72 1 d
rlabel metal1 26 92 26 92 1 x
rlabel polysilicon 31 85 31 85 1 e
rlabel metal1 26 105 26 105 5 Vdd!
rlabel metal1 -5 37 -5 37 1 GND!
rlabel polysilicon -10 43 -10 43 3 a
rlabel polysilicon -10 51 -10 51 3 b
rlabel polysilicon -10 59 -10 59 3 c
rlabel polysilicon -10 67 -10 67 3 d
rlabel polysilicon -10 75 -10 75 3 e
rlabel metal1 -5 90 -5 90 1 x
rlabel polysilicon -10 83 -10 83 3 f
rlabel polysilicon 31 98 31 98 1 f
rlabel space -14 33 -9 94 7 ^n
rlabel space 30 23 35 109 3 ^p
<< end >>
