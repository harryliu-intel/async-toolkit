//                                                                             
// File:       TLM1_classes.svh                                                 
// Creator:    kmoses1                                                         
// Time:       Thursday Jan 16, 2014 [3:40:08 pm]                              
//                                                                             
// Path:       /tmp/kmoses1/nebulon_run/1248                                   
// Arguments:  /p/com/eda/denali/blueprint/3.7.4/Linux/blueprint -cspec -fuse  
//             -html -I /p/com/eda/intel/nebulon/2.07p1/include/               
//             fusegen-Nebulon.rdl                                             
//                                                                             
// Sources:    /nfs/iil/proj/mpg/kmoses1_wa/SOCFuseGen/TLM1/fusegen-Nebulon.rdl:5b3e806ef7d09a39437507f3cfbd0ecb
//             /p/com/eda/intel/nebulon/2.07p1/generators/fuse.pm              
//             /p/com/eda/intel/nebulon/2.07p1/generators/generator_common.pm  
//             /p/com/eda/intel/nebulon/2.07p1/generators/html.pm              
//             /p/com/eda/intel/nebulon/2.07p1/include/fuse_udp.rdl:c11891ce81c95bc748bf1f2bdbde2f6f
//             /usr/intel/pkgs/perl/5.8.7/lib64/5.8.7/Digest/base.pm           
//             /usr/intel/pkgs/perl/5.8.7/lib64/site_perl/Devel/StackTrace.pm  
//                                                                             
// Blueprint:   3.7.4 (Tue Jun 23 00:17:01 PDT 2009)                           
// Machine:    ivnc0059                                                        
// OS:         Linux 2.6.16.60-0.58.1.3835.0.PTF.638363-smp                    
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2014 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY DENALI BLUEPRINT, DO NOT EDIT       
//                                                                             


//Fuse code compatible with Saola versions: v20131113 and newer 

class tlm_fuse_tlm_fuse_fuse_1_field extends slu_fuse;

    rand bit [   7:   0] cfg_val;
    logic [   7:   0] desired_val;
    bit [   7:   0] configuration_values[int unsigned];
    bit [   7:   0] configuration_value;

   `uvm_object_utils(tlm_fuse_tlm_fuse_fuse_1_field)

   function void do_print (uvm_printer printer);
      super.do_print(printer);
      printer.print_field("cfg_val", cfg_val, $bits(cfg_val));
      printer.print_field("desired_val", desired_val, $bits(desired_val));
   endfunction

   function void do_pack (uvm_packer packer);
      super.do_pack(packer);
      packer.pack_field_int(cfg_val, $bits(cfg_val));
   endfunction

    constraint default_c {cfg_val == 8'hCA;};
    constraint configuration_c { cfg_val == configuration_value; };

    function new (string name = "tlm_fuse_tlm_fuse_fuse_1_field");
        super.new(name);
        set_default();
    endfunction

    function void set_default();
        super.set_size(8);
        desired_val = 8'hCA;
        super.set_pull_once(0); 
        super.set_blk_on_dbg(0); 
        super.set_ram_address(17'h00008);
        super.set_start_bit(4'h0); 
        set_configuration_constraint(0);
        super.set_rcvraddr(8'b0);
        super.set_request_type("Group0");
        super.set_jtagrd(0);
        super.set_jtagwr(0);
        super.set_csrrd(0);
        super.set_csrwr(0);
        super.set_group_type("DF");
        super.set_rd4err(0);
        super.set_array_type("HS");
        set_lockout_valid_tag("1"); 
        set_category("IntelHVM"); 
        super.set_lldd(0);
    endfunction

    function void set_rand_mode (int mode);
        if (mode==1) cfg_val.rand_mode(1);
        else cfg_val.rand_mode(0);
    endfunction

   function void set_cfg_val (logic val[]);
      for(int i=0; i< val.size(); i++)
         this.cfg_val[i] = val[i];
   endfunction

    function void get_desired_val(ref logic val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.desired_val[i];
    endfunction

    function void get_cfg_val(ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.cfg_val[i];
    endfunction

    function void set_desired_val(logic val[]);
        for(int i=0; i< val.size(); i++)
           this.desired_val[i] = val[i];
    endfunction

    function void set_configuration_constraint(bit enable, int mode=0);
       if (!enable) configuration_c.constraint_mode(0);
       else if (has_configuration_value(mode)) begin
         bit val[];
         get_configuration_value(mode, val);
         configuration_value = {<<{val}};
         set_default_constraint(0); 
         configuration_c.constraint_mode(1);
       end //if has_configuration_value
    endfunction : set_configuration_constraint


    function void set_configuration_value(int unsigned mode, bit val[]);
        for(int i=0; i< get_size(); i++)
           this.configuration_values[mode][i] = val[i];
    endfunction


    function void get_configuration_value(int unsigned mode, ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.configuration_values[mode][i];
    endfunction


    function bit has_configuration_value(int unsigned mode);
       return(configuration_values.exists(mode));
    endfunction

    function void mirror_desired(); 
    desired_val = cfg_val;
    endfunction

    function void reset_desired();
    desired_val = 8'b0;
    endfunction

endclass

class tlm_fuse_tlm_fuse_fuse_2_field extends slu_fuse;

    rand bit [   5:   0] cfg_val;
    logic [   5:   0] desired_val;
    bit [   5:   0] configuration_values[int unsigned];
    bit [   5:   0] configuration_value;

   `uvm_object_utils(tlm_fuse_tlm_fuse_fuse_2_field)

   function void do_print (uvm_printer printer);
      super.do_print(printer);
      printer.print_field("cfg_val", cfg_val, $bits(cfg_val));
      printer.print_field("desired_val", desired_val, $bits(desired_val));
   endfunction

   function void do_pack (uvm_packer packer);
      super.do_pack(packer);
      packer.pack_field_int(cfg_val, $bits(cfg_val));
   endfunction

    constraint default_c {cfg_val == 6'b100100;};
    constraint configuration_c { cfg_val == configuration_value; };

    function new (string name = "tlm_fuse_tlm_fuse_fuse_2_field");
        super.new(name);
        set_default();
    endfunction

    function void set_default();
        super.set_size(6);
        desired_val = 6'b100100;
        super.set_pull_once(0); 
        super.set_blk_on_dbg(0); 
        super.set_ram_address(17'h00400);
        super.set_start_bit(4'h0); 
        set_configuration_constraint(0);
        super.set_rcvraddr('d1);
        super.set_request_type("Group0");
        super.set_jtagrd(0);
        super.set_jtagwr(0);
        super.set_csrrd(0);
        super.set_csrwr(0);
        super.set_group_type("DF");
        super.set_rd4err(0);
        super.set_array_type("HD");
        set_lockout_valid_tag("2"); 
        set_category("IntelHVM"); 
        super.set_lldd(0);
    endfunction

    function void set_rand_mode (int mode);
        if (mode==1) cfg_val.rand_mode(1);
        else cfg_val.rand_mode(0);
    endfunction

   function void set_cfg_val (logic val[]);
      for(int i=0; i< val.size(); i++)
         this.cfg_val[i] = val[i];
   endfunction

    function void get_desired_val(ref logic val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.desired_val[i];
    endfunction

    function void get_cfg_val(ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.cfg_val[i];
    endfunction

    function void set_desired_val(logic val[]);
        for(int i=0; i< val.size(); i++)
           this.desired_val[i] = val[i];
    endfunction

    function void set_configuration_constraint(bit enable, int mode=0);
       if (!enable) configuration_c.constraint_mode(0);
       else if (has_configuration_value(mode)) begin
         bit val[];
         get_configuration_value(mode, val);
         configuration_value = {<<{val}};
         set_default_constraint(0); 
         configuration_c.constraint_mode(1);
       end //if has_configuration_value
    endfunction : set_configuration_constraint


    function void set_configuration_value(int unsigned mode, bit val[]);
        for(int i=0; i< get_size(); i++)
           this.configuration_values[mode][i] = val[i];
    endfunction


    function void get_configuration_value(int unsigned mode, ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.configuration_values[mode][i];
    endfunction


    function bit has_configuration_value(int unsigned mode);
       return(configuration_values.exists(mode));
    endfunction

    function void mirror_desired(); 
    desired_val = cfg_val;
    endfunction

    function void reset_desired();
    desired_val = 6'b0;
    endfunction

endclass

class tlm_fuse_tlm_fuse_fuse_3_field extends slu_fuse;

    rand bit [   1:   0] cfg_val;
    logic [   1:   0] desired_val;
    bit [   1:   0] configuration_values[int unsigned];
    bit [   1:   0] configuration_value;

   `uvm_object_utils(tlm_fuse_tlm_fuse_fuse_3_field)

   function void do_print (uvm_printer printer);
      super.do_print(printer);
      printer.print_field("cfg_val", cfg_val, $bits(cfg_val));
      printer.print_field("desired_val", desired_val, $bits(desired_val));
   endfunction

   function void do_pack (uvm_packer packer);
      super.do_pack(packer);
      packer.pack_field_int(cfg_val, $bits(cfg_val));
   endfunction

    constraint default_c {cfg_val == 2'b11;};
    constraint configuration_c { cfg_val == configuration_value; };

    function new (string name = "tlm_fuse_tlm_fuse_fuse_3_field");
        super.new(name);
        set_default();
    endfunction

    function void set_default();
        super.set_size(2);
        desired_val = 2'b11;
        super.set_pull_once(0); 
        super.set_blk_on_dbg(0); 
        super.set_ram_address(17'h00400);
        super.set_start_bit('d6); 
        set_configuration_constraint(0);
        super.set_rcvraddr('d1);
        super.set_request_type("Group0");
        super.set_jtagrd(0);
        super.set_jtagwr(0);
        super.set_csrrd(0);
        super.set_csrwr(0);
        super.set_group_type("DF");
        super.set_rd4err(0);
        super.set_array_type("HD");
        set_lockout_valid_tag("2"); 
        set_category("IntelHVM"); 
        super.set_lldd(0);
    endfunction

    function void set_rand_mode (int mode);
        if (mode==1) cfg_val.rand_mode(1);
        else cfg_val.rand_mode(0);
    endfunction

   function void set_cfg_val (logic val[]);
      for(int i=0; i< val.size(); i++)
         this.cfg_val[i] = val[i];
   endfunction

    function void get_desired_val(ref logic val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.desired_val[i];
    endfunction

    function void get_cfg_val(ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.cfg_val[i];
    endfunction

    function void set_desired_val(logic val[]);
        for(int i=0; i< val.size(); i++)
           this.desired_val[i] = val[i];
    endfunction

    function void set_configuration_constraint(bit enable, int mode=0);
       if (!enable) configuration_c.constraint_mode(0);
       else if (has_configuration_value(mode)) begin
         bit val[];
         get_configuration_value(mode, val);
         configuration_value = {<<{val}};
         set_default_constraint(0); 
         configuration_c.constraint_mode(1);
       end //if has_configuration_value
    endfunction : set_configuration_constraint


    function void set_configuration_value(int unsigned mode, bit val[]);
        for(int i=0; i< get_size(); i++)
           this.configuration_values[mode][i] = val[i];
    endfunction


    function void get_configuration_value(int unsigned mode, ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.configuration_values[mode][i];
    endfunction


    function bit has_configuration_value(int unsigned mode);
       return(configuration_values.exists(mode));
    endfunction

    function void mirror_desired(); 
    desired_val = cfg_val;
    endfunction

    function void reset_desired();
    desired_val = 2'b0;
    endfunction

endclass

class tlm_fuse_tlm_fuse_fuse_4_field extends slu_fuse;

    rand bit [   7:   0] cfg_val;
    logic [   7:   0] desired_val;
    bit [   7:   0] configuration_values[int unsigned];
    bit [   7:   0] configuration_value;

   `uvm_object_utils(tlm_fuse_tlm_fuse_fuse_4_field)

   function void do_print (uvm_printer printer);
      super.do_print(printer);
      printer.print_field("cfg_val", cfg_val, $bits(cfg_val));
      printer.print_field("desired_val", desired_val, $bits(desired_val));
   endfunction

   function void do_pack (uvm_packer packer);
      super.do_pack(packer);
      packer.pack_field_int(cfg_val, $bits(cfg_val));
   endfunction

    constraint default_c {cfg_val == 8'hAD;};
    constraint configuration_c { cfg_val == configuration_value; };

    function new (string name = "tlm_fuse_tlm_fuse_fuse_4_field");
        super.new(name);
        set_default();
    endfunction

    function void set_default();
        super.set_size(8);
        desired_val = 8'hAD;
        super.set_pull_once(0); 
        super.set_blk_on_dbg(0); 
        super.set_ram_address(17'h00404);
        super.set_start_bit(4'h0); 
        set_configuration_constraint(0);
        super.set_rcvraddr('d2);
        super.set_request_type("Group1");
        super.set_jtagrd(0);
        super.set_jtagwr(0);
        super.set_csrrd(0);
        super.set_csrwr(0);
        super.set_group_type("DF");
        super.set_rd4err(0);
        super.set_array_type("HD");
        set_lockout_valid_tag("3"); 
        set_category("IntelHVM"); 
        super.set_lldd(0);
    endfunction

    function void set_rand_mode (int mode);
        if (mode==1) cfg_val.rand_mode(1);
        else cfg_val.rand_mode(0);
    endfunction

   function void set_cfg_val (logic val[]);
      for(int i=0; i< val.size(); i++)
         this.cfg_val[i] = val[i];
   endfunction

    function void get_desired_val(ref logic val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.desired_val[i];
    endfunction

    function void get_cfg_val(ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.cfg_val[i];
    endfunction

    function void set_desired_val(logic val[]);
        for(int i=0; i< val.size(); i++)
           this.desired_val[i] = val[i];
    endfunction

    function void set_configuration_constraint(bit enable, int mode=0);
       if (!enable) configuration_c.constraint_mode(0);
       else if (has_configuration_value(mode)) begin
         bit val[];
         get_configuration_value(mode, val);
         configuration_value = {<<{val}};
         set_default_constraint(0); 
         configuration_c.constraint_mode(1);
       end //if has_configuration_value
    endfunction : set_configuration_constraint


    function void set_configuration_value(int unsigned mode, bit val[]);
        for(int i=0; i< get_size(); i++)
           this.configuration_values[mode][i] = val[i];
    endfunction


    function void get_configuration_value(int unsigned mode, ref bit val[]);
        val = new[get_size()];
        for(int i=0; i<get_size(); i++)
           val[i] = this.configuration_values[mode][i];
    endfunction


    function bit has_configuration_value(int unsigned mode);
       return(configuration_values.exists(mode));
    endfunction

    function void mirror_desired(); 
    desired_val = cfg_val;
    endfunction

    function void reset_desired();
    desired_val = 8'b0;
    endfunction

endclass

class tlm_fuse_fusegroup extends slu_fuse_group;
    rand tlm_fuse_tlm_fuse_fuse_1_field tlm_fuse_tlm_fuse_fuse_1;
    rand tlm_fuse_tlm_fuse_fuse_2_field tlm_fuse_tlm_fuse_fuse_2;
    rand tlm_fuse_tlm_fuse_fuse_3_field tlm_fuse_tlm_fuse_fuse_3;
    rand tlm_fuse_tlm_fuse_fuse_4_field tlm_fuse_tlm_fuse_fuse_4;

    `uvm_object_utils(tlm_fuse_fusegroup)

    function void do_print (uvm_printer printer);
       super.do_print(printer);
        printer.print_object("tlm_fuse_tlm_fuse_fuse_1", tlm_fuse_tlm_fuse_fuse_1);
        printer.print_object("tlm_fuse_tlm_fuse_fuse_2", tlm_fuse_tlm_fuse_fuse_2);
        printer.print_object("tlm_fuse_tlm_fuse_fuse_3", tlm_fuse_tlm_fuse_fuse_3);
        printer.print_object("tlm_fuse_tlm_fuse_fuse_4", tlm_fuse_tlm_fuse_fuse_4);
    endfunction

    function void do_pack (uvm_packer packer);
       super.do_pack(packer);
       packer.pack_object(tlm_fuse_tlm_fuse_fuse_1);
       packer.pack_object(tlm_fuse_tlm_fuse_fuse_2);
       packer.pack_object(tlm_fuse_tlm_fuse_fuse_3);
       packer.pack_object(tlm_fuse_tlm_fuse_fuse_4);
    endfunction

    function new (string name = "tlm_fuse_fusegroup");
        super.new(name);
        set_default();
        this.build_phase();
    endfunction

    function void build_phase(uvm_phase phase = null);
        tlm_fuse_tlm_fuse_fuse_1 = tlm_fuse_tlm_fuse_fuse_1_field::type_id::create("tlm_fuse_tlm_fuse_fuse_1");
        tlm_fuse_tlm_fuse_fuse_1.set_group(this);
        tlm_fuse_tlm_fuse_fuse_2 = tlm_fuse_tlm_fuse_fuse_2_field::type_id::create("tlm_fuse_tlm_fuse_fuse_2");
        tlm_fuse_tlm_fuse_fuse_2.set_group(this);
        tlm_fuse_tlm_fuse_fuse_3 = tlm_fuse_tlm_fuse_fuse_3_field::type_id::create("tlm_fuse_tlm_fuse_fuse_3");
        tlm_fuse_tlm_fuse_fuse_3.set_group(this);
        tlm_fuse_tlm_fuse_fuse_4 = tlm_fuse_tlm_fuse_fuse_4_field::type_id::create("tlm_fuse_tlm_fuse_fuse_4");
        tlm_fuse_tlm_fuse_fuse_4.set_group(this);

    endfunction

    function add_fuses();
        _env.add_fuse("tlm_fuse_tlm_fuse_fuse_1", tlm_fuse_tlm_fuse_fuse_1);
        _env.add_fuse("tlm_fuse_tlm_fuse_fuse_2", tlm_fuse_tlm_fuse_fuse_2);
        _env.add_fuse("tlm_fuse_tlm_fuse_fuse_3", tlm_fuse_tlm_fuse_fuse_3);
        _env.add_fuse("tlm_fuse_tlm_fuse_fuse_4", tlm_fuse_tlm_fuse_fuse_4);
    endfunction

    function void set_default();
        super.set_size(24);
        super.set_cmplfmt('d1);
        super.set_sai(16'b0);
    endfunction

    function void pre_randomize();
        super.pre_randomize();
        if ($value$plusargs("tlm_fuse_tlm_fuse_fuse_1=%b",tlm_fuse_tlm_fuse_fuse_1.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_1.rand_mode(0);
        end
        else if(_env.get_config_int("tlm_fuse_tlm_fuse_fuse_1", tlm_fuse_tlm_fuse_fuse_1.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_1.rand_mode(0);
        end
        if ($value$plusargs("tlm_fuse_tlm_fuse_fuse_2=%b",tlm_fuse_tlm_fuse_fuse_2.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_2.rand_mode(0);
        end
        else if(_env.get_config_int("tlm_fuse_tlm_fuse_fuse_2", tlm_fuse_tlm_fuse_fuse_2.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_2.rand_mode(0);
        end
        if ($value$plusargs("tlm_fuse_tlm_fuse_fuse_3=%b",tlm_fuse_tlm_fuse_fuse_3.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_3.rand_mode(0);
        end
        else if(_env.get_config_int("tlm_fuse_tlm_fuse_fuse_3", tlm_fuse_tlm_fuse_fuse_3.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_3.rand_mode(0);
        end
        if ($value$plusargs("tlm_fuse_tlm_fuse_fuse_4=%b",tlm_fuse_tlm_fuse_fuse_4.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_4.rand_mode(0);
        end
        else if(_env.get_config_int("tlm_fuse_tlm_fuse_fuse_4", tlm_fuse_tlm_fuse_fuse_4.cfg_val)) begin
            tlm_fuse_tlm_fuse_fuse_4.rand_mode(0);
        end
    endfunction
     virtual function void print_sv_fusegroup_file();  
       $display("FuseGroup Type [%s], FuseGroup Instance [%s], SV File ---> %s", get_type_name(), get_name(), `__FILE__); 
    endfunction 

endclass : tlm_fuse_fusegroup

