///------------------------------------------------------------------------------
///                                                                              
///  INTEL CONFIDENTIAL                                                          
///                                                                              
///  Copyright 2018 Intel Corporation All Rights Reserved.                 
///                                                                              
///  The source code contained or described herein and all documents related     
///  to the source code ("Material") are owned by Intel Corporation or its    
///  suppliers or licensors. Title to the Material remains with Intel            
///  Corporation or its suppliers and licensors. The Material contains trade     
///  secrets and proprietary and confidential information of Intel or its        
///  suppliers and licensors. The Material is protected by worldwide copyright   
///  and trade secret laws and treaty provisions. No part of the Material may    
///  be used, copied, reproduced, modified, published, uploaded, posted,         
///  transmitted, distributed, or disclosed in any way without Intel's prior     
///  express written permission.                                                 
///                                                                              
///  No license under any patent, copyright, trade secret or other intellectual  
///  property right is granted to or conferred upon you by disclosure or         
///  delivery of the Materials, either expressly, by implication, inducement,    
///  estoppel or otherwise. Any license under such intellectual property rights  
///  must be express and approved by Intel in writing.                           
///                                                                              
///------------------------------------------------------------------------------
///  Auto-generated by ngen. please do not hand edit
///------------------------------------------------------------------------------
// -- Author       : Mike Jarvis <michael.a.jarvis.com> 
// -- Project Name : MBY 
// -- Description  : mgp (MeGaPort) netlist. 
// ------------------------------------------------------------------- 

module mgp (
//Input List
input                   arst_n,                                   //Asynchronous negedge reset    
input                   cclk,                                     
input                   clk,                                      
input            [7:0]  epl0_igr_rx_data_valid,                   
input         [0:7][71:0]  epl0_igr_rx_data_w_ecc,                   
input            [7:0]  epl0_igr_rx_ecc,                          
input            [2:0]  epl0_igr_rx_flow_control_tc,              
input           [23:0]  epl0_igr_rx_metadata,                     
input                   epl0_igr_rx_pfc_xoff,                     
input            [1:0]  epl0_igr_rx_port_num,                     
input           [35:0]  epl0_igr_rx_time_stamp,                   
input            [7:0]  epl1_igr_rx_data_valid,                   
input         [0:7][71:0]  epl1_igr_rx_data_w_ecc,                   
input            [7:0]  epl1_igr_rx_ecc,                          
input            [2:0]  epl1_igr_rx_flow_control_tc,              
input           [23:0]  epl1_igr_rx_metadata,                     
input                   epl1_igr_rx_pfc_xoff,                     
input            [1:0]  epl1_igr_rx_port_num,                     
input           [35:0]  epl1_igr_rx_time_stamp,                   
input            [7:0]  epl2_igr_rx_data_valid,                   
input         [0:7][71:0]  epl2_igr_rx_data_w_ecc,                   
input            [7:0]  epl2_igr_rx_ecc,                          
input            [2:0]  epl2_igr_rx_flow_control_tc,              
input           [23:0]  epl2_igr_rx_metadata,                     
input                   epl2_igr_rx_pfc_xoff,                     
input            [1:0]  epl2_igr_rx_port_num,                     
input           [35:0]  epl2_igr_rx_time_stamp,                   
input            [7:0]  epl3_igr_rx_data_valid,                   
input         [0:7][71:0]  epl3_igr_rx_data_w_ecc,                   
input            [7:0]  epl3_igr_rx_ecc,                          
input            [2:0]  epl3_igr_rx_flow_control_tc,              
input           [23:0]  epl3_igr_rx_metadata,                     
input                   epl3_igr_rx_pfc_xoff,                     
input            [1:0]  epl3_igr_rx_port_num,                     
input           [35:0]  epl3_igr_rx_time_stamp,                   
input           [19:0]  igr_vp_cpp_rx_metadata,                   
input            [7:0]  igr_vp_rx_data_valid,                     
input         [0:7][71:0]  igr_vp_rx_data_w_ecc,                     
input            [7:0]  igr_vp_rx_ecc,                            
input            [2:0]  igr_vp_rx_flow_control_tc,                
input           [23:0]  igr_vp_rx_metadata,                       
input            [1:0]  igr_vp_rx_port_num,                       
input           [35:0]  igr_vp_rx_time_stamp,                     
input                   reset,                                    
input                   rst_n,                                    //taken from HLP active low for MBY? 

//Interface List
ahb_rx_ppe_if.ppe                 ahb_rx_ppe_if,  
ahb_rx_ppe_if.ppe                 ahb_txppe0_if,  
ahb_rx_ppe_if.ppe                 ahb_txppe1_if,  
egr_ahb_if.egr                    egr_ahb_if,  //EGR-AHB and DFx Interface 
egr_epl_if.egr                    egr_epl0_if,  //EGR-EPL 0 Interface 
egr_epl_if.egr                    egr_epl1_if,  //EGR-EPL 1 Interface 
egr_epl_if.egr                    egr_epl2_if,  //EGR-EPL 2 Interface 
egr_epl_if.egr                    egr_epl3_if,  //EGR-EPL 3 Interface 
egr_igr_if.egr                    egr_igr_if,  //EGR-IGR Pointer Interface 
egr_mc_table_if.egr               egr_mc_table_if0,  //EGR-MultiCast Shared Table 0 Interface 
egr_mc_table_if.egr               egr_mc_table_if1,  //EGR-MultiCast Shared Table 1 Interface 
egr_pod_if.egr                    egr_pod_if,  //EGR-Pod Ring Interface 
egr_ppe_stm_if.egr                egr_ppestm_if0,  //EGR-PPE Shared Table Memory 0 Interface  
egr_ppe_stm_if.egr                egr_ppestm_if1,  //EGR-PPE Shared Table Memory 1 Interface 
egr_smm_readarb_if.egr            egr_smm_readarb_if,  //EGR-SMM_Read_Arb Interface 
egr_smm_writearb_if.egr           egr_smm_writearb_if,  //EGR-SMM_Write_Arb Interface 
egr_statsmgmt_if.egr              egr_statsmgmt_if,  //EGR-Stats Management Interface 
egr_tagring_if.egr                egr_tagring_if,  //EGR-Tag Ring Interface 
egr_vp_if.egr                     egr_vp_if0,  //EGR-VP0 Interface 
egr_vp_if.egr                     egr_vp_if1,  //EGR-VP1 Interface 
glb_rx_ppe_if.ppe                 glb_rx_ppe_if,  
glb_rx_ppe_if.ppe                 glb_txppe0_if,  
glb_rx_ppe_if.ppe                 glb_txppe1_if,  
rx_ppe_ppe_stm_if.ppe             rx_ppe_ppe_stm_if,  

//Output List
output                  igr_vp_tx_pfc_xoff                        //FIXME should this be [1:0] for 2 VP  
);

egr_tx_ppe_if                    egr_txppe0_if();
egr_tx_ppe_if                    egr_txppe1_if();
igr_rx_ppe_if                    igr_rx_ppe_if();
rx_ppe_igr_if                    rx_ppe_igr_if();


// module igr    from igr_top using igr.map 
igr_top    igr(
/* input  logic                */ .clk                         (clk),                                   
/* input  logic                */ .rst_n                       (rst_n),                                 //taken from HLP active low for MBY? 
/* input  logic          [7:0] */ .grp_A_rx_ecc                (epl0_igr_rx_ecc),                       
/* input  logic          [7:0] */ .grp_B_rx_ecc                (epl1_igr_rx_ecc),                       
/* input  logic          [7:0] */ .grp_C_rx_ecc                (epl2_igr_rx_ecc),                       
/* input  logic          [7:0] */ .grp_D_rx_ecc                (epl3_igr_rx_ecc),                       
/* input  logic          [1:0] */ .grp_A_rx_port_num           (epl0_igr_rx_port_num),                  
/* input  logic          [1:0] */ .grp_B_rx_port_num           (epl1_igr_rx_port_num),                  
/* input  logic          [1:0] */ .grp_C_rx_port_num           (epl2_igr_rx_port_num),                  
/* input  logic          [1:0] */ .grp_D_rx_port_num           (epl3_igr_rx_port_num),                  
/* input  logic          [7:0] */ .grp_A_rx_data_valid         (epl0_igr_rx_data_valid),                
/* input  logic          [7:0] */ .grp_B_rx_data_valid         (epl1_igr_rx_data_valid),                
/* input  logic          [7:0] */ .grp_C_rx_data_valid         (epl2_igr_rx_data_valid),                
/* input  logic          [7:0] */ .grp_D_rx_data_valid         (epl3_igr_rx_data_valid),                
/* input  logic         [23:0] */ .grp_A_rx_metadata           (epl0_igr_rx_metadata),                  
/* input  logic         [23:0] */ .grp_B_rx_metadata           (epl1_igr_rx_metadata),                  
/* input  logic         [23:0] */ .grp_C_rx_metadata           (epl2_igr_rx_metadata),                  
/* input  logic         [23:0] */ .grp_D_rx_metadata           (epl3_igr_rx_metadata),                  
/* input  logic         [35:0] */ .grp_A_rx_time_stamp         (epl0_igr_rx_time_stamp),                
/* input  logic         [35:0] */ .grp_B_rx_time_stamp         (epl1_igr_rx_time_stamp),                
/* input  logic         [35:0] */ .grp_C_rx_time_stamp         (epl2_igr_rx_time_stamp),                
/* input  logic         [35:0] */ .grp_D_rx_time_stamp         (epl3_igr_rx_time_stamp),                
/* input  logic    [0:7][71:0] */ .grp_A_rx_data_w_ecc         (epl0_igr_rx_data_w_ecc),                
/* input  logic    [0:7][71:0] */ .grp_B_rx_data_w_ecc         (epl1_igr_rx_data_w_ecc),                
/* input  logic    [0:7][71:0] */ .grp_C_rx_data_w_ecc         (epl2_igr_rx_data_w_ecc),                
/* input  logic    [0:7][71:0] */ .grp_D_rx_data_w_ecc         (epl3_igr_rx_data_w_ecc),                
/* input  logic                */ .grp_A_rx_pfc_xoff           (epl0_igr_rx_pfc_xoff),                  
/* input  logic                */ .grp_B_rx_pfc_xoff           (epl1_igr_rx_pfc_xoff),                  
/* input  logic                */ .grp_C_rx_pfc_xoff           (epl2_igr_rx_pfc_xoff),                  
/* input  logic                */ .grp_D_rx_pfc_xoff           (epl3_igr_rx_pfc_xoff),                  
/* input  logic          [2:0] */ .grp_A_rx_flow_control_tc    (epl0_igr_rx_flow_control_tc),           
/* input  logic          [2:0] */ .grp_B_rx_flow_control_tc    (epl1_igr_rx_flow_control_tc),           
/* input  logic          [2:0] */ .grp_C_rx_flow_control_tc    (epl2_igr_rx_flow_control_tc),           
/* input  logic          [2:0] */ .grp_D_rx_flow_control_tc    (epl3_igr_rx_flow_control_tc),           
/* input  logic          [7:0] */ .vp_rx_ecc                   (igr_vp_rx_ecc),                         
/* input  logic          [1:0] */ .vp_rx_port_num              (igr_vp_rx_port_num),                    
/* input  logic          [7:0] */ .vp_rx_data_valid            (igr_vp_rx_data_valid),                  
/* input  logic         [23:0] */ .vp_rx_metadata              (igr_vp_rx_metadata),                    
/* input  logic         [35:0] */ .vp_rx_time_stamp            (igr_vp_rx_time_stamp),                  
/* input  logic         [19:0] */ .vp_cpp_rx_metadata          (igr_vp_cpp_rx_metadata),                
/* input  logic    [0:7][71:0] */ .vp_rx_data_w_ecc            (igr_vp_rx_data_w_ecc),                  
/* input  logic          [2:0] */ .vp_rx_flow_control_tc       (igr_vp_rx_flow_control_tc),             
/* output logic                */ .vp_tx_pfc_xoff              (igr_vp_tx_pfc_xoff),                    //FIXME should this be [1:0] for 2 VP  
/* Interface rx_ppe_igr_if.igr */ .rx_ppe_igr                  (rx_ppe_igr_if),                         
/* Interface igr_rx_ppe_if.igr */ .igr_rx_ppe                  (igr_rx_ppe_if));                         
// End of module igr from igr_top


// module egr    from egr_top using egr.map 
egr_top    egr(
/* input  logic                      */ .clk                         (clk),                                   
/* input  logic                      */ .arst_n                      (arst_n),                                //Asynchronous negedge reset    
/* Interface egr_igr_if.egr          */ .igr_if                      (egr_igr_if),                            
/* Interface egr_pod_if.egr          */ .pod_if                      (egr_pod_if),                            
/* Interface egr_ahb_if.egr          */ .ahb_if                      (egr_ahb_if),                            
/* Interface egr_smm_writearb_if.egr */ .smm_writearb_if             (egr_smm_writearb_if),                   
/* Interface egr_smm_readarb_if.egr  */ .smm_readarb_if              (egr_smm_readarb_if),                    
/* Interface egr_tagring_if.egr      */ .tagring_if                  (egr_tagring_if),                        
/* Interface egr_statsmgmt_if.egr    */ .statsmgmt_if                (egr_statsmgmt_if),                      
/* Interface egr_tx_ppe_if.egr       */ .tx_ppe_if0                  (egr_txppe0_if),                         
/* Interface egr_tx_ppe_if.egr       */ .tx_ppe_if1                  (egr_txppe1_if),                         
/* Interface egr_ppe_stm_if.egr      */ .ppe_stm_if0                 (egr_ppestm_if0),                        
/* Interface egr_ppe_stm_if.egr      */ .ppe_stm_if1                 (egr_ppestm_if1),                        
/* Interface egr_epl_if.egr          */ .epl_if0                     (egr_epl0_if),                           
/* Interface egr_epl_if.egr          */ .epl_if1                     (egr_epl1_if),                           
/* Interface egr_epl_if.egr          */ .epl_if2                     (egr_epl2_if),                           
/* Interface egr_epl_if.egr          */ .epl_if3                     (egr_epl3_if),                           
/* Interface egr_vp_if.egr           */ .vp_if0                      (egr_vp_if0),                            
/* Interface egr_vp_if.egr           */ .vp_if1                      (egr_vp_if1),                            
/* Interface egr_mc_table_if.egr     */ .mc_table_if0                (egr_mc_table_if0),                      
/* Interface egr_mc_table_if.egr     */ .mc_table_if1                (egr_mc_table_if1));                      
// End of module egr from egr_top


// module rxppe    from rx_ppe using rxppe.map 
rx_ppe    rxppe(
/* Interface rx_ppe_ppe_stm_if.ppe */ .rx_ppe_ppe_stm_if           (rx_ppe_ppe_stm_if),                     
/* Interface rx_ppe_igr_if.ppe     */ .rx_ppe_igr_if               (rx_ppe_igr_if),                         
/* input  logic                    */ .cclk                        (cclk),                                  
/* input  logic                    */ .reset                       (reset),                                 
/* Interface ahb_rx_ppe_if.ppe     */ .ahb_rx_ppe_if               (ahb_rx_ppe_if),                         
/* Interface glb_rx_ppe_if.ppe     */ .glb_rx_ppe_if               (glb_rx_ppe_if),                         
/* Interface igr_rx_ppe_if.ppe     */ .igr_rx_ppe_if               (igr_rx_ppe_if));                         
// End of module rxppe from rx_ppe


// module txppe0    from tx_ppe using txppe.map 0
tx_ppe    txppe0(
/* input  logic                */ .cclk                        (cclk),                                  
/* input  logic                */ .reset                       (reset),                                 
/* Interface ahb_rx_ppe_if.ppe */ .ahb_tx_ppe_if               (ahb_txppe0_if),                         
/* Interface glb_rx_ppe_if.ppe */ .glb_tx_ppe_if               (glb_txppe0_if),                         
/* Interface egr_tx_ppe_if.ppe */ .egr_tx_ppe_if               (egr_txppe0_if));                         
// End of module txppe0 from tx_ppe


// module txppe1    from tx_ppe using txppe.map 1
tx_ppe    txppe1(
/* input  logic                */ .cclk                        (cclk),                                  
/* input  logic                */ .reset                       (reset),                                 
/* Interface ahb_rx_ppe_if.ppe */ .ahb_tx_ppe_if               (ahb_txppe1_if),                         
/* Interface glb_rx_ppe_if.ppe */ .glb_tx_ppe_if               (glb_txppe1_if),                         
/* Interface egr_tx_ppe_if.ppe */ .egr_tx_ppe_if               (egr_txppe1_if));                         
// End of module txppe1 from tx_ppe

endmodule // mgp
