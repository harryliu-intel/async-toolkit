magic
tech scmos
timestamp 965071057
<< ndiffusion >>
rect -16 56 -8 57
rect -16 48 -8 53
rect -16 44 -8 45
<< pdiffusion >>
rect 8 61 16 62
rect 8 57 16 58
rect 16 49 24 54
rect 8 48 24 49
rect 8 44 24 45
<< ntransistor >>
rect -16 53 -8 56
rect -16 45 -8 48
<< ptransistor >>
rect 8 58 16 61
rect 8 45 24 48
<< polysilicon >>
rect 3 58 8 61
rect 16 58 20 61
rect 3 56 6 58
rect -20 53 -16 56
rect -8 53 6 56
rect -20 45 -16 48
rect -8 45 -4 48
rect 4 45 8 48
rect 24 45 28 48
<< ndcontact >>
rect -16 57 -8 65
rect -16 36 -8 44
<< pdcontact >>
rect 8 62 16 70
rect 8 49 16 57
rect 8 36 24 44
<< metal1 >>
rect -16 57 0 65
rect 8 62 16 70
rect -8 49 16 57
rect -16 36 -8 44
rect 8 36 24 44
<< labels >>
rlabel pdcontact 12 40 12 40 5 Vdd!
rlabel ndcontact -12 61 -12 61 4 x
rlabel ndcontact -12 40 -12 40 5 GND!
rlabel space -21 36 -16 65 7 ^n
rlabel polysilicon 17 60 17 60 7 a
rlabel pdcontact 12 66 12 66 5 Vdd!
rlabel pdcontact 12 53 12 53 7 x
rlabel polysilicon -17 54 -17 54 3 a
rlabel polysilicon -17 46 -17 46 3 _SReset!
rlabel polysilicon 25 46 25 46 1 _PReset!
rlabel space 16 56 21 70 3 ^p
<< end >>
