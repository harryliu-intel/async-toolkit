// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

// vim: noai : ts=3 : sw=3 : expandtab : ft=systemverilog

//------------------------------------------------------------------------------
//
// INTEL CONFIDENTIAL
//
// Copyright 2018 Intel Corporation All Rights Reserved.
//
// The source code contained or described herein and all documents related to
// the source code ("Material") are owned by Intel Corporation or its suppliers
// or licensors. Title to the Material remains with Intel Corporation or its
// suppliers and licensors. The Material contains trade secrets and proprietary
// and confidential information of Intel or its suppliers and licensors.  The
// Material is protected by worldwide copyright and trade secret laws and
// treaty provisions. No part of the Material may be used, copied, reproduced,
// modified, published, uploaded, posted, transmitted, distributed, or
// disclosed in any way without Intel's prior express written permission.
//
// No license under any patent, copyright, trade secret or other intellectual
// property right is granted to or conferred upon you by disclosure or delivery
// of the Materials, either expressly, by implication, inducement, estoppel or
// otherwise. Any license under such intellectual property rights must be
// express and approved by Intel in writing.
//
//------------------------------------------------------------------------------
//   Author        : Akshay Kotian
//   Project       : Madison Bay
//------------------------------------------------------------------------------

//   Class:    mby_rx_ppe_base_test
//
//   This is the Base Test file.


`ifndef MBY_RX_PPE_BASE_TEST__SV
`define MBY_RX_PPE_BASE_TEST__SV

`ifndef __INSIDE_MBY_RX_PPE_TEST_LIB
`error "Attempt to include file outside of mby_rx_ppe_test_lib."
`endif

class mby_rx_ppe_base_test extends shdv_base_test;

   // Variable: cfg
   // Top level rx_ppe env configuration
   mby_rx_ppe_tb_top_cfg cfg;

   // Variable: env
   // Top level ENV
   mby_rx_ppe_env    env;

   `uvm_component_utils_begin(mby_rx_ppe_base_test)
      `uvm_field_object(cfg,  UVM_DEFAULT)
      `uvm_field_object(env,      UVM_DEFAULT)
   `uvm_component_utils_end

   //------------------------------------------------------------------------------
   // Constructor: new
   // Configure the TimeFormat - $timeformat(-9, 0, "ns", 10);
   //
   //  Arguments:
   //  name   - rx_ppe base test object name.
   //  parent - Component parent object.
   //------------------------------------------------------------------------------
   function      new(string name = "mby_rx_ppe_base_test", uvm_component parent = null);
      super.new (name, parent);
      $timeformat(-9, 0, "ns", 10);
   endfunction: new

   //------------------------------------------------------------------------------
   // Function: report_phase
   // Checks the Global report server as well as the Test for Errors.  Indicates End_of_Test PASS or FAIL
   //
   //  Arguments:
   //  phase - uvm_phase object.
   //------------------------------------------------------------------------------
   virtual function void report_phase(uvm_phase phase);
      uvm_report_server foo;
      int err_cnt;
      super.report_phase(phase);
      foo = uvm_top.get_report_server();

      // sum num of errors from sequences (use global report server)
      err_cnt = foo.get_severity_count(UVM_ERROR) + foo.get_severity_count(UVM_FATAL);

      // sum num of errors from this test.
      foo = get_report_server();
      err_cnt += (foo.get_severity_count(UVM_ERROR) + foo.get_severity_count(UVM_FATAL));

      if (err_cnt == 0) begin
         uvm_report_info(get_full_name(),  "                                                    ", UVM_LOG);
         uvm_report_info(get_full_name(),  "         _______  _______  _______  _______         ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |       ||   _   ||       ||       |        ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |    _  ||  |_|  ||  _____||  _____|        ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |   |_| ||       || |_____ | |_____         ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |    ___||       ||_____  ||_____  |        ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |   |    |   _   | _____| | _____| |        ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |___|    |__| |__||_______||_______|        ", UVM_LOG);
         uvm_report_info(get_full_name(),  "                                                    ", UVM_LOG);
      end
      else begin
         uvm_report_info(get_full_name(),  "                                                    ", UVM_LOG);
         uvm_report_info(get_full_name(),  "         _______  _______  ___   ___                ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |       ||   _   ||   | |   |               ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |    ___||  |_|  ||   | |   |               ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |   |___ |       ||   | |   |               ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |    ___||       ||   | |   |___            ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |   |    |   _   ||   | |       |           ", UVM_LOG);
         uvm_report_info(get_full_name(),  "        |___|    |__| |__||___| |_______|           ", UVM_LOG);
         uvm_report_info(get_full_name(),  "                                                    ", UVM_LOG);
         uvm_report_info(get_full_name(),  "                                                    ", UVM_LOG);
      end
   endfunction

   //------------------------------------------------------------------------------
   // Function: build_phase
   // Creates cfg, then Randomizes cfg's. Sets the cfg object. Then creates the mby_rx_ppe_env.
   //
   //  Arguments:
   //  phase - uvm_phase object.
   //------------------------------------------------------------------------------
   virtual function void build_phase(uvm_phase phase);
      uvm_report_info(get_full_name(),"Build", UVM_LOG);

      cfg = mby_rx_ppe_tb_top_cfg::type_id::create("cfg", this);                      // Create a Top-Level Configuration object

      randomize_cfg();                                                                // Randomize the Top_Config

      set_config_object("env", "mby_rx_ppe_tb_top_cfg", cfg, 0);

      env     = mby_rx_ppe_env::type_id::create("env",this);                          // Create the Top Environment object
   endfunction : build_phase


   //------------------------------------------------------------------------------
   // Function: connect_phase
   //
   //  Arguments:
   //  phase - uvm_phase object.
   //------------------------------------------------------------------------------
   virtual function void connect_phase(uvm_phase phase);
      super.connect_phase(phase);
      set_default_sequences();

   endfunction : connect_phase

   //-----------------------------------------------------------------------------
   // Function: set_default_sequences()
   //-----------------------------------------------------------------------------
   virtual function void set_default_sequences();        
       
      // Specifying reset phase sequence
      uvm_config_db#(uvm_object_wrapper)::set(this,
         "env.tb_seqr.reset_phase",
         "default_sequence",
         mby_rx_ppe_seq_lib::mby_rx_ppe_hard_reset_seq::type_id::get());

      // Specifying configure phase sequence
      uvm_config_db#(uvm_object_wrapper)::set(this,
         "env.tb_seqr.configure_phase",
         "default_sequence",
         mby_rx_ppe_seq_lib::mby_rx_ppe_env_cfg_seq::type_id::get());

      // Specifying shutdown phase sequence
      uvm_config_db#(uvm_object_wrapper)::set(this,
         "env.tb_seqr.shutdown_phase",
         "default_sequence",
         mby_rx_ppe_seq_lib::mby_rx_ppe_env_shutdown_seq::type_id::get());

   endfunction : set_default_sequences


   //------------------------------------------------------------------------------
   // Function: randomize_cfg()
   // Randomizes the Top_cfg, which will randomizes any sub-level cfg as well.
   //------------------------------------------------------------------------------
   virtual function void randomize_cfg();
      `uvm_info(get_name(), "mby_rx_ppe_base_test randomize_cfg was called!", UVM_HIGH);
      if (!this.randomize(cfg)) begin
         `uvm_fatal(get_name, "randomization of mby_rx_ppe_tb_top_cfg failed");
      end

   endfunction : randomize_cfg

endclass : mby_rx_ppe_base_test

`endif // MBY_RX_PPE_BASE_TEST__SV
