magic
tech scmos
timestamp 962801301
<< ndiffusion >>
rect 5 144 13 145
rect 35 144 43 145
rect 5 136 13 141
rect -17 123 -9 128
rect 5 132 13 133
rect 5 123 13 124
rect 35 136 43 141
rect 35 132 43 133
rect 35 123 43 124
rect -17 112 -9 120
rect 5 115 13 120
rect 35 115 43 120
rect 5 111 13 112
rect 5 102 13 103
rect 35 111 43 112
rect 5 94 13 99
rect 35 94 43 95
rect -25 88 -17 89
rect -25 84 -17 85
rect 5 86 13 91
rect 35 86 43 91
rect 5 82 13 83
rect 5 73 13 74
rect 5 65 13 70
rect 35 82 43 83
rect 35 73 43 74
rect 35 65 43 70
rect 5 57 13 62
rect 35 61 43 62
rect 5 53 13 54
rect 5 44 13 45
rect 35 44 43 45
rect -17 36 -9 44
rect 5 36 13 41
rect 35 36 43 41
rect -17 28 -9 33
rect 5 32 13 33
rect 5 23 13 24
rect 5 15 13 20
rect 35 32 43 33
rect 35 23 43 24
rect 35 15 43 20
rect 5 11 13 12
rect 35 11 43 12
<< pdiffusion >>
rect 59 144 67 145
rect 88 144 100 145
rect 114 144 126 145
rect 59 136 67 141
rect 88 136 100 141
rect 114 140 126 141
rect 59 132 67 133
rect 59 123 67 124
rect 59 115 67 120
rect 88 132 100 133
rect 88 123 100 124
rect 122 135 126 140
rect 88 115 100 120
rect 59 111 67 112
rect 88 111 100 112
rect 59 94 67 95
rect 113 101 129 102
rect 88 94 100 95
rect 113 97 129 98
rect 113 92 118 97
rect 59 86 67 91
rect 59 82 67 83
rect 59 73 67 74
rect 88 86 100 91
rect 126 92 129 97
rect 88 82 100 83
rect 88 73 100 74
rect 59 65 67 70
rect 88 65 100 70
rect 122 66 126 71
rect 114 65 126 66
rect 59 61 67 62
rect 59 44 67 45
rect 88 61 100 62
rect 114 61 126 62
rect 88 44 100 45
rect 59 36 67 41
rect 59 32 67 33
rect 59 23 67 24
rect 88 36 100 41
rect 88 32 100 33
rect 88 23 100 24
rect 59 15 67 20
rect 88 15 100 20
rect 122 16 126 21
rect 114 15 126 16
rect 59 11 67 12
rect 88 11 100 12
rect 114 11 126 12
<< ntransistor >>
rect 5 141 13 144
rect 35 141 43 144
rect 5 133 13 136
rect 35 133 43 136
rect -17 120 -9 123
rect 5 120 13 123
rect 35 120 43 123
rect 5 112 13 115
rect 35 112 43 115
rect 5 99 13 102
rect 5 91 13 94
rect 35 91 43 94
rect -25 85 -17 88
rect 5 83 13 86
rect 35 83 43 86
rect 5 70 13 73
rect 35 70 43 73
rect 5 62 13 65
rect 35 62 43 65
rect 5 54 13 57
rect 5 41 13 44
rect 35 41 43 44
rect -17 33 -9 36
rect 5 33 13 36
rect 35 33 43 36
rect 5 20 13 23
rect 35 20 43 23
rect 5 12 13 15
rect 35 12 43 15
<< ptransistor >>
rect 59 141 67 144
rect 88 141 100 144
rect 114 141 126 144
rect 59 133 67 136
rect 88 133 100 136
rect 59 120 67 123
rect 88 120 100 123
rect 59 112 67 115
rect 88 112 100 115
rect 59 91 67 94
rect 113 98 129 101
rect 88 91 100 94
rect 59 83 67 86
rect 88 83 100 86
rect 59 70 67 73
rect 88 70 100 73
rect 59 62 67 65
rect 88 62 100 65
rect 114 62 126 65
rect 59 41 67 44
rect 88 41 100 44
rect 59 33 67 36
rect 88 33 100 36
rect 59 20 67 23
rect 88 20 100 23
rect 59 12 67 15
rect 88 12 100 15
rect 114 12 126 15
<< polysilicon >>
rect 1 141 5 144
rect 13 141 35 144
rect 43 141 59 144
rect 67 141 88 144
rect 100 141 104 144
rect 110 141 114 144
rect 126 141 131 144
rect 1 133 5 136
rect 13 133 18 136
rect 1 128 3 133
rect 0 123 3 128
rect 23 123 26 141
rect 31 133 35 136
rect 43 133 59 136
rect 67 133 79 136
rect 84 133 88 136
rect 100 133 104 136
rect -19 120 -17 123
rect -9 120 -5 123
rect 0 120 5 123
rect 13 120 18 123
rect 23 120 35 123
rect 43 120 59 123
rect 67 120 71 123
rect 76 115 79 133
rect 102 128 104 133
rect 128 128 131 141
rect 102 123 105 128
rect 84 120 88 123
rect 100 120 105 123
rect 126 125 131 128
rect 1 112 5 115
rect 13 112 35 115
rect 43 112 59 115
rect 67 112 88 115
rect 100 112 104 115
rect 1 99 5 102
rect 13 99 18 102
rect 1 91 5 94
rect 13 91 35 94
rect 43 91 59 94
rect 67 91 74 94
rect 109 98 113 101
rect 129 98 133 101
rect 82 91 88 94
rect 100 91 104 94
rect -29 85 -25 88
rect -17 85 -13 88
rect 0 83 5 86
rect 13 83 18 86
rect 23 83 35 86
rect 43 83 59 86
rect 67 83 71 86
rect 0 78 3 83
rect 1 73 3 78
rect 1 70 5 73
rect 13 70 18 73
rect 23 65 26 83
rect 76 73 79 91
rect 84 83 88 86
rect 100 83 105 86
rect 102 78 105 83
rect 126 78 131 81
rect 102 73 104 78
rect 31 70 35 73
rect 43 70 59 73
rect 67 70 79 73
rect 84 70 88 73
rect 100 70 104 73
rect 128 65 131 78
rect -19 62 5 65
rect 13 62 35 65
rect 43 62 59 65
rect 67 62 88 65
rect 100 62 104 65
rect 110 62 114 65
rect 126 62 131 65
rect 1 54 5 57
rect 13 54 18 57
rect 1 41 5 44
rect 13 41 35 44
rect 43 41 59 44
rect 67 41 88 44
rect 100 41 104 44
rect -19 33 -17 36
rect -9 33 -5 36
rect 0 33 5 36
rect 13 33 18 36
rect 23 33 35 36
rect 43 33 59 36
rect 67 33 71 36
rect 0 28 3 33
rect 1 23 3 28
rect 1 20 5 23
rect 13 20 18 23
rect 23 15 26 33
rect 76 23 79 41
rect 84 33 88 36
rect 100 33 105 36
rect 102 28 105 33
rect 126 28 131 31
rect 102 23 104 28
rect 31 20 35 23
rect 43 20 59 23
rect 67 20 79 23
rect 84 20 88 23
rect 100 20 104 23
rect 128 15 131 28
rect 1 12 5 15
rect 13 12 35 15
rect 43 12 59 15
rect 67 12 88 15
rect 100 12 104 15
rect 110 12 114 15
rect 126 12 131 15
<< ndcontact >>
rect 5 145 13 153
rect 35 145 43 153
rect -17 128 -9 136
rect 5 124 13 132
rect 35 124 43 132
rect -17 104 -9 112
rect 5 103 13 111
rect -25 89 -17 97
rect 35 95 43 111
rect -25 76 -17 84
rect 5 74 13 82
rect 35 74 43 82
rect -17 44 -9 52
rect 5 45 13 53
rect 35 45 43 61
rect -17 20 -9 28
rect 5 24 13 32
rect 35 24 43 32
rect 5 3 13 11
rect 35 3 43 11
<< pdcontact >>
rect 59 145 67 153
rect 88 145 100 153
rect 114 145 126 153
rect 59 124 67 132
rect 88 124 100 132
rect 114 132 122 140
rect 59 95 67 111
rect 88 95 100 111
rect 113 102 129 110
rect 59 74 67 82
rect 118 89 126 97
rect 88 74 100 82
rect 114 66 122 74
rect 59 45 67 61
rect 88 45 100 61
rect 114 53 126 61
rect 59 24 67 32
rect 88 24 100 32
rect 114 16 122 24
rect 59 3 67 11
rect 88 3 100 11
rect 114 3 126 11
<< polycontact >>
rect -7 128 1 136
rect -27 116 -19 124
rect 104 128 112 136
rect 118 120 126 128
rect 74 91 82 99
rect -13 83 -5 91
rect -7 70 1 78
rect -27 62 -19 70
rect 118 78 126 86
rect 104 70 112 78
rect -27 32 -19 40
rect -7 20 1 28
rect 118 28 126 36
rect 104 20 112 28
<< metal1 >>
rect 5 145 43 153
rect 59 145 126 153
rect -4 140 118 141
rect -4 136 122 140
rect -17 128 1 136
rect 104 132 122 136
rect 5 124 100 132
rect 104 128 112 132
rect 118 124 126 128
rect -27 116 13 124
rect -17 111 -9 112
rect -25 104 43 111
rect -25 89 -17 104
rect 5 103 43 104
rect 35 95 43 103
rect 48 91 54 124
rect 96 120 126 124
rect 59 110 100 111
rect 59 103 129 110
rect 59 95 67 103
rect 74 91 82 99
rect 88 95 100 103
rect 113 102 129 103
rect -13 89 -5 91
rect -25 78 -17 84
rect -13 83 13 89
rect 48 86 79 91
rect 118 86 126 97
rect 5 82 13 83
rect 96 82 126 86
rect -25 76 1 78
rect -24 74 1 76
rect 5 74 100 82
rect 118 78 126 82
rect 104 74 112 78
rect -7 70 1 74
rect 104 70 122 74
rect -27 62 -19 70
rect -4 66 122 70
rect -4 65 118 66
rect -27 40 -21 62
rect 35 53 43 61
rect 5 52 43 53
rect -17 45 43 52
rect 59 53 126 61
rect 59 45 67 53
rect 88 45 100 53
rect -17 44 -9 45
rect -27 32 13 40
rect 96 32 126 36
rect -17 20 1 28
rect 5 24 100 32
rect 118 28 126 32
rect 104 24 112 28
rect 104 20 122 24
rect -4 16 122 20
rect -4 15 118 16
rect 5 3 43 11
rect 59 3 126 11
<< labels >>
rlabel metal1 94 149 94 149 5 Vdd!
rlabel metal1 9 149 9 149 5 GND!
rlabel metal1 63 149 63 149 5 Vdd!
rlabel metal1 39 149 39 149 5 GND!
rlabel metal1 94 28 94 28 1 _ab
rlabel metal1 63 28 63 28 1 _ab
rlabel metal1 39 28 39 28 1 _ab
rlabel metal1 9 28 9 28 1 _ab
rlabel polysilicon 101 42 101 42 1 b
rlabel polysilicon 4 13 4 13 1 a
rlabel metal1 120 7 120 7 1 Vdd!
rlabel metal1 94 7 94 7 1 Vdd!
rlabel metal1 9 7 9 7 1 GND!
rlabel metal1 63 7 63 7 1 Vdd!
rlabel metal1 39 7 39 7 1 GND!
rlabel metal1 9 49 9 49 1 GND!
rlabel metal1 39 49 39 49 1 GND!
rlabel metal1 9 107 9 107 5 GND!
rlabel metal1 39 107 39 107 5 GND!
rlabel metal1 122 82 122 82 1 x
rlabel polysilicon 4 55 4 55 1 _SReset!
rlabel polysilicon 4 100 4 100 1 _SReset!
rlabel metal1 120 57 120 57 1 Vdd!
rlabel metal1 94 57 94 57 1 Vdd!
rlabel metal1 94 78 94 78 5 x
rlabel metal1 9 78 9 78 1 x
rlabel metal1 63 57 63 57 1 Vdd!
rlabel metal1 63 78 63 78 1 x
rlabel metal1 39 78 39 78 1 x
rlabel metal1 94 107 94 107 5 Vdd!
rlabel metal1 63 107 63 107 5 Vdd!
rlabel polysilicon 4 143 4 143 5 c
rlabel polysilicon 101 114 101 114 5 d
rlabel metal1 39 128 39 128 5 _cd
rlabel metal1 9 128 9 128 5 _cd
rlabel metal1 63 128 63 128 5 _cd
rlabel metal1 94 128 94 128 5 _cd
rlabel metal1 120 149 120 149 1 Vdd!
rlabel metal1 118 107 118 107 1 Vdd!
rlabel metal1 78 95 78 95 1 _cd
rlabel metal1 -9 87 -9 87 5 x
rlabel ndcontact -13 108 -13 108 5 GND!
rlabel metal1 -21 93 -21 93 1 GND!
rlabel metal1 -23 66 -23 66 1 _ab
rlabel metal1 -13 48 -13 48 1 GND!
rlabel polysilicon 130 99 130 99 7 _PReset!
rlabel space -30 2 36 154 7 ^n
rlabel space 66 2 134 154 3 ^p
rlabel space 67 10 80 46 7 ^pab
rlabel space 22 10 35 46 3 ^nab
rlabel space 22 60 35 96 3 ^nx
rlabel space 67 60 83 100 7 ^px
rlabel space 22 110 35 146 3 ^ncd
rlabel space 67 110 80 146 7 ^pcd
<< end >>
