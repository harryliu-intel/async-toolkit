magic
tech scmos
timestamp 988943070
<< nselect >>
rect -34 483 0 528
<< pselect >>
rect 0 475 46 528
<< ndiffusion >>
rect -28 516 -8 517
rect -28 508 -8 513
rect -28 500 -8 505
rect -28 496 -8 497
<< pdiffusion >>
rect 8 516 40 517
rect 8 512 40 513
rect 8 503 40 504
rect 8 499 40 500
rect 28 491 40 499
rect 8 490 40 491
rect 8 486 40 487
<< ntransistor >>
rect -28 513 -8 516
rect -28 505 -8 508
rect -28 497 -8 500
<< ptransistor >>
rect 8 513 40 516
rect 8 500 40 503
rect 8 487 40 490
<< polysilicon >>
rect -32 513 -28 516
rect -8 513 8 516
rect 40 513 44 516
rect -32 505 -28 508
rect -8 505 6 508
rect 3 503 6 505
rect 3 500 8 503
rect 40 500 44 503
rect -32 497 -28 500
rect -8 497 -2 500
rect -5 490 -2 497
rect -5 487 8 490
rect 40 487 44 490
<< ndcontact >>
rect -28 517 -8 525
rect -28 488 -8 496
<< pdcontact >>
rect 8 517 40 525
rect 8 504 40 512
rect 8 491 28 499
rect 8 478 40 486
<< metal1 >>
rect -28 517 40 525
rect -4 499 4 517
rect 8 504 40 512
rect -28 488 -8 496
rect -4 491 28 499
rect 32 486 40 504
rect 8 478 40 486
<< labels >>
rlabel space -35 475 -28 528 7 ^n
rlabel space 28 475 47 528 3 ^p
rlabel metal1 -28 488 -8 496 1 GND!|pin|s|0
rlabel metal1 32 478 40 512 1 Vdd!|pin|s|1
rlabel metal1 -4 491 4 525 1 x|pin|s|2
rlabel metal1 -28 517 40 525 1 x|pin|s|2
rlabel metal1 -4 491 28 499 1 x|pin|s|2
rlabel polysilicon 40 487 44 490 1 a|pin|w|3|poly
rlabel polysilicon -2 487 2 490 1 a|pin|w|3|poly
rlabel polysilicon -32 497 -28 500 1 a|pin|w|3|poly
rlabel polysilicon -32 505 -28 508 1 b|pin|w|4|poly
rlabel polysilicon 40 500 44 503 1 b|pin|w|4|poly
rlabel polysilicon 40 513 44 516 1 c|pin|w|5|poly
rlabel polysilicon -1 513 3 516 1 c|pin|w|5|poly
rlabel polysilicon -32 513 -28 516 1 c|pin|w|5|poly
rlabel metal1 8 478 40 486 1 Vdd!|pin|s|1
rlabel metal1 8 504 40 512 1 Vdd!|pin|s|1
<< end >>
