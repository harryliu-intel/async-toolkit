package mby_mesh_bfm_pkg;

   `include "uvm_macros.svh"
   `include "slu_macros.svh"
   import uvm_pkg::*;
   import shdv_base_pkg::*;

   `include "mby_mesh_defines.svh"
   `include "mby_mesh_mem_crdt_io.sv"
   `include "mby_mesh_flow_ctrl.sv"
   `include "mby_mesh_agent_cfg.sv"
   `include "mby_mesh_req_agent_cfg.sv"
   `include "mby_mesh_req_seq_item.sv"
   `include "mby_mesh_rdreq_drv.sv"
   `include "mby_mesh_rdreq_mon.sv"
   `include "mby_mesh_rdreq_agent.sv"
   `include "mby_mesh_wrreq_drv.sv"
   `include "mby_mesh_wrreq_mon.sv"
   `include "mby_mesh_wrreq_agent.sv"
   `include "mby_mesh_rdrsp_drv.sv"
   `include "mby_mesh_rdrsp_mon.sv"
   `include "mby_mesh_rdrsp_agent.sv"
   `include "mby_mesh_agent.sv"
   `include "mby_mesh_bfm.sv"

endpackage