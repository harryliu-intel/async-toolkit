///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_modify_map.sv                                      
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_modify_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_FF
`define RTLGEN_MBY_PPE_MODIFY_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_FF

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF
`define RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_MODIFY_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_FF_RSTD


module rtlgen_mby_ppe_modify_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_modify_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_MODIFY_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_MODIFY_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_MODIFY_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_MODIFY_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_PH2_FF
`define RTLGEN_MBY_PPE_MODIFY_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_MODIFY_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_MODIFY_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_LATCH
`define RTLGEN_MBY_PPE_MODIFY_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_MODIFY_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_MODIFY_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_modify_map ( //lintra s-2096
    // Clocks
    gated_clk,

    // Resets
    rst_n,


    // Register Inputs
    handcode_reg_rdata_MOD_CSUM_CFG1,
    handcode_reg_rdata_MOD_CSUM_CFG2,
    handcode_reg_rdata_MOD_MAP,
    handcode_reg_rdata_MOD_MAP_CFG,
    handcode_reg_rdata_MOD_MAP_DUAL,
    handcode_reg_rdata_MOD_MAP_DUAL_CFG,
    handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE0,
    handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE1,
    handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE2,
    handcode_reg_rdata_MOD_PROFILE_COMMAND,
    handcode_reg_rdata_MOD_PROFILE_FIELD,
    handcode_reg_rdata_MOD_PROFILE_GROUP,

    handcode_rvalid_MOD_CSUM_CFG1,
    handcode_rvalid_MOD_CSUM_CFG2,
    handcode_rvalid_MOD_MAP,
    handcode_rvalid_MOD_MAP_CFG,
    handcode_rvalid_MOD_MAP_DUAL,
    handcode_rvalid_MOD_MAP_DUAL_CFG,
    handcode_rvalid_MOD_MIRROR_PROFILE_TABLE0,
    handcode_rvalid_MOD_MIRROR_PROFILE_TABLE1,
    handcode_rvalid_MOD_MIRROR_PROFILE_TABLE2,
    handcode_rvalid_MOD_PROFILE_COMMAND,
    handcode_rvalid_MOD_PROFILE_FIELD,
    handcode_rvalid_MOD_PROFILE_GROUP,

    handcode_wvalid_MOD_CSUM_CFG1,
    handcode_wvalid_MOD_CSUM_CFG2,
    handcode_wvalid_MOD_MAP,
    handcode_wvalid_MOD_MAP_CFG,
    handcode_wvalid_MOD_MAP_DUAL,
    handcode_wvalid_MOD_MAP_DUAL_CFG,
    handcode_wvalid_MOD_MIRROR_PROFILE_TABLE0,
    handcode_wvalid_MOD_MIRROR_PROFILE_TABLE1,
    handcode_wvalid_MOD_MIRROR_PROFILE_TABLE2,
    handcode_wvalid_MOD_PROFILE_COMMAND,
    handcode_wvalid_MOD_PROFILE_FIELD,
    handcode_wvalid_MOD_PROFILE_GROUP,

    handcode_error_MOD_CSUM_CFG1,
    handcode_error_MOD_CSUM_CFG2,
    handcode_error_MOD_MAP,
    handcode_error_MOD_MAP_CFG,
    handcode_error_MOD_MAP_DUAL,
    handcode_error_MOD_MAP_DUAL_CFG,
    handcode_error_MOD_MIRROR_PROFILE_TABLE0,
    handcode_error_MOD_MIRROR_PROFILE_TABLE1,
    handcode_error_MOD_MIRROR_PROFILE_TABLE2,
    handcode_error_MOD_PROFILE_COMMAND,
    handcode_error_MOD_PROFILE_FIELD,
    handcode_error_MOD_PROFILE_GROUP,


    // Register Outputs
    MOD_CSUM_EN_CFG,


    // Register signals for HandCoded registers
    handcode_reg_wdata_MOD_CSUM_CFG1,
    handcode_reg_wdata_MOD_CSUM_CFG2,
    handcode_reg_wdata_MOD_MAP,
    handcode_reg_wdata_MOD_MAP_CFG,
    handcode_reg_wdata_MOD_MAP_DUAL,
    handcode_reg_wdata_MOD_MAP_DUAL_CFG,
    handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE0,
    handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE1,
    handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE2,
    handcode_reg_wdata_MOD_PROFILE_COMMAND,
    handcode_reg_wdata_MOD_PROFILE_FIELD,
    handcode_reg_wdata_MOD_PROFILE_GROUP,

    we_MOD_CSUM_CFG1,
    we_MOD_CSUM_CFG2,
    we_MOD_MAP,
    we_MOD_MAP_CFG,
    we_MOD_MAP_DUAL,
    we_MOD_MAP_DUAL_CFG,
    we_MOD_MIRROR_PROFILE_TABLE0,
    we_MOD_MIRROR_PROFILE_TABLE1,
    we_MOD_MIRROR_PROFILE_TABLE2,
    we_MOD_PROFILE_COMMAND,
    we_MOD_PROFILE_FIELD,
    we_MOD_PROFILE_GROUP,

    re_MOD_CSUM_CFG1,
    re_MOD_CSUM_CFG2,
    re_MOD_MAP,
    re_MOD_MAP_CFG,
    re_MOD_MAP_DUAL,
    re_MOD_MAP_DUAL_CFG,
    re_MOD_MIRROR_PROFILE_TABLE0,
    re_MOD_MIRROR_PROFILE_TABLE1,
    re_MOD_MIRROR_PROFILE_TABLE2,
    re_MOD_PROFILE_COMMAND,
    re_MOD_PROFILE_FIELD,
    re_MOD_PROFILE_GROUP,




    // Config Access
    req,
    ack
    

);

import mby_ppe_modify_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:0] MBY_PPE_MODIFY_MAP_OFFSET = {MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] MODIFY_SB_BAR = 3'b0;
parameter [7:0] MODIFY_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
localparam [MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] MOD_CSUM_EN_CFG_DECODE_ADDR = MOD_CSUM_EN_CFG_CR_ADDR[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_MODIFY_MAP_OFFSET[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];

    // Clocks
input logic  gated_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input MOD_CSUM_CFG1_t  handcode_reg_rdata_MOD_CSUM_CFG1;
input MOD_CSUM_CFG2_t  handcode_reg_rdata_MOD_CSUM_CFG2;
input MOD_MAP_t  handcode_reg_rdata_MOD_MAP;
input MOD_MAP_CFG_t  handcode_reg_rdata_MOD_MAP_CFG;
input MOD_MAP_DUAL_t  handcode_reg_rdata_MOD_MAP_DUAL;
input MOD_MAP_DUAL_CFG_t  handcode_reg_rdata_MOD_MAP_DUAL_CFG;
input MOD_MIRROR_PROFILE_TABLE0_t  handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE0;
input MOD_MIRROR_PROFILE_TABLE1_t  handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE1;
input MOD_MIRROR_PROFILE_TABLE2_t  handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE2;
input MOD_PROFILE_COMMAND_t  handcode_reg_rdata_MOD_PROFILE_COMMAND;
input MOD_PROFILE_FIELD_t  handcode_reg_rdata_MOD_PROFILE_FIELD;
input MOD_PROFILE_GROUP_t  handcode_reg_rdata_MOD_PROFILE_GROUP;

input handcode_rvalid_MOD_CSUM_CFG1_t  handcode_rvalid_MOD_CSUM_CFG1;
input handcode_rvalid_MOD_CSUM_CFG2_t  handcode_rvalid_MOD_CSUM_CFG2;
input handcode_rvalid_MOD_MAP_t  handcode_rvalid_MOD_MAP;
input handcode_rvalid_MOD_MAP_CFG_t  handcode_rvalid_MOD_MAP_CFG;
input handcode_rvalid_MOD_MAP_DUAL_t  handcode_rvalid_MOD_MAP_DUAL;
input handcode_rvalid_MOD_MAP_DUAL_CFG_t  handcode_rvalid_MOD_MAP_DUAL_CFG;
input handcode_rvalid_MOD_MIRROR_PROFILE_TABLE0_t  handcode_rvalid_MOD_MIRROR_PROFILE_TABLE0;
input handcode_rvalid_MOD_MIRROR_PROFILE_TABLE1_t  handcode_rvalid_MOD_MIRROR_PROFILE_TABLE1;
input handcode_rvalid_MOD_MIRROR_PROFILE_TABLE2_t  handcode_rvalid_MOD_MIRROR_PROFILE_TABLE2;
input handcode_rvalid_MOD_PROFILE_COMMAND_t  handcode_rvalid_MOD_PROFILE_COMMAND;
input handcode_rvalid_MOD_PROFILE_FIELD_t  handcode_rvalid_MOD_PROFILE_FIELD;
input handcode_rvalid_MOD_PROFILE_GROUP_t  handcode_rvalid_MOD_PROFILE_GROUP;

input handcode_wvalid_MOD_CSUM_CFG1_t  handcode_wvalid_MOD_CSUM_CFG1;
input handcode_wvalid_MOD_CSUM_CFG2_t  handcode_wvalid_MOD_CSUM_CFG2;
input handcode_wvalid_MOD_MAP_t  handcode_wvalid_MOD_MAP;
input handcode_wvalid_MOD_MAP_CFG_t  handcode_wvalid_MOD_MAP_CFG;
input handcode_wvalid_MOD_MAP_DUAL_t  handcode_wvalid_MOD_MAP_DUAL;
input handcode_wvalid_MOD_MAP_DUAL_CFG_t  handcode_wvalid_MOD_MAP_DUAL_CFG;
input handcode_wvalid_MOD_MIRROR_PROFILE_TABLE0_t  handcode_wvalid_MOD_MIRROR_PROFILE_TABLE0;
input handcode_wvalid_MOD_MIRROR_PROFILE_TABLE1_t  handcode_wvalid_MOD_MIRROR_PROFILE_TABLE1;
input handcode_wvalid_MOD_MIRROR_PROFILE_TABLE2_t  handcode_wvalid_MOD_MIRROR_PROFILE_TABLE2;
input handcode_wvalid_MOD_PROFILE_COMMAND_t  handcode_wvalid_MOD_PROFILE_COMMAND;
input handcode_wvalid_MOD_PROFILE_FIELD_t  handcode_wvalid_MOD_PROFILE_FIELD;
input handcode_wvalid_MOD_PROFILE_GROUP_t  handcode_wvalid_MOD_PROFILE_GROUP;

input handcode_error_MOD_CSUM_CFG1_t  handcode_error_MOD_CSUM_CFG1;
input handcode_error_MOD_CSUM_CFG2_t  handcode_error_MOD_CSUM_CFG2;
input handcode_error_MOD_MAP_t  handcode_error_MOD_MAP;
input handcode_error_MOD_MAP_CFG_t  handcode_error_MOD_MAP_CFG;
input handcode_error_MOD_MAP_DUAL_t  handcode_error_MOD_MAP_DUAL;
input handcode_error_MOD_MAP_DUAL_CFG_t  handcode_error_MOD_MAP_DUAL_CFG;
input handcode_error_MOD_MIRROR_PROFILE_TABLE0_t  handcode_error_MOD_MIRROR_PROFILE_TABLE0;
input handcode_error_MOD_MIRROR_PROFILE_TABLE1_t  handcode_error_MOD_MIRROR_PROFILE_TABLE1;
input handcode_error_MOD_MIRROR_PROFILE_TABLE2_t  handcode_error_MOD_MIRROR_PROFILE_TABLE2;
input handcode_error_MOD_PROFILE_COMMAND_t  handcode_error_MOD_PROFILE_COMMAND;
input handcode_error_MOD_PROFILE_FIELD_t  handcode_error_MOD_PROFILE_FIELD;
input handcode_error_MOD_PROFILE_GROUP_t  handcode_error_MOD_PROFILE_GROUP;


    // Register Outputs
output MOD_CSUM_EN_CFG_t  MOD_CSUM_EN_CFG;


    // Register signals for HandCoded registers
output MOD_CSUM_CFG1_t  handcode_reg_wdata_MOD_CSUM_CFG1;
output MOD_CSUM_CFG2_t  handcode_reg_wdata_MOD_CSUM_CFG2;
output MOD_MAP_t  handcode_reg_wdata_MOD_MAP;
output MOD_MAP_CFG_t  handcode_reg_wdata_MOD_MAP_CFG;
output MOD_MAP_DUAL_t  handcode_reg_wdata_MOD_MAP_DUAL;
output MOD_MAP_DUAL_CFG_t  handcode_reg_wdata_MOD_MAP_DUAL_CFG;
output MOD_MIRROR_PROFILE_TABLE0_t  handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE0;
output MOD_MIRROR_PROFILE_TABLE1_t  handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE1;
output MOD_MIRROR_PROFILE_TABLE2_t  handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE2;
output MOD_PROFILE_COMMAND_t  handcode_reg_wdata_MOD_PROFILE_COMMAND;
output MOD_PROFILE_FIELD_t  handcode_reg_wdata_MOD_PROFILE_FIELD;
output MOD_PROFILE_GROUP_t  handcode_reg_wdata_MOD_PROFILE_GROUP;

output we_MOD_CSUM_CFG1_t  we_MOD_CSUM_CFG1;
output we_MOD_CSUM_CFG2_t  we_MOD_CSUM_CFG2;
output we_MOD_MAP_t  we_MOD_MAP;
output we_MOD_MAP_CFG_t  we_MOD_MAP_CFG;
output we_MOD_MAP_DUAL_t  we_MOD_MAP_DUAL;
output we_MOD_MAP_DUAL_CFG_t  we_MOD_MAP_DUAL_CFG;
output we_MOD_MIRROR_PROFILE_TABLE0_t  we_MOD_MIRROR_PROFILE_TABLE0;
output we_MOD_MIRROR_PROFILE_TABLE1_t  we_MOD_MIRROR_PROFILE_TABLE1;
output we_MOD_MIRROR_PROFILE_TABLE2_t  we_MOD_MIRROR_PROFILE_TABLE2;
output we_MOD_PROFILE_COMMAND_t  we_MOD_PROFILE_COMMAND;
output we_MOD_PROFILE_FIELD_t  we_MOD_PROFILE_FIELD;
output we_MOD_PROFILE_GROUP_t  we_MOD_PROFILE_GROUP;

output re_MOD_CSUM_CFG1_t  re_MOD_CSUM_CFG1;
output re_MOD_CSUM_CFG2_t  re_MOD_CSUM_CFG2;
output re_MOD_MAP_t  re_MOD_MAP;
output re_MOD_MAP_CFG_t  re_MOD_MAP_CFG;
output re_MOD_MAP_DUAL_t  re_MOD_MAP_DUAL;
output re_MOD_MAP_DUAL_CFG_t  re_MOD_MAP_DUAL_CFG;
output re_MOD_MIRROR_PROFILE_TABLE0_t  re_MOD_MIRROR_PROFILE_TABLE0;
output re_MOD_MIRROR_PROFILE_TABLE1_t  re_MOD_MIRROR_PROFILE_TABLE1;
output re_MOD_MIRROR_PROFILE_TABLE2_t  re_MOD_MIRROR_PROFILE_TABLE2;
output re_MOD_PROFILE_COMMAND_t  re_MOD_PROFILE_COMMAND;
output re_MOD_PROFILE_FIELD_t  re_MOD_PROFILE_FIELD;
output re_MOD_PROFILE_GROUP_t  re_MOD_PROFILE_GROUP;




    // Config Access
input mby_ppe_modify_map_cr_req_t  req;
output mby_ppe_modify_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_modify_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_MODIFY_MAP_MEM;
assign case_req_addr_MBY_PPE_MODIFY_MAP_MEM = req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_modify;
always_comb begin : sb_fid_cond_modify_BLOCK
    unique casez (req_fid) 
		MODIFY_SB_FID: sb_fid_cond_modify = 1;
		default: sb_fid_cond_modify = 0;
    endcase 
end


logic sb_bar_cond_modify;
always_comb begin : sb_bar_cond_modify_BLOCK
    unique casez (req_bar) 
		MODIFY_SB_BAR: sb_bar_cond_modify = 1;
		default: sb_bar_cond_modify = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// MOD_PROFILE_COMMAND using HANDCODED_REG template.
logic addr_decode_MOD_PROFILE_COMMAND;
logic write_req_MOD_PROFILE_COMMAND;
logic read_req_MOD_PROFILE_COMMAND;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'b0?,8'h??,1'b?}: 
         addr_decode_MOD_PROFILE_COMMAND = req.valid;
      default: 
         addr_decode_MOD_PROFILE_COMMAND = 1'b0; 
   endcase
end

always_comb write_req_MOD_PROFILE_COMMAND = f_IsMEMWr(req_opcode) && addr_decode_MOD_PROFILE_COMMAND ;
always_comb read_req_MOD_PROFILE_COMMAND  = f_IsMEMRd(req_opcode) && addr_decode_MOD_PROFILE_COMMAND ;

always_comb we_MOD_PROFILE_COMMAND = {8{write_req_MOD_PROFILE_COMMAND}} & be;
always_comb re_MOD_PROFILE_COMMAND = {8{read_req_MOD_PROFILE_COMMAND}} & be;
always_comb handcode_reg_wdata_MOD_PROFILE_COMMAND = write_data;


// ----------------------------------------------------------------------
// MOD_PROFILE_FIELD using HANDCODED_REG template.
logic addr_decode_MOD_PROFILE_FIELD;
logic write_req_MOD_PROFILE_FIELD;
logic read_req_MOD_PROFILE_FIELD;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h2??,1'b?}: 
         addr_decode_MOD_PROFILE_FIELD = req.valid;
      default: 
         addr_decode_MOD_PROFILE_FIELD = 1'b0; 
   endcase
end

always_comb write_req_MOD_PROFILE_FIELD = f_IsMEMWr(req_opcode) && addr_decode_MOD_PROFILE_FIELD ;
always_comb read_req_MOD_PROFILE_FIELD  = f_IsMEMRd(req_opcode) && addr_decode_MOD_PROFILE_FIELD ;

always_comb we_MOD_PROFILE_FIELD = {8{write_req_MOD_PROFILE_FIELD}} & be;
always_comb re_MOD_PROFILE_FIELD = {8{read_req_MOD_PROFILE_FIELD}} & be;
always_comb handcode_reg_wdata_MOD_PROFILE_FIELD = write_data;


// ----------------------------------------------------------------------
// MOD_MAP_DUAL using HANDCODED_REG template.
logic addr_decode_MOD_MAP_DUAL;
logic write_req_MOD_MAP_DUAL;
logic read_req_MOD_MAP_DUAL;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h1???,1'b?}: 
         addr_decode_MOD_MAP_DUAL = req.valid;
      default: 
         addr_decode_MOD_MAP_DUAL = 1'b0; 
   endcase
end

always_comb write_req_MOD_MAP_DUAL = f_IsMEMWr(req_opcode) && addr_decode_MOD_MAP_DUAL ;
always_comb read_req_MOD_MAP_DUAL  = f_IsMEMRd(req_opcode) && addr_decode_MOD_MAP_DUAL ;

always_comb we_MOD_MAP_DUAL = {8{write_req_MOD_MAP_DUAL}} & be;
always_comb re_MOD_MAP_DUAL = {8{read_req_MOD_MAP_DUAL}} & be;
always_comb handcode_reg_wdata_MOD_MAP_DUAL = write_data;


// ----------------------------------------------------------------------
// MOD_MAP using HANDCODED_REG template.
logic addr_decode_MOD_MAP;
logic write_req_MOD_MAP;
logic read_req_MOD_MAP;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h2,4'b00??,8'h??,1'b?}: 
         addr_decode_MOD_MAP = req.valid;
      default: 
         addr_decode_MOD_MAP = 1'b0; 
   endcase
end

always_comb write_req_MOD_MAP = f_IsMEMWr(req_opcode) && addr_decode_MOD_MAP ;
always_comb read_req_MOD_MAP  = f_IsMEMRd(req_opcode) && addr_decode_MOD_MAP ;

always_comb we_MOD_MAP = {8{write_req_MOD_MAP}} & be;
always_comb re_MOD_MAP = {8{read_req_MOD_MAP}} & be;
always_comb handcode_reg_wdata_MOD_MAP = write_data;


// ----------------------------------------------------------------------
// MOD_PROFILE_GROUP using HANDCODED_REG template.
logic addr_decode_MOD_PROFILE_GROUP;
logic write_req_MOD_PROFILE_GROUP;
logic read_req_MOD_PROFILE_GROUP;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h24,4'b000?,4'h?,1'b?}: 
         addr_decode_MOD_PROFILE_GROUP = req.valid;
      default: 
         addr_decode_MOD_PROFILE_GROUP = 1'b0; 
   endcase
end

always_comb write_req_MOD_PROFILE_GROUP = f_IsMEMWr(req_opcode) && addr_decode_MOD_PROFILE_GROUP ;
always_comb read_req_MOD_PROFILE_GROUP  = f_IsMEMRd(req_opcode) && addr_decode_MOD_PROFILE_GROUP ;

always_comb we_MOD_PROFILE_GROUP = {8{write_req_MOD_PROFILE_GROUP}} & be;
always_comb re_MOD_PROFILE_GROUP = {8{read_req_MOD_PROFILE_GROUP}} & be;
always_comb handcode_reg_wdata_MOD_PROFILE_GROUP = write_data;


// ----------------------------------------------------------------------
// MOD_MIRROR_PROFILE_TABLE0 using HANDCODED_REG template.
logic addr_decode_MOD_MIRROR_PROFILE_TABLE0;
logic write_req_MOD_MIRROR_PROFILE_TABLE0;
logic read_req_MOD_MIRROR_PROFILE_TABLE0;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h24,4'b001?,4'h?,1'b?}: 
         addr_decode_MOD_MIRROR_PROFILE_TABLE0 = req.valid;
      default: 
         addr_decode_MOD_MIRROR_PROFILE_TABLE0 = 1'b0; 
   endcase
end

always_comb write_req_MOD_MIRROR_PROFILE_TABLE0 = f_IsMEMWr(req_opcode) && addr_decode_MOD_MIRROR_PROFILE_TABLE0 ;
always_comb read_req_MOD_MIRROR_PROFILE_TABLE0  = f_IsMEMRd(req_opcode) && addr_decode_MOD_MIRROR_PROFILE_TABLE0 ;

always_comb we_MOD_MIRROR_PROFILE_TABLE0 = {8{write_req_MOD_MIRROR_PROFILE_TABLE0}} & be;
always_comb re_MOD_MIRROR_PROFILE_TABLE0 = {8{read_req_MOD_MIRROR_PROFILE_TABLE0}} & be;
always_comb handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE0 = write_data;


// ----------------------------------------------------------------------
// MOD_MIRROR_PROFILE_TABLE1 using HANDCODED_REG template.
logic addr_decode_MOD_MIRROR_PROFILE_TABLE1;
logic write_req_MOD_MIRROR_PROFILE_TABLE1;
logic read_req_MOD_MIRROR_PROFILE_TABLE1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h24,4'b010?,4'h?,1'b?}: 
         addr_decode_MOD_MIRROR_PROFILE_TABLE1 = req.valid;
      default: 
         addr_decode_MOD_MIRROR_PROFILE_TABLE1 = 1'b0; 
   endcase
end

always_comb write_req_MOD_MIRROR_PROFILE_TABLE1 = f_IsMEMWr(req_opcode) && addr_decode_MOD_MIRROR_PROFILE_TABLE1 ;
always_comb read_req_MOD_MIRROR_PROFILE_TABLE1  = f_IsMEMRd(req_opcode) && addr_decode_MOD_MIRROR_PROFILE_TABLE1 ;

always_comb we_MOD_MIRROR_PROFILE_TABLE1 = {8{write_req_MOD_MIRROR_PROFILE_TABLE1}} & be;
always_comb re_MOD_MIRROR_PROFILE_TABLE1 = {8{read_req_MOD_MIRROR_PROFILE_TABLE1}} & be;
always_comb handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE1 = write_data;


// ----------------------------------------------------------------------
// MOD_MIRROR_PROFILE_TABLE2 using HANDCODED_REG template.
logic addr_decode_MOD_MIRROR_PROFILE_TABLE2;
logic write_req_MOD_MIRROR_PROFILE_TABLE2;
logic read_req_MOD_MIRROR_PROFILE_TABLE2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h24,4'b011?,4'h?,1'b?}: 
         addr_decode_MOD_MIRROR_PROFILE_TABLE2 = req.valid;
      default: 
         addr_decode_MOD_MIRROR_PROFILE_TABLE2 = 1'b0; 
   endcase
end

always_comb write_req_MOD_MIRROR_PROFILE_TABLE2 = f_IsMEMWr(req_opcode) && addr_decode_MOD_MIRROR_PROFILE_TABLE2 ;
always_comb read_req_MOD_MIRROR_PROFILE_TABLE2  = f_IsMEMRd(req_opcode) && addr_decode_MOD_MIRROR_PROFILE_TABLE2 ;

always_comb we_MOD_MIRROR_PROFILE_TABLE2 = {8{write_req_MOD_MIRROR_PROFILE_TABLE2}} & be;
always_comb re_MOD_MIRROR_PROFILE_TABLE2 = {8{read_req_MOD_MIRROR_PROFILE_TABLE2}} & be;
always_comb handcode_reg_wdata_MOD_MIRROR_PROFILE_TABLE2 = write_data;


// ----------------------------------------------------------------------
// MOD_MAP_CFG using HANDCODED_REG template.
logic addr_decode_MOD_MAP_CFG;
logic write_req_MOD_MAP_CFG;
logic read_req_MOD_MAP_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {40'h248,4'b000?,1'b?}: 
         addr_decode_MOD_MAP_CFG = req.valid;
      default: 
         addr_decode_MOD_MAP_CFG = 1'b0; 
   endcase
end

always_comb write_req_MOD_MAP_CFG = f_IsMEMWr(req_opcode) && addr_decode_MOD_MAP_CFG ;
always_comb read_req_MOD_MAP_CFG  = f_IsMEMRd(req_opcode) && addr_decode_MOD_MAP_CFG ;

always_comb we_MOD_MAP_CFG = {8{write_req_MOD_MAP_CFG}} & be;
always_comb re_MOD_MAP_CFG = {8{read_req_MOD_MAP_CFG}} & be;
always_comb handcode_reg_wdata_MOD_MAP_CFG = write_data;


// ----------------------------------------------------------------------
// MOD_MAP_DUAL_CFG using HANDCODED_REG template.
logic addr_decode_MOD_MAP_DUAL_CFG;
logic write_req_MOD_MAP_DUAL_CFG;
logic read_req_MOD_MAP_DUAL_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h2482,1'b0}: 
         addr_decode_MOD_MAP_DUAL_CFG = req.valid;
      default: 
         addr_decode_MOD_MAP_DUAL_CFG = 1'b0; 
   endcase
end

always_comb write_req_MOD_MAP_DUAL_CFG = f_IsMEMWr(req_opcode) && addr_decode_MOD_MAP_DUAL_CFG ;
always_comb read_req_MOD_MAP_DUAL_CFG  = f_IsMEMRd(req_opcode) && addr_decode_MOD_MAP_DUAL_CFG ;

always_comb we_MOD_MAP_DUAL_CFG = {8{write_req_MOD_MAP_DUAL_CFG}} & be;
always_comb re_MOD_MAP_DUAL_CFG = {8{read_req_MOD_MAP_DUAL_CFG}} & be;
always_comb handcode_reg_wdata_MOD_MAP_DUAL_CFG = write_data;


// ----------------------------------------------------------------------
// MOD_CSUM_CFG1 using HANDCODED_REG template.
logic addr_decode_MOD_CSUM_CFG1;
logic write_req_MOD_CSUM_CFG1;
logic read_req_MOD_CSUM_CFG1;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h2482,1'b1}: 
         addr_decode_MOD_CSUM_CFG1 = req.valid;
      default: 
         addr_decode_MOD_CSUM_CFG1 = 1'b0; 
   endcase
end

always_comb write_req_MOD_CSUM_CFG1 = f_IsMEMWr(req_opcode) && addr_decode_MOD_CSUM_CFG1 ;
always_comb read_req_MOD_CSUM_CFG1  = f_IsMEMRd(req_opcode) && addr_decode_MOD_CSUM_CFG1 ;

always_comb we_MOD_CSUM_CFG1 = {8{write_req_MOD_CSUM_CFG1}} & be;
always_comb re_MOD_CSUM_CFG1 = {8{read_req_MOD_CSUM_CFG1}} & be;
always_comb handcode_reg_wdata_MOD_CSUM_CFG1 = write_data;


// ----------------------------------------------------------------------
// MOD_CSUM_CFG2 using HANDCODED_REG template.
logic addr_decode_MOD_CSUM_CFG2;
logic write_req_MOD_CSUM_CFG2;
logic read_req_MOD_CSUM_CFG2;

always_comb begin 
   unique casez (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {44'h2483,1'b0}: 
         addr_decode_MOD_CSUM_CFG2 = req.valid;
      default: 
         addr_decode_MOD_CSUM_CFG2 = 1'b0; 
   endcase
end

always_comb write_req_MOD_CSUM_CFG2 = f_IsMEMWr(req_opcode) && addr_decode_MOD_CSUM_CFG2 ;
always_comb read_req_MOD_CSUM_CFG2  = f_IsMEMRd(req_opcode) && addr_decode_MOD_CSUM_CFG2 ;

always_comb we_MOD_CSUM_CFG2 = {8{write_req_MOD_CSUM_CFG2}} & be;
always_comb re_MOD_CSUM_CFG2 = {8{read_req_MOD_CSUM_CFG2}} & be;
always_comb handcode_reg_wdata_MOD_CSUM_CFG2 = write_data;


//---------------------------------------------------------------------
// MOD_CSUM_EN_CFG Address Decode
logic  addr_decode_MOD_CSUM_EN_CFG;
logic  write_req_MOD_CSUM_EN_CFG;
always_comb begin
   addr_decode_MOD_CSUM_EN_CFG = (req_addr[MBY_PPE_MODIFY_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == MOD_CSUM_EN_CFG_DECODE_ADDR) && req.valid ;
   write_req_MOD_CSUM_EN_CFG = IsMEMWr && addr_decode_MOD_CSUM_EN_CFG && sb_fid_cond_modify && sb_bar_cond_modify;
end

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D0_IPV4_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D0_IPV4_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D0_IPV4_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D0_IPV4_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D0_IPV4_EN = write_data[0:0];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D0_IPV4_EN[0], nxt_MOD_CSUM_EN_CFG_D0_IPV4_EN[0:0], MOD_CSUM_EN_CFG.D0_IPV4_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D1_IPV4_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D1_IPV4_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D1_IPV4_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D1_IPV4_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D1_IPV4_EN = write_data[1:1];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D1_IPV4_EN[0], nxt_MOD_CSUM_EN_CFG_D1_IPV4_EN[0:0], MOD_CSUM_EN_CFG.D1_IPV4_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D2_IPV4_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D2_IPV4_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D2_IPV4_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D2_IPV4_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D2_IPV4_EN = write_data[2:2];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D2_IPV4_EN[0], nxt_MOD_CSUM_EN_CFG_D2_IPV4_EN[0:0], MOD_CSUM_EN_CFG.D2_IPV4_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D0_IPV6_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D0_IPV6_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D0_IPV6_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D0_IPV6_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D0_IPV6_EN = write_data[3:3];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D0_IPV6_EN[0], nxt_MOD_CSUM_EN_CFG_D0_IPV6_EN[0:0], MOD_CSUM_EN_CFG.D0_IPV6_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D1_IPV6_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D1_IPV6_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D1_IPV6_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D1_IPV6_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D1_IPV6_EN = write_data[4:4];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D1_IPV6_EN[0], nxt_MOD_CSUM_EN_CFG_D1_IPV6_EN[0:0], MOD_CSUM_EN_CFG.D1_IPV6_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D2_IPV6_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D2_IPV6_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D2_IPV6_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D2_IPV6_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D2_IPV6_EN = write_data[5:5];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D2_IPV6_EN[0], nxt_MOD_CSUM_EN_CFG_D2_IPV6_EN[0:0], MOD_CSUM_EN_CFG.D2_IPV6_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D0_UDP_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D0_UDP_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D0_UDP_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D0_UDP_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D0_UDP_EN = write_data[6:6];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D0_UDP_EN[0], nxt_MOD_CSUM_EN_CFG_D0_UDP_EN[0:0], MOD_CSUM_EN_CFG.D0_UDP_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D1_UDP_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D1_UDP_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D1_UDP_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[0:0]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D1_UDP_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D1_UDP_EN = write_data[7:7];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D1_UDP_EN[0], nxt_MOD_CSUM_EN_CFG_D1_UDP_EN[0:0], MOD_CSUM_EN_CFG.D1_UDP_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D0_TCP_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D0_TCP_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D0_TCP_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[1:1]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D0_TCP_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D0_TCP_EN = write_data[8:8];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D0_TCP_EN[0], nxt_MOD_CSUM_EN_CFG_D0_TCP_EN[0:0], MOD_CSUM_EN_CFG.D0_TCP_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.D1_TCP_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_D1_TCP_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_D1_TCP_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[1:1]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_D1_TCP_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_D1_TCP_EN = write_data[9:9];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_D1_TCP_EN[0], nxt_MOD_CSUM_EN_CFG_D1_TCP_EN[0:0], MOD_CSUM_EN_CFG.D1_TCP_EN[0:0])

// ----------------------------------------------------------------------
// MOD_CSUM_EN_CFG.SCTP_EN x1 RW, using RW template.
logic [0:0] up_MOD_CSUM_EN_CFG_SCTP_EN;
always_comb begin
 up_MOD_CSUM_EN_CFG_SCTP_EN =
    ({1{write_req_MOD_CSUM_EN_CFG }} &
    be[1:1]);
end

logic [0:0] nxt_MOD_CSUM_EN_CFG_SCTP_EN;
always_comb begin
 nxt_MOD_CSUM_EN_CFG_SCTP_EN = write_data[10:10];

end


`RTLGEN_MBY_PPE_MODIFY_MAP_EN_FF(gated_clk, rst_n, 1'h1, up_MOD_CSUM_EN_CFG_SCTP_EN[0], nxt_MOD_CSUM_EN_CFG_SCTP_EN[0:0], MOD_CSUM_EN_CFG.SCTP_EN[0:0])

// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_MODIFY_MAP_MEM) 
           {36'b0?,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_PROFILE_COMMAND;
                    ack.read_miss = handcode_error_MOD_PROFILE_COMMAND;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h2??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_PROFILE_FIELD;
                    ack.read_miss = handcode_error_MOD_PROFILE_FIELD;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_MAP_DUAL;
                    ack.read_miss = handcode_error_MOD_MAP_DUAL;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h2,4'b00??,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_MAP;
                    ack.read_miss = handcode_error_MOD_MAP;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h24,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_PROFILE_GROUP;
                    ack.read_miss = handcode_error_MOD_PROFILE_GROUP;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h24,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_MIRROR_PROFILE_TABLE0;
                    ack.read_miss = handcode_error_MOD_MIRROR_PROFILE_TABLE0;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h24,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_MIRROR_PROFILE_TABLE1;
                    ack.read_miss = handcode_error_MOD_MIRROR_PROFILE_TABLE1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h24,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_MIRROR_PROFILE_TABLE2;
                    ack.read_miss = handcode_error_MOD_MIRROR_PROFILE_TABLE2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {40'h248,4'b000?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_MAP_CFG;
                    ack.read_miss = handcode_error_MOD_MAP_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h2482,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_MAP_DUAL_CFG;
                    ack.read_miss = handcode_error_MOD_MAP_DUAL_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h2482,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_CSUM_CFG1;
                    ack.read_miss = handcode_error_MOD_CSUM_CFG1;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {44'h2483,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_MOD_CSUM_CFG2;
                    ack.read_miss = handcode_error_MOD_CSUM_CFG2;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           MOD_CSUM_EN_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_MODIFY_MAP_MEM) 
           {36'b0?,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_PROFILE_COMMAND;
                    ack.write_miss = handcode_error_MOD_PROFILE_COMMAND;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h2??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_PROFILE_FIELD;
                    ack.write_miss = handcode_error_MOD_PROFILE_FIELD;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_MAP_DUAL;
                    ack.write_miss = handcode_error_MOD_MAP_DUAL;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h2,4'b00??,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_MAP;
                    ack.write_miss = handcode_error_MOD_MAP;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h24,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_PROFILE_GROUP;
                    ack.write_miss = handcode_error_MOD_PROFILE_GROUP;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h24,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_MIRROR_PROFILE_TABLE0;
                    ack.write_miss = handcode_error_MOD_MIRROR_PROFILE_TABLE0;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h24,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_MIRROR_PROFILE_TABLE1;
                    ack.write_miss = handcode_error_MOD_MIRROR_PROFILE_TABLE1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h24,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_MIRROR_PROFILE_TABLE2;
                    ack.write_miss = handcode_error_MOD_MIRROR_PROFILE_TABLE2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {40'h248,4'b000?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_MAP_CFG;
                    ack.write_miss = handcode_error_MOD_MAP_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h2482,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_MAP_DUAL_CFG;
                    ack.write_miss = handcode_error_MOD_MAP_DUAL_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h2482,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_CSUM_CFG1;
                    ack.write_miss = handcode_error_MOD_CSUM_CFG1;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {44'h2483,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_MOD_CSUM_CFG2;
                    ack.write_miss = handcode_error_MOD_CSUM_CFG2;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           MOD_CSUM_EN_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_MODIFY_MAP_MEM) 
           {36'b0?,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_PROFILE_COMMAND;
                 default: read_data = '0;
              endcase
           end
           {44'h2??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_PROFILE_FIELD;
                 default: read_data = '0;
              endcase
           end
           {44'h1???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_MAP_DUAL;
                 default: read_data = '0;
              endcase
           end
           {32'h2,4'b00??,8'h??,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_MAP;
                 default: read_data = '0;
              endcase
           end
           {36'h24,4'b000?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_PROFILE_GROUP;
                 default: read_data = '0;
              endcase
           end
           {36'h24,4'b001?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE0;
                 default: read_data = '0;
              endcase
           end
           {36'h24,4'b010?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE1;
                 default: read_data = '0;
              endcase
           end
           {36'h24,4'b011?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_MIRROR_PROFILE_TABLE2;
                 default: read_data = '0;
              endcase
           end
           {40'h248,4'b000?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_MAP_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'h2482,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_MAP_DUAL_CFG;
                 default: read_data = '0;
              endcase
           end
           {44'h2482,1'b1}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_CSUM_CFG1;
                 default: read_data = '0;
              endcase
           end
           {44'h2483,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = handcode_reg_rdata_MOD_CSUM_CFG2;
                 default: read_data = '0;
              endcase
           end
           MOD_CSUM_EN_CFG_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {MODIFY_SB_FID,MODIFY_SB_BAR}: read_data = {MOD_CSUM_EN_CFG};
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    MOD_CSUM_EN_CFG.reserved0 = '0;
end

// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
