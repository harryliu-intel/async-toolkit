magic
tech scmos
timestamp 969760391
<< ndiffusion >>
rect -50 33 -42 34
rect -20 33 -12 34
rect -50 25 -42 30
rect -20 25 -12 30
rect -50 21 -42 22
rect -50 12 -42 13
rect -50 4 -42 9
rect -20 21 -12 22
rect -20 12 -12 13
rect 67 16 75 17
rect -20 4 -12 9
rect 67 12 75 13
rect 67 3 75 4
rect -50 0 -42 1
rect -20 0 -12 1
rect 67 -1 75 0
<< pdiffusion >>
rect 4 33 12 34
rect 33 33 45 34
rect 4 25 12 30
rect 4 21 12 22
rect 4 12 12 13
rect 33 25 45 30
rect 33 21 45 22
rect 33 12 45 13
rect 91 16 99 17
rect 4 4 12 9
rect 33 4 45 9
rect 91 12 99 13
rect 91 3 99 4
rect 4 0 12 1
rect 33 0 45 1
rect 91 -1 99 0
<< ntransistor >>
rect -50 30 -42 33
rect -20 30 -12 33
rect -50 22 -42 25
rect -20 22 -12 25
rect -50 9 -42 12
rect -20 9 -12 12
rect 67 13 75 16
rect -50 1 -42 4
rect -20 1 -12 4
rect 67 0 75 3
<< ptransistor >>
rect 4 30 12 33
rect 33 30 45 33
rect 4 22 12 25
rect 33 22 45 25
rect 4 9 12 12
rect 33 9 45 12
rect 91 13 99 16
rect 4 1 12 4
rect 33 1 45 4
rect 91 0 99 3
<< polysilicon >>
rect -54 30 -50 33
rect -42 30 -20 33
rect -12 30 4 33
rect 12 30 33 33
rect 45 30 49 33
rect -55 22 -50 25
rect -42 22 -37 25
rect -32 22 -20 25
rect -12 22 4 25
rect 12 22 16 25
rect -55 17 -52 22
rect -54 12 -52 17
rect -54 9 -50 12
rect -42 9 -37 12
rect -32 4 -29 22
rect 21 12 24 30
rect 29 22 33 25
rect 45 22 50 25
rect 47 17 50 22
rect 47 12 49 17
rect -24 9 -20 12
rect -12 9 4 12
rect 12 9 24 12
rect 29 9 33 12
rect 45 9 49 12
rect 62 13 67 16
rect 75 13 91 16
rect 99 13 104 16
rect -54 1 -50 4
rect -42 1 -20 4
rect -12 1 4 4
rect 12 1 33 4
rect 45 1 49 4
rect 62 3 65 13
rect 101 3 104 13
rect 62 0 67 3
rect 75 0 91 3
rect 99 0 104 3
<< ndcontact >>
rect -50 34 -42 42
rect -20 34 -12 42
rect -50 13 -42 21
rect -20 13 -12 21
rect 67 17 75 25
rect 67 4 75 12
rect -50 -8 -42 0
rect -20 -8 -12 0
rect 67 -9 75 -1
<< pdcontact >>
rect 4 34 12 42
rect 33 34 45 42
rect 4 13 12 21
rect 33 13 45 21
rect 91 17 99 25
rect 91 4 99 12
rect 4 -8 12 0
rect 33 -8 45 0
rect 91 -9 99 -1
<< polycontact >>
rect -62 9 -54 17
rect 49 9 57 17
<< metal1 >>
rect -50 34 -12 42
rect 4 34 45 42
rect -62 9 -54 17
rect -50 13 45 21
rect 67 17 75 25
rect 91 17 99 25
rect 49 9 57 17
rect -59 4 54 9
rect 67 4 99 12
rect -50 -8 -12 0
rect 4 -8 45 0
rect 67 -9 75 -1
rect 91 -9 99 -1
<< labels >>
rlabel metal1 -16 38 -16 38 5 GND!
rlabel metal1 8 38 8 38 5 Vdd!
rlabel metal1 -16 -4 -16 -4 1 GND!
rlabel metal1 8 -4 8 -4 1 Vdd!
rlabel metal1 -46 38 -46 38 5 GND!
rlabel metal1 -46 -4 -46 -4 1 GND!
rlabel polysilicon -51 31 -51 31 3 b
rlabel polysilicon -51 2 -51 2 3 a
rlabel polysilicon 46 3 46 3 7 a
rlabel polysilicon 46 32 46 32 7 b
rlabel metal1 39 38 39 38 5 Vdd!
rlabel metal1 39 -4 39 -4 1 Vdd!
rlabel metal1 -46 17 -46 17 1 _x
rlabel metal1 -16 17 -16 17 1 _x
rlabel metal1 8 17 8 17 1 _x
rlabel metal1 39 17 39 17 1 _x
rlabel metal1 53 13 53 13 1 x
rlabel metal1 -58 13 -58 13 1 x
rlabel ndcontact 71 8 71 8 1 x
rlabel pdcontact 95 8 95 8 1 x
rlabel ndcontact 71 -5 71 -5 1 GND!
rlabel pdcontact 95 -5 95 -5 1 Vdd!
rlabel pdcontact 95 21 95 21 5 Vdd!
rlabel ndcontact 71 21 71 21 5 GND!
rlabel polysilicon 66 14 66 14 1 _x
rlabel polysilicon 66 1 66 1 1 _x
rlabel polysilicon 100 14 100 14 1 _x
rlabel polysilicon 100 1 100 1 1 _x
rlabel space -63 -9 -19 43 7 ^n1
rlabel space 10 -9 58 43 3 ^p1
rlabel space 61 -10 68 26 7 ^n2
rlabel space 98 -10 105 26 3 ^p2
<< end >>
