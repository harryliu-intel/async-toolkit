///
///  INTEL CONFIDENTIAL
///
///  Copyright 2018 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            mby_ppe_cgrp_b_nested_map.sv                               
// Creator:         solson                                                     
// Time:            Wednesday Dec 12, 2018 [10:52:23 am]                       
//                                                                             
// Path:            /tmp/solson/nebulon_run/4706538284_2018-12-12.10:40:08     
// Arguments:       -I                                                         
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/tools/srdl
//                  -sv_no_sai_checks -sverilog -xml -chdr -crif -ovm -input   
//                  mby_top_map.rdl -timeout 60000 -out_dir                    
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby
//                  -rtlgencomp -log_file                                      
//                  /nfs/site/disks/slx_1593/solson/mby/work_root/mby-mby-x0_WW5018a/MockTurnin/target/GenRTL/regflow/mby/nebulon_sv_output.log
//                                                                             
// MRE:             5.2018.2                                                   
// Machine:         scci79110                                                  
// OS:              Linux 3.0.101-108.13.1.14249.0.PTF-default                 
// Nebulon version: d18ww24.4                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2018 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d18ww24.4/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_mby_top_map.vh"
`include "rtlgen_pkg_mby_top_map.vh"
`include "mby_ppe_cgrp_b_nested_map_pkg.vh"

//lintra push -68094


// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_RSTD
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_RSTD


module rtlgen_mby_ppe_cgrp_b_nested_map_en_ff_rstd(rtl_clk_var, rst_n_var, rst_val_var, en_var, d_var, q_var);
parameter DATA_WIDTH=1;
input logic rtl_clk_var, rst_n_var, en_var;
input logic [DATA_WIDTH-1:0] rst_val_var, d_var;
output logic [DATA_WIDTH-1:0] q_var;

   genvar gen_var ; 
   generate 
      if (1) begin : rtlgen_en_ff_rstd
         logic [DATA_WIDTH-1:0] rst_vec, set_vec, d_vec, q_vec; 
         assign rst_vec = !rst_n_var ? ~rst_val_var : '0; 
         assign set_vec = !rst_n_var ? rst_val_var : '0; 
         assign d_vec = d_var; 
         assign q_var = q_vec; 
         for ( gen_var = 0 ; gen_var < DATA_WIDTH; gen_var = gen_var + 1)  
            always_ff @(posedge rtl_clk_var, posedge rst_vec[ gen_var ], posedge set_vec[ gen_var ]) 
               if (rst_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '0; 
               else if (set_vec[ gen_var ]) 
                  q_vec[ gen_var ] <= '1; 
               else if (en_var)  
                  q_vec[ gen_var ] <= d_vec[ gen_var ]; 
      end 
   endgenerate       

endmodule 

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_RSTD
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
rtlgen_mby_ppe_cgrp_b_nested_map_en_ff_rstd #(.DATA_WIDTH($bits(q))) \``d``_en_ff_rstd (.rtl_clk_var(rtl_clk), .rst_n_var(rst_n), .rst_val_var(rst_val), .en_var(en), .d_var(d), .q_var(q));
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_RSTD


`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_SYNCRST

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_FF_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_LOW
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_LOW

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_PH2_FF
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) q <= d;
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_PH2_FF

// Can't be override
`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_LOW_ASSIGN
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_PH2_FF_ASSIGN
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_PH2_FF_ASSIGN(n) \
   `RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_PH2_FF_ASSIGN

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_SYNCRST

`ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH_SYNCRST
`define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_LATCH_BOTHRST
// 
// `ifndef RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH_BOTHRST
// `define RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_LATCH_BOTHRST


//lintra pop

module mby_ppe_cgrp_b_nested_map ( //lintra s-2096
    // Clocks
    gated_clk,
    rtl_clk,

    // Resets
    rst_n,


    // Register Inputs
    load_WCM_IP,

    new_WCM_IP,

    handcode_reg_rdata_EM_HASH_LOOKUP,
    handcode_reg_rdata_IDX,
    handcode_reg_rdata_WCM_ACTION,
    handcode_reg_rdata_WCM_ACTION_CFG_EN,
    handcode_reg_rdata_WCM_TCAM,
    handcode_reg_rdata_WCM_TCAM_CFG,

    handcode_rvalid_EM_HASH_LOOKUP,
    handcode_rvalid_IDX,
    handcode_rvalid_WCM_ACTION,
    handcode_rvalid_WCM_ACTION_CFG_EN,
    handcode_rvalid_WCM_TCAM,
    handcode_rvalid_WCM_TCAM_CFG,

    handcode_wvalid_EM_HASH_LOOKUP,
    handcode_wvalid_IDX,
    handcode_wvalid_WCM_ACTION,
    handcode_wvalid_WCM_ACTION_CFG_EN,
    handcode_wvalid_WCM_TCAM,
    handcode_wvalid_WCM_TCAM_CFG,

    handcode_error_EM_HASH_LOOKUP,
    handcode_error_IDX,
    handcode_error_WCM_ACTION,
    handcode_error_WCM_ACTION_CFG_EN,
    handcode_error_WCM_TCAM,
    handcode_error_WCM_TCAM_CFG,


    // Register Outputs
    WCM_IM,
    WCM_IP,


    // Register signals for HandCoded registers
    handcode_reg_wdata_EM_HASH_LOOKUP,
    handcode_reg_wdata_IDX,
    handcode_reg_wdata_WCM_ACTION,
    handcode_reg_wdata_WCM_ACTION_CFG_EN,
    handcode_reg_wdata_WCM_TCAM,
    handcode_reg_wdata_WCM_TCAM_CFG,

    we_EM_HASH_LOOKUP,
    we_IDX,
    we_WCM_ACTION,
    we_WCM_ACTION_CFG_EN,
    we_WCM_TCAM,
    we_WCM_TCAM_CFG,

    re_EM_HASH_LOOKUP,
    re_IDX,
    re_WCM_ACTION,
    re_WCM_ACTION_CFG_EN,
    re_WCM_TCAM,
    re_WCM_TCAM_CFG,




    // Config Access
    req,
    ack
    

);

import mby_ppe_cgrp_b_nested_map_pkg::*;
import rtlgen_pkg_mby_top_map::*;

parameter  MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB = 47;
parameter [MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:0] MBY_PPE_CGRP_B_NESTED_MAP_OFFSET = {MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB+1{1'b0}};
parameter [2:0] B_SB_BAR = 3'b0;
parameter [7:0] B_SB_FID = 8'b0;
localparam  ADDR_LSB_BUS_ALIGN = 3;
localparam [MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] WCM_IP_DECODE_ADDR = WCM_IP_CR_ADDR[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CGRP_B_NESTED_MAP_OFFSET[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] WCM_IM_DECODE_ADDR = WCM_IM_CR_ADDR[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MBY_PPE_CGRP_B_NESTED_MAP_OFFSET[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];

    // Clocks
input logic  gated_clk;
input logic  rtl_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input load_WCM_IP_t  load_WCM_IP;

input new_WCM_IP_t  new_WCM_IP;

input EM_HASH_LOOKUP_t  handcode_reg_rdata_EM_HASH_LOOKUP;
input IDX_t  handcode_reg_rdata_IDX;
input WCM_ACTION_t  handcode_reg_rdata_WCM_ACTION;
input WCM_ACTION_CFG_EN_t  handcode_reg_rdata_WCM_ACTION_CFG_EN;
input WCM_TCAM_t  handcode_reg_rdata_WCM_TCAM;
input WCM_TCAM_CFG_t  handcode_reg_rdata_WCM_TCAM_CFG;

input handcode_rvalid_EM_HASH_LOOKUP_t  handcode_rvalid_EM_HASH_LOOKUP;
input handcode_rvalid_IDX_t  handcode_rvalid_IDX;
input handcode_rvalid_WCM_ACTION_t  handcode_rvalid_WCM_ACTION;
input handcode_rvalid_WCM_ACTION_CFG_EN_t  handcode_rvalid_WCM_ACTION_CFG_EN;
input handcode_rvalid_WCM_TCAM_t  handcode_rvalid_WCM_TCAM;
input handcode_rvalid_WCM_TCAM_CFG_t  handcode_rvalid_WCM_TCAM_CFG;

input handcode_wvalid_EM_HASH_LOOKUP_t  handcode_wvalid_EM_HASH_LOOKUP;
input handcode_wvalid_IDX_t  handcode_wvalid_IDX;
input handcode_wvalid_WCM_ACTION_t  handcode_wvalid_WCM_ACTION;
input handcode_wvalid_WCM_ACTION_CFG_EN_t  handcode_wvalid_WCM_ACTION_CFG_EN;
input handcode_wvalid_WCM_TCAM_t  handcode_wvalid_WCM_TCAM;
input handcode_wvalid_WCM_TCAM_CFG_t  handcode_wvalid_WCM_TCAM_CFG;

input handcode_error_EM_HASH_LOOKUP_t  handcode_error_EM_HASH_LOOKUP;
input handcode_error_IDX_t  handcode_error_IDX;
input handcode_error_WCM_ACTION_t  handcode_error_WCM_ACTION;
input handcode_error_WCM_ACTION_CFG_EN_t  handcode_error_WCM_ACTION_CFG_EN;
input handcode_error_WCM_TCAM_t  handcode_error_WCM_TCAM;
input handcode_error_WCM_TCAM_CFG_t  handcode_error_WCM_TCAM_CFG;


    // Register Outputs
output WCM_IM_t  WCM_IM;
output WCM_IP_t  WCM_IP;


    // Register signals for HandCoded registers
output EM_HASH_LOOKUP_t  handcode_reg_wdata_EM_HASH_LOOKUP;
output IDX_t  handcode_reg_wdata_IDX;
output WCM_ACTION_t  handcode_reg_wdata_WCM_ACTION;
output WCM_ACTION_CFG_EN_t  handcode_reg_wdata_WCM_ACTION_CFG_EN;
output WCM_TCAM_t  handcode_reg_wdata_WCM_TCAM;
output WCM_TCAM_CFG_t  handcode_reg_wdata_WCM_TCAM_CFG;

output we_EM_HASH_LOOKUP_t  we_EM_HASH_LOOKUP;
output we_IDX_t  we_IDX;
output we_WCM_ACTION_t  we_WCM_ACTION;
output we_WCM_ACTION_CFG_EN_t  we_WCM_ACTION_CFG_EN;
output we_WCM_TCAM_t  we_WCM_TCAM;
output we_WCM_TCAM_CFG_t  we_WCM_TCAM_CFG;

output re_EM_HASH_LOOKUP_t  re_EM_HASH_LOOKUP;
output re_IDX_t  re_IDX;
output re_WCM_ACTION_t  re_WCM_ACTION;
output re_WCM_ACTION_CFG_EN_t  re_WCM_ACTION_CFG_EN;
output re_WCM_TCAM_t  re_WCM_TCAM;
output re_WCM_TCAM_CFG_t  re_WCM_TCAM_CFG;




    // Config Access
input mby_ppe_cgrp_b_nested_map_cr_req_t  req;
output mby_ppe_cgrp_b_nested_map_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input mby_ppe_cgrp_b_nested_map_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;

logic [7:0] req_fid;
assign req_fid = req.fid;
logic [2:0] req_bar;
assign req_bar = req.bar;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_MBY_PPE_CGRP_B_NESTED_MAP_MEM;
assign case_req_addr_MBY_PPE_CGRP_B_NESTED_MAP_MEM = req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;



logic sb_fid_cond_b;
always_comb begin : sb_fid_cond_b_BLOCK
    unique casez (req_fid) 
		B_SB_FID: sb_fid_cond_b = 1;
		default: sb_fid_cond_b = 0;
    endcase 
end


logic sb_bar_cond_b;
always_comb begin : sb_bar_cond_b_BLOCK
    unique casez (req_bar) 
		B_SB_BAR: sb_bar_cond_b = 1;
		default: sb_bar_cond_b = 0;
    endcase 
end


// ======================================================================
// begin register logic section {

// ----------------------------------------------------------------------
// EM_HASH_LOOKUP using HANDCODED_REG template.
logic addr_decode_EM_HASH_LOOKUP;
logic write_req_EM_HASH_LOOKUP;
logic read_req_EM_HASH_LOOKUP;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b0?,12'h???,1'b0}: 
         addr_decode_EM_HASH_LOOKUP = req.valid;
      default: 
         addr_decode_EM_HASH_LOOKUP = 1'b0; 
   endcase
end

always_comb write_req_EM_HASH_LOOKUP = f_IsMEMWr(req_opcode) && addr_decode_EM_HASH_LOOKUP ;
always_comb read_req_EM_HASH_LOOKUP  = f_IsMEMRd(req_opcode) && addr_decode_EM_HASH_LOOKUP ;

always_comb we_EM_HASH_LOOKUP = {16{write_req_EM_HASH_LOOKUP}} & req.be[15:0];
always_comb re_EM_HASH_LOOKUP = {16{read_req_EM_HASH_LOOKUP}} & req.be[15:0];
always_comb handcode_reg_wdata_EM_HASH_LOOKUP = req.data[127:0];


// ----------------------------------------------------------------------
// WCM_TCAM using HANDCODED_REG template.
logic addr_decode_WCM_TCAM;
logic write_req_WCM_TCAM;
logic read_req_WCM_TCAM;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'b10??,12'h???,1'b0},
      {44'hC???,1'b0}:
          addr_decode_WCM_TCAM = req.valid;
      default: 
         addr_decode_WCM_TCAM = 1'b0; 
   endcase
end

always_comb write_req_WCM_TCAM = f_IsMEMWr(req_opcode) && addr_decode_WCM_TCAM ;
always_comb read_req_WCM_TCAM  = f_IsMEMRd(req_opcode) && addr_decode_WCM_TCAM ;

always_comb we_WCM_TCAM = {16{write_req_WCM_TCAM}} & req.be[15:0];
always_comb re_WCM_TCAM = {16{read_req_WCM_TCAM}} & req.be[15:0];
always_comb handcode_reg_wdata_WCM_TCAM = req.data[127:0];


// ----------------------------------------------------------------------
// WCM_ACTION using HANDCODED_REG template.
logic addr_decode_WCM_ACTION;
logic write_req_WCM_ACTION;
logic read_req_WCM_ACTION;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {28'h1,4'b000?,12'h???,1'b?},
      {44'h12???,1'b?}:
          addr_decode_WCM_ACTION = req.valid;
      default: 
         addr_decode_WCM_ACTION = 1'b0; 
   endcase
end

always_comb write_req_WCM_ACTION = f_IsMEMWr(req_opcode) && addr_decode_WCM_ACTION ;
always_comb read_req_WCM_ACTION  = f_IsMEMRd(req_opcode) && addr_decode_WCM_ACTION ;

always_comb we_WCM_ACTION = {8{write_req_WCM_ACTION}} & be;
always_comb re_WCM_ACTION = {8{read_req_WCM_ACTION}} & be;
always_comb handcode_reg_wdata_WCM_ACTION = write_data;


// ----------------------------------------------------------------------
// WCM_TCAM_CFG using HANDCODED_REG template.
logic addr_decode_WCM_TCAM_CFG;
logic write_req_WCM_TCAM_CFG;
logic read_req_WCM_TCAM_CFG;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {32'h13,4'b000?,8'h??,1'b?},
      {36'h132,4'b0???,4'h?,1'b?}:
          addr_decode_WCM_TCAM_CFG = req.valid;
      default: 
         addr_decode_WCM_TCAM_CFG = 1'b0; 
   endcase
end

always_comb write_req_WCM_TCAM_CFG = f_IsMEMWr(req_opcode) && addr_decode_WCM_TCAM_CFG ;
always_comb read_req_WCM_TCAM_CFG  = f_IsMEMRd(req_opcode) && addr_decode_WCM_TCAM_CFG ;

always_comb we_WCM_TCAM_CFG = {8{write_req_WCM_TCAM_CFG}} & be;
always_comb re_WCM_TCAM_CFG = {8{read_req_WCM_TCAM_CFG}} & be;
always_comb handcode_reg_wdata_WCM_TCAM_CFG = write_data;


// ----------------------------------------------------------------------
// WCM_ACTION_CFG_EN using HANDCODED_REG template.
logic addr_decode_WCM_ACTION_CFG_EN;
logic write_req_WCM_ACTION_CFG_EN;
logic read_req_WCM_ACTION_CFG_EN;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h132,4'b100?,4'h?,1'b?}: 
         addr_decode_WCM_ACTION_CFG_EN = req.valid;
      default: 
         addr_decode_WCM_ACTION_CFG_EN = 1'b0; 
   endcase
end

always_comb write_req_WCM_ACTION_CFG_EN = f_IsMEMWr(req_opcode) && addr_decode_WCM_ACTION_CFG_EN ;
always_comb read_req_WCM_ACTION_CFG_EN  = f_IsMEMRd(req_opcode) && addr_decode_WCM_ACTION_CFG_EN ;

always_comb we_WCM_ACTION_CFG_EN = {8{write_req_WCM_ACTION_CFG_EN}} & be;
always_comb re_WCM_ACTION_CFG_EN = {8{read_req_WCM_ACTION_CFG_EN}} & be;
always_comb handcode_reg_wdata_WCM_ACTION_CFG_EN = write_data;


// ----------------------------------------------------------------------
// IDX using HANDCODED_REG template.
logic addr_decode_IDX;
logic write_req_IDX;
logic read_req_IDX;

always_comb begin 
   unique casez (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN]) 
      {36'h132,4'b11??,4'h?,1'b?}: 
         addr_decode_IDX = req.valid;
      default: 
         addr_decode_IDX = 1'b0; 
   endcase
end

always_comb write_req_IDX = f_IsMEMWr(req_opcode) && addr_decode_IDX ;
always_comb read_req_IDX  = f_IsMEMRd(req_opcode) && addr_decode_IDX ;

always_comb we_IDX = {8{write_req_IDX}} & be;
always_comb re_IDX = {8{read_req_IDX}} & be;
always_comb handcode_reg_wdata_IDX = write_data;


//---------------------------------------------------------------------
// WCM_IP Address Decode
logic  addr_decode_WCM_IP;
logic  write_req_WCM_IP;
always_comb begin
   addr_decode_WCM_IP = (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == WCM_IP_DECODE_ADDR) && req.valid ;
   write_req_WCM_IP = IsMEMWr && addr_decode_WCM_IP && sb_fid_cond_b && sb_bar_cond_b;
end

// ----------------------------------------------------------------------
// WCM_IP.FCMN_SHELL_CTRL_ERR x1 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [0:0] req_up_WCM_IP_FCMN_SHELL_CTRL_ERR;
always_comb begin
 req_up_WCM_IP_FCMN_SHELL_CTRL_ERR[0:0] = 
   {1{write_req_WCM_IP & be[0]}}
;
end

logic [0:0] clr_WCM_IP_FCMN_SHELL_CTRL_ERR;
always_comb begin
 clr_WCM_IP_FCMN_SHELL_CTRL_ERR = write_data[0:0] & req_up_WCM_IP_FCMN_SHELL_CTRL_ERR;

end
logic [0:0] swwr_WCM_IP_FCMN_SHELL_CTRL_ERR;
logic [0:0] sw_nxt_WCM_IP_FCMN_SHELL_CTRL_ERR;
always_comb begin
 swwr_WCM_IP_FCMN_SHELL_CTRL_ERR = clr_WCM_IP_FCMN_SHELL_CTRL_ERR;
 sw_nxt_WCM_IP_FCMN_SHELL_CTRL_ERR = {1{1'b0}};

end
logic [0:0] up_WCM_IP_FCMN_SHELL_CTRL_ERR;
logic [0:0] nxt_WCM_IP_FCMN_SHELL_CTRL_ERR;
always_comb begin
 up_WCM_IP_FCMN_SHELL_CTRL_ERR = 
   swwr_WCM_IP_FCMN_SHELL_CTRL_ERR | {1{load_WCM_IP.FCMN_SHELL_CTRL_ERR}};
end
always_comb begin
 nxt_WCM_IP_FCMN_SHELL_CTRL_ERR[0] = 
    load_WCM_IP.FCMN_SHELL_CTRL_ERR ?
    new_WCM_IP.FCMN_SHELL_CTRL_ERR[0] :
    sw_nxt_WCM_IP_FCMN_SHELL_CTRL_ERR[0];
end



`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_FCMN_SHELL_CTRL_ERR[0], nxt_WCM_IP_FCMN_SHELL_CTRL_ERR[0], WCM_IP.FCMN_SHELL_CTRL_ERR[0])

// ----------------------------------------------------------------------
// WCM_IP.TCAM_SWEEP_ERR x1 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [0:0] req_up_WCM_IP_TCAM_SWEEP_ERR;
always_comb begin
 req_up_WCM_IP_TCAM_SWEEP_ERR[0:0] = 
   {1{write_req_WCM_IP & be[0]}}
;
end

logic [0:0] clr_WCM_IP_TCAM_SWEEP_ERR;
always_comb begin
 clr_WCM_IP_TCAM_SWEEP_ERR = write_data[1:1] & req_up_WCM_IP_TCAM_SWEEP_ERR;

end
logic [0:0] swwr_WCM_IP_TCAM_SWEEP_ERR;
logic [0:0] sw_nxt_WCM_IP_TCAM_SWEEP_ERR;
always_comb begin
 swwr_WCM_IP_TCAM_SWEEP_ERR = clr_WCM_IP_TCAM_SWEEP_ERR;
 sw_nxt_WCM_IP_TCAM_SWEEP_ERR = {1{1'b0}};

end
logic [0:0] up_WCM_IP_TCAM_SWEEP_ERR;
logic [0:0] nxt_WCM_IP_TCAM_SWEEP_ERR;
always_comb begin
 up_WCM_IP_TCAM_SWEEP_ERR = 
   swwr_WCM_IP_TCAM_SWEEP_ERR | {1{load_WCM_IP.TCAM_SWEEP_ERR}};
end
always_comb begin
 nxt_WCM_IP_TCAM_SWEEP_ERR[0] = 
    load_WCM_IP.TCAM_SWEEP_ERR ?
    new_WCM_IP.TCAM_SWEEP_ERR[0] :
    sw_nxt_WCM_IP_TCAM_SWEEP_ERR[0];
end



`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_TCAM_SWEEP_ERR[0], nxt_WCM_IP_TCAM_SWEEP_ERR[0], WCM_IP.TCAM_SWEEP_ERR[0])

// ----------------------------------------------------------------------
// WCM_IP.FGRP_ERR x3 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [2:0] req_up_WCM_IP_FGRP_ERR;
always_comb begin
 req_up_WCM_IP_FGRP_ERR[2:0] = 
   {3{write_req_WCM_IP & be[0]}}
;
end

logic [2:0] clr_WCM_IP_FGRP_ERR;
always_comb begin
 clr_WCM_IP_FGRP_ERR = write_data[4:2] & req_up_WCM_IP_FGRP_ERR;

end
logic [2:0] swwr_WCM_IP_FGRP_ERR;
logic [2:0] sw_nxt_WCM_IP_FGRP_ERR;
always_comb begin
 swwr_WCM_IP_FGRP_ERR = clr_WCM_IP_FGRP_ERR;
 sw_nxt_WCM_IP_FGRP_ERR = {3{1'b0}};

end
logic [2:0] up_WCM_IP_FGRP_ERR;
logic [2:0] nxt_WCM_IP_FGRP_ERR;
always_comb begin
 up_WCM_IP_FGRP_ERR = 
   swwr_WCM_IP_FGRP_ERR | {3{load_WCM_IP.FGRP_ERR}};
end
always_comb begin
 nxt_WCM_IP_FGRP_ERR[0] = 
    load_WCM_IP.FGRP_ERR ?
    new_WCM_IP.FGRP_ERR[0] :
    sw_nxt_WCM_IP_FGRP_ERR[0];
 nxt_WCM_IP_FGRP_ERR[1] = 
    load_WCM_IP.FGRP_ERR ?
    new_WCM_IP.FGRP_ERR[1] :
    sw_nxt_WCM_IP_FGRP_ERR[1];
 nxt_WCM_IP_FGRP_ERR[2] = 
    load_WCM_IP.FGRP_ERR ?
    new_WCM_IP.FGRP_ERR[2] :
    sw_nxt_WCM_IP_FGRP_ERR[2];
end



`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_FGRP_ERR[0], nxt_WCM_IP_FGRP_ERR[0], WCM_IP.FGRP_ERR[0])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_FGRP_ERR[1], nxt_WCM_IP_FGRP_ERR[1], WCM_IP.FGRP_ERR[1])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_FGRP_ERR[2], nxt_WCM_IP_FGRP_ERR[2], WCM_IP.FGRP_ERR[2])

// ----------------------------------------------------------------------
// WCM_IP.FGHASH_ERR x3 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [2:0] req_up_WCM_IP_FGHASH_ERR;
always_comb begin
 req_up_WCM_IP_FGHASH_ERR[2:0] = 
   {3{write_req_WCM_IP & be[0]}}
;
end

logic [2:0] clr_WCM_IP_FGHASH_ERR;
always_comb begin
 clr_WCM_IP_FGHASH_ERR = write_data[7:5] & req_up_WCM_IP_FGHASH_ERR;

end
logic [2:0] swwr_WCM_IP_FGHASH_ERR;
logic [2:0] sw_nxt_WCM_IP_FGHASH_ERR;
always_comb begin
 swwr_WCM_IP_FGHASH_ERR = clr_WCM_IP_FGHASH_ERR;
 sw_nxt_WCM_IP_FGHASH_ERR = {3{1'b0}};

end
logic [2:0] up_WCM_IP_FGHASH_ERR;
logic [2:0] nxt_WCM_IP_FGHASH_ERR;
always_comb begin
 up_WCM_IP_FGHASH_ERR = 
   swwr_WCM_IP_FGHASH_ERR | {3{load_WCM_IP.FGHASH_ERR}};
end
always_comb begin
 nxt_WCM_IP_FGHASH_ERR[0] = 
    load_WCM_IP.FGHASH_ERR ?
    new_WCM_IP.FGHASH_ERR[0] :
    sw_nxt_WCM_IP_FGHASH_ERR[0];
 nxt_WCM_IP_FGHASH_ERR[1] = 
    load_WCM_IP.FGHASH_ERR ?
    new_WCM_IP.FGHASH_ERR[1] :
    sw_nxt_WCM_IP_FGHASH_ERR[1];
 nxt_WCM_IP_FGHASH_ERR[2] = 
    load_WCM_IP.FGHASH_ERR ?
    new_WCM_IP.FGHASH_ERR[2] :
    sw_nxt_WCM_IP_FGHASH_ERR[2];
end



`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_FGHASH_ERR[0], nxt_WCM_IP_FGHASH_ERR[0], WCM_IP.FGHASH_ERR[0])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_FGHASH_ERR[1], nxt_WCM_IP_FGHASH_ERR[1], WCM_IP.FGHASH_ERR[1])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_FGHASH_ERR[2], nxt_WCM_IP_FGHASH_ERR[2], WCM_IP.FGHASH_ERR[2])

// ----------------------------------------------------------------------
// WCM_IP.HASH_ENTRY_RAM_U_ERR x4 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [3:0] req_up_WCM_IP_HASH_ENTRY_RAM_U_ERR;
always_comb begin
 req_up_WCM_IP_HASH_ENTRY_RAM_U_ERR[3:0] = 
   {4{write_req_WCM_IP & be[1]}}
;
end

logic [3:0] clr_WCM_IP_HASH_ENTRY_RAM_U_ERR;
always_comb begin
 clr_WCM_IP_HASH_ENTRY_RAM_U_ERR = write_data[11:8] & req_up_WCM_IP_HASH_ENTRY_RAM_U_ERR;

end
logic [3:0] swwr_WCM_IP_HASH_ENTRY_RAM_U_ERR;
logic [3:0] sw_nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR;
always_comb begin
 swwr_WCM_IP_HASH_ENTRY_RAM_U_ERR = clr_WCM_IP_HASH_ENTRY_RAM_U_ERR;
 sw_nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR = {4{1'b0}};

end
logic [3:0] up_WCM_IP_HASH_ENTRY_RAM_U_ERR;
logic [3:0] nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR;
always_comb begin
 up_WCM_IP_HASH_ENTRY_RAM_U_ERR = 
   swwr_WCM_IP_HASH_ENTRY_RAM_U_ERR | {4{load_WCM_IP.HASH_ENTRY_RAM_U_ERR}};
end
always_comb begin
 nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[0] = 
    load_WCM_IP.HASH_ENTRY_RAM_U_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_U_ERR[0] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[0];
 nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[1] = 
    load_WCM_IP.HASH_ENTRY_RAM_U_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_U_ERR[1] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[1];
 nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[2] = 
    load_WCM_IP.HASH_ENTRY_RAM_U_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_U_ERR[2] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[2];
 nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[3] = 
    load_WCM_IP.HASH_ENTRY_RAM_U_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_U_ERR[3] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[3];
end



`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_U_ERR[0], nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[0], WCM_IP.HASH_ENTRY_RAM_U_ERR[0])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_U_ERR[1], nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[1], WCM_IP.HASH_ENTRY_RAM_U_ERR[1])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_U_ERR[2], nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[2], WCM_IP.HASH_ENTRY_RAM_U_ERR[2])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_U_ERR[3], nxt_WCM_IP_HASH_ENTRY_RAM_U_ERR[3], WCM_IP.HASH_ENTRY_RAM_U_ERR[3])

// ----------------------------------------------------------------------
// WCM_IP.HASH_ENTRY_RAM_C_ERR x4 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [3:0] req_up_WCM_IP_HASH_ENTRY_RAM_C_ERR;
always_comb begin
 req_up_WCM_IP_HASH_ENTRY_RAM_C_ERR[3:0] = 
   {4{write_req_WCM_IP & be[1]}}
;
end

logic [3:0] clr_WCM_IP_HASH_ENTRY_RAM_C_ERR;
always_comb begin
 clr_WCM_IP_HASH_ENTRY_RAM_C_ERR = write_data[15:12] & req_up_WCM_IP_HASH_ENTRY_RAM_C_ERR;

end
logic [3:0] swwr_WCM_IP_HASH_ENTRY_RAM_C_ERR;
logic [3:0] sw_nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR;
always_comb begin
 swwr_WCM_IP_HASH_ENTRY_RAM_C_ERR = clr_WCM_IP_HASH_ENTRY_RAM_C_ERR;
 sw_nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR = {4{1'b0}};

end
logic [3:0] up_WCM_IP_HASH_ENTRY_RAM_C_ERR;
logic [3:0] nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR;
always_comb begin
 up_WCM_IP_HASH_ENTRY_RAM_C_ERR = 
   swwr_WCM_IP_HASH_ENTRY_RAM_C_ERR | {4{load_WCM_IP.HASH_ENTRY_RAM_C_ERR}};
end
always_comb begin
 nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[0] = 
    load_WCM_IP.HASH_ENTRY_RAM_C_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_C_ERR[0] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[0];
 nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[1] = 
    load_WCM_IP.HASH_ENTRY_RAM_C_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_C_ERR[1] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[1];
 nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[2] = 
    load_WCM_IP.HASH_ENTRY_RAM_C_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_C_ERR[2] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[2];
 nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[3] = 
    load_WCM_IP.HASH_ENTRY_RAM_C_ERR ?
    new_WCM_IP.HASH_ENTRY_RAM_C_ERR[3] :
    sw_nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[3];
end



`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_C_ERR[0], nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[0], WCM_IP.HASH_ENTRY_RAM_C_ERR[0])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_C_ERR[1], nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[1], WCM_IP.HASH_ENTRY_RAM_C_ERR[1])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_C_ERR[2], nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[2], WCM_IP.HASH_ENTRY_RAM_C_ERR[2])
`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(rtl_clk, rst_n, 1'h0, up_WCM_IP_HASH_ENTRY_RAM_C_ERR[3], nxt_WCM_IP_HASH_ENTRY_RAM_C_ERR[3], WCM_IP.HASH_ENTRY_RAM_C_ERR[3])

//---------------------------------------------------------------------
// WCM_IM Address Decode
logic  addr_decode_WCM_IM;
logic  write_req_WCM_IM;
always_comb begin
   addr_decode_WCM_IM = (req_addr[MBY_PPE_CGRP_B_NESTED_MAP_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == WCM_IM_DECODE_ADDR) && req.valid ;
   write_req_WCM_IM = IsMEMWr && addr_decode_WCM_IM && sb_fid_cond_b && sb_bar_cond_b;
end

// ----------------------------------------------------------------------
// WCM_IM.FCMN_SHELL_CTRL_ERR x1 RW, using RW template.
logic [0:0] up_WCM_IM_FCMN_SHELL_CTRL_ERR;
always_comb begin
 up_WCM_IM_FCMN_SHELL_CTRL_ERR =
    ({1{write_req_WCM_IM }} &
    be[0:0]);
end

logic [0:0] nxt_WCM_IM_FCMN_SHELL_CTRL_ERR;
always_comb begin
 nxt_WCM_IM_FCMN_SHELL_CTRL_ERR = write_data[0:0];

end


`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_WCM_IM_FCMN_SHELL_CTRL_ERR[0], nxt_WCM_IM_FCMN_SHELL_CTRL_ERR[0:0], WCM_IM.FCMN_SHELL_CTRL_ERR[0:0])

// ----------------------------------------------------------------------
// WCM_IM.TCAM_SWEEP_ERR x1 RW, using RW template.
logic [0:0] up_WCM_IM_TCAM_SWEEP_ERR;
always_comb begin
 up_WCM_IM_TCAM_SWEEP_ERR =
    ({1{write_req_WCM_IM }} &
    be[0:0]);
end

logic [0:0] nxt_WCM_IM_TCAM_SWEEP_ERR;
always_comb begin
 nxt_WCM_IM_TCAM_SWEEP_ERR = write_data[1:1];

end


`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(gated_clk, rst_n, 1'h0, up_WCM_IM_TCAM_SWEEP_ERR[0], nxt_WCM_IM_TCAM_SWEEP_ERR[0:0], WCM_IM.TCAM_SWEEP_ERR[0:0])

// ----------------------------------------------------------------------
// WCM_IM.FGRP_ERR x3 RW, using RW template.
logic [0:0] up_WCM_IM_FGRP_ERR;
always_comb begin
 up_WCM_IM_FGRP_ERR =
    ({1{write_req_WCM_IM }} &
    be[0:0]);
end

logic [2:0] nxt_WCM_IM_FGRP_ERR;
always_comb begin
 nxt_WCM_IM_FGRP_ERR = write_data[4:2];

end


`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(gated_clk, rst_n, 3'h0, up_WCM_IM_FGRP_ERR[0], nxt_WCM_IM_FGRP_ERR[2:0], WCM_IM.FGRP_ERR[2:0])

// ----------------------------------------------------------------------
// WCM_IM.FGHASH_ERR x3 RW, using RW template.
logic [0:0] up_WCM_IM_FGHASH_ERR;
always_comb begin
 up_WCM_IM_FGHASH_ERR =
    ({1{write_req_WCM_IM }} &
    be[0:0]);
end

logic [2:0] nxt_WCM_IM_FGHASH_ERR;
always_comb begin
 nxt_WCM_IM_FGHASH_ERR = write_data[7:5];

end


`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(gated_clk, rst_n, 3'h0, up_WCM_IM_FGHASH_ERR[0], nxt_WCM_IM_FGHASH_ERR[2:0], WCM_IM.FGHASH_ERR[2:0])

// ----------------------------------------------------------------------
// WCM_IM.HASH_ENTRY_RAM_U_ERR x4 RW, using RW template.
logic [0:0] up_WCM_IM_HASH_ENTRY_RAM_U_ERR;
always_comb begin
 up_WCM_IM_HASH_ENTRY_RAM_U_ERR =
    ({1{write_req_WCM_IM }} &
    be[1:1]);
end

logic [3:0] nxt_WCM_IM_HASH_ENTRY_RAM_U_ERR;
always_comb begin
 nxt_WCM_IM_HASH_ENTRY_RAM_U_ERR = write_data[11:8];

end


`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(gated_clk, rst_n, 4'h0, up_WCM_IM_HASH_ENTRY_RAM_U_ERR[0], nxt_WCM_IM_HASH_ENTRY_RAM_U_ERR[3:0], WCM_IM.HASH_ENTRY_RAM_U_ERR[3:0])

// ----------------------------------------------------------------------
// WCM_IM.HASH_ENTRY_RAM_C_ERR x4 RW, using RW template.
logic [0:0] up_WCM_IM_HASH_ENTRY_RAM_C_ERR;
always_comb begin
 up_WCM_IM_HASH_ENTRY_RAM_C_ERR =
    ({1{write_req_WCM_IM }} &
    be[1:1]);
end

logic [3:0] nxt_WCM_IM_HASH_ENTRY_RAM_C_ERR;
always_comb begin
 nxt_WCM_IM_HASH_ENTRY_RAM_C_ERR = write_data[15:12];

end


`RTLGEN_MBY_PPE_CGRP_B_NESTED_MAP_EN_FF(gated_clk, rst_n, 4'h0, up_WCM_IM_HASH_ENTRY_RAM_C_ERR[0], nxt_WCM_IM_HASH_ENTRY_RAM_C_ERR[3:0], WCM_IM.HASH_ENTRY_RAM_C_ERR[3:0])

// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_MBY_PPE_CGRP_B_NESTED_MAP_MEM) 
           {32'b0?,12'h???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_EM_HASH_LOOKUP;
                    ack.read_miss = handcode_error_EM_HASH_LOOKUP;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'b10??,12'h???,1'b0},
           {44'hC???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_WCM_TCAM;
                    ack.read_miss = handcode_error_WCM_TCAM;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {28'h1,4'b000?,12'h???,1'b?},
           {44'h12???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_WCM_ACTION;
                    ack.read_miss = handcode_error_WCM_ACTION;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {32'h13,4'b000?,8'h??,1'b?},
           {36'h132,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_WCM_TCAM_CFG;
                    ack.read_miss = handcode_error_WCM_TCAM_CFG;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h132,4'b100?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_WCM_ACTION_CFG_EN;
                    ack.read_miss = handcode_error_WCM_ACTION_CFG_EN;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           {36'h132,4'b11??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.read_valid = req.valid && handcode_rvalid_IDX;
                    ack.read_miss = handcode_error_IDX;
                 end
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           WCM_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
           WCM_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: ack.read_miss = 1'b0;
                 default: ack.read_miss = ack.read_valid;
              endcase
           end
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_MBY_PPE_CGRP_B_NESTED_MAP_MEM) 
           {32'b0?,12'h???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_EM_HASH_LOOKUP;
                    ack.write_miss = handcode_error_EM_HASH_LOOKUP;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'b10??,12'h???,1'b0},
           {44'hC???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_WCM_TCAM;
                    ack.write_miss = handcode_error_WCM_TCAM;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {28'h1,4'b000?,12'h???,1'b?},
           {44'h12???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_WCM_ACTION;
                    ack.write_miss = handcode_error_WCM_ACTION;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {32'h13,4'b000?,8'h??,1'b?},
           {36'h132,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_WCM_TCAM_CFG;
                    ack.write_miss = handcode_error_WCM_TCAM_CFG;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h132,4'b100?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_WCM_ACTION_CFG_EN;
                    ack.write_miss = handcode_error_WCM_ACTION_CFG_EN;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           {36'h132,4'b11??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: begin
                    ack.write_valid = req.valid && handcode_wvalid_IDX;
                    ack.write_miss = handcode_error_IDX;
                 end
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           WCM_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
           WCM_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: ack.write_miss = 1'b0;
                 default: ack.write_miss = ack.write_valid;
              endcase
           end
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

assign sai_successfull_per_byte = {8{1'b1}};

always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      MRD:
         unique casez (case_req_addr_MBY_PPE_CGRP_B_NESTED_MAP_MEM) 
           {32'b0?,12'h???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = handcode_reg_rdata_EM_HASH_LOOKUP;
                 default: read_data = '0;
              endcase
           end
           {32'b10??,12'h???,1'b0},
           {44'hC???,1'b0}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = handcode_reg_rdata_WCM_TCAM;
                 default: read_data = '0;
              endcase
           end
           {28'h1,4'b000?,12'h???,1'b?},
           {44'h12???,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = handcode_reg_rdata_WCM_ACTION;
                 default: read_data = '0;
              endcase
           end
           {32'h13,4'b000?,8'h??,1'b?},
           {36'h132,4'b0???,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = handcode_reg_rdata_WCM_TCAM_CFG;
                 default: read_data = '0;
              endcase
           end
           {36'h132,4'b100?,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = handcode_reg_rdata_WCM_ACTION_CFG_EN;
                 default: read_data = '0;
              endcase
           end
           {36'h132,4'b11??,4'h?,1'b?}: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = handcode_reg_rdata_IDX;
                 default: read_data = '0;
              endcase
           end
           WCM_IP_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = {WCM_IP};
                 default: read_data = '0;
              endcase
           end
           WCM_IM_DECODE_ADDR: begin
              unique casez ({req_fid,req_bar})
                 {B_SB_FID,B_SB_BAR}: read_data = {WCM_IM};
                 default: read_data = '0;
              endcase
           end
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    WCM_IP.reserved0 = '0;
    WCM_IM.reserved0 = '0;
end

// end register RSVD init section }

// ======================================================================
// begin unit parity section {

// end unit parity section }


endmodule
//lintra pop
//lintra pop
