magic
tech scmos
timestamp 988943070
<< nselect >>
rect -87 15 0 86
<< pselect >>
rect 0 15 93 80
<< ndiffusion >>
rect -57 74 -49 75
rect -28 74 -8 75
rect -57 66 -49 71
rect -28 66 -8 71
rect -57 58 -49 63
rect -28 58 -8 63
rect -57 54 -49 55
rect -57 45 -49 46
rect -28 54 -8 55
rect -81 37 -73 38
rect -57 37 -49 42
rect -28 45 -8 46
rect -28 37 -8 42
rect -81 33 -73 34
rect -57 29 -49 34
rect -28 29 -8 34
rect -57 25 -49 26
rect -28 25 -8 26
<< pdiffusion >>
rect 8 66 28 67
rect 49 66 61 67
rect 75 66 87 67
rect 8 58 28 63
rect 8 54 28 55
rect 49 58 61 63
rect 75 62 87 63
rect 8 45 28 46
rect 49 54 61 55
rect 49 45 61 46
rect 83 57 87 62
rect 8 37 28 42
rect 49 37 61 42
rect 8 33 28 34
rect 49 33 61 34
rect 67 30 79 35
rect 67 29 87 30
rect 67 25 87 26
<< ntransistor >>
rect -57 71 -49 74
rect -28 71 -8 74
rect -57 63 -49 66
rect -28 63 -8 66
rect -57 55 -49 58
rect -28 55 -8 58
rect -57 42 -49 45
rect -28 42 -8 45
rect -81 34 -73 37
rect -57 34 -49 37
rect -28 34 -8 37
rect -57 26 -49 29
rect -28 26 -8 29
<< ptransistor >>
rect 8 63 28 66
rect 49 63 61 66
rect 75 63 87 66
rect 8 55 28 58
rect 49 55 61 58
rect 8 42 28 45
rect 49 42 61 45
rect 8 34 28 37
rect 49 34 61 37
rect 67 26 87 29
<< polysilicon >>
rect -61 71 -57 74
rect -49 71 -28 74
rect -8 71 -4 74
rect -61 63 -57 66
rect -49 63 -28 66
rect -8 63 8 66
rect 28 63 49 66
rect 61 63 65 66
rect 71 63 75 66
rect 87 63 92 66
rect -86 50 -82 53
rect -62 55 -57 58
rect -49 55 -45 58
rect -62 50 -59 55
rect -86 37 -83 50
rect -61 45 -59 50
rect -32 55 -28 58
rect -8 55 8 58
rect 28 55 32 58
rect -61 42 -57 45
rect -49 42 -45 45
rect -40 37 -37 50
rect 37 50 40 63
rect 45 55 49 58
rect 61 55 65 58
rect -32 42 -28 45
rect -8 42 8 45
rect 28 42 32 45
rect 63 50 65 55
rect 89 50 92 63
rect 63 45 66 50
rect 45 42 49 45
rect 61 42 66 45
rect 87 47 92 50
rect -86 34 -81 37
rect -73 34 -69 37
rect -61 34 -57 37
rect -49 34 -28 37
rect -8 34 8 37
rect 28 34 49 37
rect 61 34 65 37
rect -61 26 -57 29
rect -49 26 -28 29
rect -8 26 -4 29
rect 63 26 67 29
rect 87 26 91 29
<< ndcontact >>
rect -57 75 -49 83
rect -28 75 -8 83
rect -81 38 -73 46
rect -57 46 -49 54
rect -28 46 -8 54
rect -81 25 -73 33
rect -57 17 -49 25
rect -28 17 -8 25
<< pdcontact >>
rect 8 67 28 75
rect 49 67 61 75
rect 75 67 87 75
rect 8 46 28 54
rect 49 46 61 54
rect 75 54 83 62
rect 8 25 28 33
rect 49 25 61 33
rect 79 30 87 38
rect 67 17 87 25
<< polycontact >>
rect -82 50 -74 58
rect -69 42 -61 50
rect -40 50 -32 58
rect 32 42 40 50
rect 65 50 73 58
rect 79 42 87 50
<< metal1 >>
rect -57 75 -8 83
rect 8 67 87 75
rect -2 58 83 62
rect -82 54 -53 58
rect -82 50 -74 54
rect -69 46 -61 50
rect -57 46 -49 54
rect -40 50 -32 58
rect -28 46 -8 54
rect -81 42 -61 46
rect -2 42 2 58
rect 65 54 83 58
rect 8 46 28 54
rect 32 42 40 50
rect 49 46 61 54
rect 65 50 73 54
rect 79 46 87 50
rect 57 42 87 46
rect -81 38 2 42
rect -81 29 -52 33
rect -81 25 -73 29
rect -57 25 -52 29
rect 8 25 74 33
rect 79 30 87 42
rect -57 17 -8 25
rect 67 17 87 25
<< labels >>
rlabel metal1 -40 50 -32 58 1 a
rlabel metal1 32 42 40 50 1 b
rlabel space -88 15 -28 86 7 ^n
rlabel space 28 15 94 80 3 ^p
rlabel metal1 -81 25 -73 33 1 GND!|pin|s|0
rlabel metal1 8 25 74 33 1 Vdd!|pin|s|1
rlabel metal1 67 17 87 25 1 Vdd!|pin|s|1
rlabel polysilicon -61 26 -57 29 1 _SReset!|pin|w|3|poly
rlabel polysilicon -8 26 -4 29 1 _SReset!|pin|w|3|poly
rlabel polysilicon -61 71 -57 74 1 _SReset!|pin|w|4|poly
rlabel polysilicon -8 71 -4 74 1 _SReset!|pin|w|4|poly
rlabel polysilicon 87 26 91 29 1 _PReset!|pin|w|5|poly
rlabel metal1 -57 75 -8 83 1 GND!|pin|s|1
rlabel metal1 8 67 87 75 1 Vdd!|pin|s|2
rlabel metal1 -82 50 -74 58 1 x|pin|s|0
rlabel metal1 -82 54 -53 58 1 x|pin|s|0
rlabel metal1 -28 46 -8 54 1 x|pin|s|1
rlabel metal1 8 46 28 54 1 x|pin|s|2
rlabel metal1 57 42 87 46 1 x|pin|s|3
rlabel metal1 79 42 87 50 1 x|pin|s|3
rlabel metal1 49 46 61 54 1 x|pin|s|3
rlabel metal1 -57 46 -49 54 1 x|pin|s|0
rlabel metal1 -57 17 -8 25 1 GND!|pin|s|0
<< end >>
