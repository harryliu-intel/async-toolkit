// Copyright (c) 2025 Intel Corporation.  All rights reserved.  See the file COPYRIGHT for more information.
// SPDX-License-Identifier: Apache-2.0

task delay_cclk(int n);
    repeat(n) @(posedge cclk);
endtask
