magic
tech scmos
timestamp 970030046
<< ndiffusion >>
rect -53 75 -45 76
rect -24 75 -8 76
rect -53 67 -45 72
rect -24 67 -8 72
rect -53 59 -45 64
rect -24 59 -8 64
rect -53 55 -45 56
rect -53 46 -45 47
rect -24 55 -8 56
rect -77 38 -69 39
rect -53 38 -45 43
rect -24 46 -8 47
rect -24 38 -8 43
rect -77 34 -69 35
rect -53 30 -45 35
rect -24 30 -8 35
rect -53 26 -45 27
rect -24 26 -8 27
<< pdiffusion >>
rect 8 67 24 68
rect 45 67 57 68
rect 71 67 83 68
rect 8 59 24 64
rect 8 55 24 56
rect 45 59 57 64
rect 71 63 83 64
rect 8 46 24 47
rect 45 55 57 56
rect 45 46 57 47
rect 79 58 83 63
rect 8 38 24 43
rect 45 38 57 43
rect 8 34 24 35
rect 45 34 57 35
rect 63 31 75 36
rect 63 30 83 31
rect 63 26 83 27
<< ntransistor >>
rect -53 72 -45 75
rect -24 72 -8 75
rect -53 64 -45 67
rect -24 64 -8 67
rect -53 56 -45 59
rect -24 56 -8 59
rect -53 43 -45 46
rect -24 43 -8 46
rect -77 35 -69 38
rect -53 35 -45 38
rect -24 35 -8 38
rect -53 27 -45 30
rect -24 27 -8 30
<< ptransistor >>
rect 8 64 24 67
rect 45 64 57 67
rect 71 64 83 67
rect 8 56 24 59
rect 45 56 57 59
rect 8 43 24 46
rect 45 43 57 46
rect 8 35 24 38
rect 45 35 57 38
rect 63 27 83 30
<< polysilicon >>
rect -57 72 -53 75
rect -45 72 -24 75
rect -8 72 -4 75
rect -57 64 -53 67
rect -45 64 -24 67
rect -8 64 8 67
rect 24 64 45 67
rect 57 64 61 67
rect 67 64 71 67
rect 83 64 88 67
rect -82 51 -78 54
rect -58 56 -53 59
rect -45 56 -41 59
rect -58 51 -55 56
rect -82 38 -79 51
rect -57 46 -55 51
rect -28 56 -24 59
rect -8 56 8 59
rect 24 56 28 59
rect -57 43 -53 46
rect -45 43 -41 46
rect -36 38 -33 51
rect 33 51 36 64
rect 41 56 45 59
rect 57 56 61 59
rect -28 43 -24 46
rect -8 43 8 46
rect 24 43 28 46
rect 59 51 61 56
rect 85 51 88 64
rect 59 46 62 51
rect 41 43 45 46
rect 57 43 62 46
rect 83 48 88 51
rect -82 35 -77 38
rect -69 35 -65 38
rect -57 35 -53 38
rect -45 35 -24 38
rect -8 35 8 38
rect 24 35 45 38
rect 57 35 61 38
rect -60 27 -53 30
rect -45 27 -24 30
rect -8 27 -4 30
rect -60 26 -57 27
rect 59 27 63 30
rect 83 27 87 30
<< ndcontact >>
rect -53 76 -45 84
rect -24 76 -8 84
rect -77 39 -69 47
rect -53 47 -45 55
rect -24 47 -8 55
rect -77 26 -69 34
rect -53 18 -45 26
rect -24 18 -8 26
<< pdcontact >>
rect 8 68 24 76
rect 45 68 57 76
rect 71 68 83 76
rect 8 47 24 55
rect 45 47 57 55
rect 71 55 79 63
rect 8 26 24 34
rect 45 26 57 34
rect 75 31 83 39
rect 63 18 83 26
<< psubstratepcontact >>
rect -77 64 -69 72
<< nsubstratencontact >>
rect 92 68 100 76
<< polycontact >>
rect -65 72 -57 80
rect -78 51 -70 59
rect -65 43 -57 51
rect -36 51 -28 59
rect 28 43 36 51
rect 61 51 69 59
rect 75 43 83 51
rect -65 18 -57 26
rect 87 22 95 30
<< metal1 >>
rect -65 72 -57 78
rect -53 78 -21 84
rect -53 76 -8 78
rect 8 76 21 78
rect -77 68 -69 72
rect -53 68 -49 76
rect 8 68 100 76
rect -77 64 -49 68
rect -78 55 -49 59
rect -78 51 -70 55
rect -53 54 -45 55
rect -65 47 -57 51
rect -36 51 -28 60
rect -2 59 79 63
rect -24 54 -8 55
rect -53 47 -45 48
rect -24 47 -8 48
rect -77 43 -57 47
rect -2 43 2 59
rect 61 55 79 59
rect 8 54 24 55
rect 45 54 57 55
rect 8 47 24 48
rect -77 39 2 43
rect 28 42 36 51
rect 53 48 57 54
rect 61 51 69 55
rect 45 47 57 48
rect 75 47 83 51
rect 53 43 83 47
rect -77 30 -48 34
rect -77 26 -69 30
rect -53 26 -48 30
rect 8 32 24 34
rect 45 32 70 34
rect 8 26 70 32
rect 75 31 83 43
rect -65 24 -57 26
rect -53 24 -8 26
rect 8 24 21 26
rect -53 18 -21 24
rect 63 18 83 26
rect 87 24 95 30
<< m2contact >>
rect -65 78 -57 84
rect -21 78 -3 84
rect 3 78 21 84
rect -36 60 -28 66
rect -53 48 -45 54
rect -24 48 -8 54
rect 8 48 24 54
rect 45 48 53 54
rect 28 36 36 42
rect -65 18 -57 24
rect -21 18 -3 24
rect 3 18 21 24
rect 87 18 95 24
<< metal2 >>
rect -65 78 -27 84
rect -36 60 0 66
rect -53 48 53 54
rect 0 36 36 42
rect -65 18 -27 24
rect 27 18 95 24
<< m3contact >>
rect -21 78 -3 84
rect 3 78 21 84
rect -21 18 -3 24
rect 3 18 21 24
<< metal3 >>
rect -21 15 -3 87
rect 3 15 21 87
<< labels >>
rlabel metal1 12 72 12 72 5 Vdd!
rlabel metal1 12 30 12 30 1 Vdd!
rlabel m2contact -12 80 -12 80 5 GND!
rlabel m2contact -12 22 -12 22 1 GND!
rlabel metal1 -49 80 -49 80 5 GND!
rlabel polysilicon -54 73 -54 73 1 _SReset!
rlabel metal1 -49 22 -49 22 1 GND!
rlabel polysilicon -54 28 -54 28 1 _SReset!
rlabel metal1 51 72 51 72 5 Vdd!
rlabel metal1 51 30 51 30 1 Vdd!
rlabel polysilicon -54 65 -54 65 3 b
rlabel polysilicon -54 36 -54 36 3 a
rlabel metal1 77 72 77 72 5 Vdd!
rlabel metal1 75 22 75 22 5 Vdd!
rlabel polysilicon 84 29 84 29 7 _PReset!
rlabel metal1 79 47 79 47 5 x
rlabel polysilicon 58 65 58 65 7 b
rlabel polysilicon 58 36 58 36 7 a
rlabel metal2 0 36 0 42 3 b
rlabel metal2 0 60 0 66 7 a
rlabel metal2 91 21 91 21 7 _PReset!
rlabel metal2 -61 81 -61 81 1 _SReset!
rlabel metal1 96 72 96 72 7 Vdd!
rlabel metal1 -73 30 -73 30 1 GND!
rlabel metal2 -61 21 -61 21 1 _SReset!
rlabel metal1 -73 68 -73 68 1 GND!
rlabel metal1 -74 55 -74 55 3 x
rlabel space -83 17 -24 85 7 ^n
rlabel space 24 17 101 77 3 ^p
rlabel metal2 27 18 27 24 7 ^p
rlabel metal2 -27 18 -27 24 3 ^n
rlabel metal2 -27 78 -27 84 3 ^n
rlabel metal2 -32 63 -32 63 1 a
rlabel metal2 49 51 49 51 1 x
rlabel metal2 16 51 16 51 1 x
rlabel metal2 -16 51 -16 51 1 x
rlabel metal2 -49 51 -49 51 1 x
rlabel metal2 32 39 32 39 1 b
<< end >>
